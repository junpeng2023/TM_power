module netlist_1 (clk,
    in0,
    in1,
    in10,
    in11,
    in12,
    in13,
    in14,
    in15,
    in16,
    in17,
    in18,
    in19,
    in2,
    in20,
    in21,
    in22,
    in23,
    in24,
    in3,
    in4,
    in5,
    in6,
    in7,
    in8,
    in9,
    out0,
    out1,
    out10,
    out11,
    out12,
    out13,
    out14,
    out15,
    out16,
    out17,
    out18,
    out19,
    out2,
    out20,
    out21,
    out22,
    out23,
    out24,
    out3,
    out4,
    out5,
    out6,
    out7,
    out8,
    out9,
    rst);
 input clk;
 input in0;
 input in1;
 input in10;
 input in11;
 input in12;
 input in13;
 input in14;
 input in15;
 input in16;
 input in17;
 input in18;
 input in19;
 input in2;
 input in20;
 input in21;
 input in22;
 input in23;
 input in24;
 input in3;
 input in4;
 input in5;
 input in6;
 input in7;
 input in8;
 input in9;
 output out0;
 output out1;
 output out10;
 output out11;
 output out12;
 output out13;
 output out14;
 output out15;
 output out16;
 output out17;
 output out18;
 output out19;
 output out2;
 output out20;
 output out21;
 output out22;
 output out23;
 output out24;
 output out3;
 output out4;
 output out5;
 output out6;
 output out7;
 output out8;
 output out9;
 input rst;

 wire net0;
 wire net1;
 wire net10;
 wire net100;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net101;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net102;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net103;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net63;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net64;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net65;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net66;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net67;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net68;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net69;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net7;
 wire net70;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net71;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net72;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net73;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net74;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net75;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net76;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net77;
 wire net770;
 wire net771;
 wire net772;
 wire net774;
 wire net775;
 wire net776;
 wire net778;
 wire net779;
 wire net78;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net79;
 wire net790;
 wire net791;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net8;
 wire net80;
 wire net800;
 wire net802;
 wire net803;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net81;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net82;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net83;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net84;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net85;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net86;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net87;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net88;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net89;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net9;
 wire net90;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net91;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net92;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net93;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net94;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net95;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net96;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net97;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net98;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net99;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net773;
 wire net777;
 wire net792;
 wire net801;
 wire net804;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire clknet_leaf_0_clk;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire clknet_0_net1028;
 wire clknet_1_0__leaf_net1028;
 wire clknet_1_1__leaf_net1028;
 wire clknet_0_net805;
 wire clknet_1_0__leaf_net805;
 wire clknet_1_1__leaf_net805;
 wire clknet_0_net723;
 wire clknet_1_0__leaf_net723;
 wire clknet_1_1__leaf_net723;
 wire clknet_0_net727;
 wire clknet_1_0__leaf_net727;
 wire clknet_1_1__leaf_net727;
 wire clknet_0_net729;
 wire clknet_1_0__leaf_net729;
 wire clknet_1_1__leaf_net729;
 wire clknet_0_net722;
 wire clknet_1_0__leaf_net722;
 wire clknet_1_1__leaf_net722;
 wire clknet_0_net725;
 wire clknet_1_0__leaf_net725;
 wire clknet_1_1__leaf_net725;
 wire clknet_0_net768;
 wire clknet_1_0__leaf_net768;
 wire clknet_1_1__leaf_net768;
 wire clknet_0_net755;
 wire clknet_1_0__leaf_net755;
 wire clknet_1_1__leaf_net755;
 wire clknet_0_net756;
 wire clknet_1_0__leaf_net756;
 wire clknet_1_1__leaf_net756;
 wire clknet_0_net1026;
 wire clknet_1_0__leaf_net1026;
 wire clknet_1_1__leaf_net1026;
 wire clknet_0_net759;
 wire clknet_1_0__leaf_net759;
 wire clknet_1_1__leaf_net759;
 wire clknet_0_net628;
 wire clknet_1_0__leaf_net628;
 wire clknet_1_1__leaf_net628;
 wire clknet_0_net747;
 wire clknet_1_0__leaf_net747;
 wire clknet_1_1__leaf_net747;
 wire clknet_0_net728;
 wire clknet_1_0__leaf_net728;
 wire clknet_1_1__leaf_net728;
 wire clknet_0_net1027;
 wire clknet_1_0__leaf_net1027;
 wire clknet_1_1__leaf_net1027;
 wire clknet_0_net313;
 wire clknet_1_0__leaf_net313;
 wire clknet_1_1__leaf_net313;
 wire clknet_0_net911;
 wire clknet_1_0__leaf_net911;
 wire clknet_1_1__leaf_net911;
 wire clknet_0_net450;
 wire clknet_1_0__leaf_net450;
 wire clknet_1_1__leaf_net450;
 wire clknet_0_net462;
 wire clknet_1_0__leaf_net462;
 wire clknet_1_1__leaf_net462;
 wire clknet_0_net454;
 wire clknet_1_0__leaf_net454;
 wire clknet_1_1__leaf_net454;
 wire clknet_0_net451;
 wire clknet_1_0__leaf_net451;
 wire clknet_1_1__leaf_net451;
 wire clknet_0_net910;
 wire clknet_1_0__leaf_net910;
 wire clknet_1_1__leaf_net910;
 wire clknet_0_net909;
 wire clknet_1_0__leaf_net909;
 wire clknet_1_1__leaf_net909;
 wire clknet_0_net1007;
 wire clknet_1_0__leaf_net1007;
 wire clknet_1_1__leaf_net1007;
 wire clknet_0_net379;
 wire clknet_1_0__leaf_net379;
 wire clknet_1_1__leaf_net379;
 wire clknet_0_net376;
 wire clknet_1_0__leaf_net376;
 wire clknet_1_1__leaf_net376;
 wire clknet_0_net377;
 wire clknet_1_0__leaf_net377;
 wire clknet_1_1__leaf_net377;
 wire clknet_0_net987;
 wire clknet_1_0__leaf_net987;
 wire clknet_1_1__leaf_net987;
 wire clknet_0_net700;
 wire clknet_1_0__leaf_net700;
 wire clknet_1_1__leaf_net700;
 wire clknet_0_net720;
 wire clknet_1_0__leaf_net720;
 wire clknet_1_1__leaf_net720;
 wire clknet_0_net705;
 wire clknet_1_0__leaf_net705;
 wire clknet_1_1__leaf_net705;
 wire clknet_0_net702;
 wire clknet_1_0__leaf_net702;
 wire clknet_1_1__leaf_net702;
 wire clknet_0_net701;
 wire clknet_1_0__leaf_net701;
 wire clknet_1_1__leaf_net701;
 wire clknet_0_net609;
 wire clknet_1_0__leaf_net609;
 wire clknet_1_1__leaf_net609;
 wire clknet_0_net613;
 wire clknet_1_0__leaf_net613;
 wire clknet_1_1__leaf_net613;
 wire clknet_0_net622;
 wire clknet_1_0__leaf_net622;
 wire clknet_1_1__leaf_net622;
 wire clknet_0_net615;
 wire clknet_1_0__leaf_net615;
 wire clknet_1_1__leaf_net615;
 wire clknet_0_net610;
 wire clknet_1_0__leaf_net610;
 wire clknet_1_1__leaf_net610;
 wire clknet_0_net626;
 wire clknet_1_0__leaf_net626;
 wire clknet_1_1__leaf_net626;
 wire clknet_0_net611;
 wire clknet_1_0__leaf_net611;
 wire clknet_1_1__leaf_net611;
 wire clknet_0_net950;
 wire clknet_1_0__leaf_net950;
 wire clknet_1_1__leaf_net950;
 wire clknet_0_net536;
 wire clknet_1_0__leaf_net536;
 wire clknet_1_1__leaf_net536;
 wire clknet_0_net1055;
 wire clknet_1_0__leaf_net1055;
 wire clknet_1_1__leaf_net1055;
 wire clknet_0_net1057;
 wire clknet_1_0__leaf_net1057;
 wire clknet_1_1__leaf_net1057;
 wire clknet_0_net533;
 wire clknet_1_0__leaf_net533;
 wire clknet_1_1__leaf_net533;
 wire clknet_0_net526;
 wire clknet_1_0__leaf_net526;
 wire clknet_1_1__leaf_net526;
 wire clknet_0_net520;
 wire clknet_1_0__leaf_net520;
 wire clknet_1_1__leaf_net520;
 wire clknet_0_net523;
 wire clknet_1_0__leaf_net523;
 wire clknet_1_1__leaf_net523;
 wire clknet_0_net948;
 wire clknet_1_0__leaf_net948;
 wire clknet_1_1__leaf_net948;
 wire clknet_0_net633;
 wire clknet_1_0__leaf_net633;
 wire clknet_1_1__leaf_net633;
 wire clknet_0_net639;
 wire clknet_1_0__leaf_net639;
 wire clknet_1_1__leaf_net639;
 wire clknet_0_net518;
 wire clknet_1_0__leaf_net518;
 wire clknet_1_1__leaf_net518;
 wire clknet_0_net931;
 wire clknet_1_0__leaf_net931;
 wire clknet_1_1__leaf_net931;
 wire clknet_0_net549;
 wire clknet_1_0__leaf_net549;
 wire clknet_1_1__leaf_net549;
 wire clknet_0_net556;
 wire clknet_1_0__leaf_net556;
 wire clknet_1_1__leaf_net556;
 wire clknet_0_net550;
 wire clknet_1_0__leaf_net550;
 wire clknet_1_1__leaf_net550;
 wire clknet_0_net560;
 wire clknet_1_0__leaf_net560;
 wire clknet_1_1__leaf_net560;
 wire clknet_0_net553;
 wire clknet_1_0__leaf_net553;
 wire clknet_1_1__leaf_net553;
 wire clknet_0_net545;
 wire clknet_1_0__leaf_net545;
 wire clknet_1_1__leaf_net545;
 wire clknet_0_net541;
 wire clknet_1_0__leaf_net541;
 wire clknet_1_1__leaf_net541;
 wire clknet_0_net544;
 wire clknet_1_0__leaf_net544;
 wire clknet_1_1__leaf_net544;
 wire clknet_0_net543;
 wire clknet_1_0__leaf_net543;
 wire clknet_1_1__leaf_net543;
 wire clknet_0_net538;
 wire clknet_1_0__leaf_net538;
 wire clknet_1_1__leaf_net538;
 wire clknet_0_net540;
 wire clknet_1_0__leaf_net540;
 wire clknet_1_1__leaf_net540;
 wire clknet_0_net539;
 wire clknet_1_0__leaf_net539;
 wire clknet_1_1__leaf_net539;
 wire clknet_0_net930;
 wire clknet_1_0__leaf_net930;
 wire clknet_1_1__leaf_net930;
 wire clknet_0_net929;
 wire clknet_1_0__leaf_net929;
 wire clknet_1_1__leaf_net929;
 wire clknet_0_net141;
 wire clknet_1_0__leaf_net141;
 wire clknet_1_1__leaf_net141;
 wire clknet_0_net890;
 wire clknet_1_0__leaf_net890;
 wire clknet_1_1__leaf_net890;
 wire clknet_0_net262;
 wire clknet_1_0__leaf_net262;
 wire clknet_1_1__leaf_net262;
 wire clknet_0_net137;
 wire clknet_1_0__leaf_net137;
 wire clknet_1_1__leaf_net137;
 wire clknet_0_net139;
 wire clknet_1_0__leaf_net139;
 wire clknet_1_1__leaf_net139;
 wire clknet_0_net138;
 wire clknet_1_0__leaf_net138;
 wire clknet_1_1__leaf_net138;
 wire clknet_0_net873;
 wire clknet_1_0__leaf_net873;
 wire clknet_1_1__leaf_net873;
 wire clknet_0_net60;
 wire clknet_1_0__leaf_net60;
 wire clknet_1_1__leaf_net60;
 wire clknet_0_net872;
 wire clknet_1_0__leaf_net872;
 wire clknet_1_1__leaf_net872;
 wire clknet_0_net67;
 wire clknet_1_0__leaf_net67;
 wire clknet_1_1__leaf_net67;
 wire clknet_0_net70;
 wire clknet_1_0__leaf_net70;
 wire clknet_1_1__leaf_net70;
 wire clknet_0_net68;
 wire clknet_1_0__leaf_net68;
 wire clknet_1_1__leaf_net68;
 wire clknet_0_net75;
 wire clknet_1_0__leaf_net75;
 wire clknet_1_1__leaf_net75;
 wire clknet_0_net69;
 wire clknet_1_0__leaf_net69;
 wire clknet_1_1__leaf_net69;
 wire clknet_0_net48;
 wire clknet_1_0__leaf_net48;
 wire clknet_1_1__leaf_net48;
 wire clknet_0_net159;
 wire clknet_1_0__leaf_net159;
 wire clknet_1_1__leaf_net159;
 wire clknet_0_net167;
 wire clknet_1_0__leaf_net167;
 wire clknet_1_1__leaf_net167;
 wire clknet_0_net161;
 wire clknet_1_0__leaf_net161;
 wire clknet_1_1__leaf_net161;
 wire clknet_0_net160;
 wire clknet_1_0__leaf_net160;
 wire clknet_1_1__leaf_net160;
 wire clknet_0_net871;
 wire clknet_1_0__leaf_net871;
 wire clknet_1_1__leaf_net871;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;

 sky130_fd_sc_hd__mux4_1 c100 (.A0(net86),
    .A1(net66),
    .A2(net74),
    .A3(clknet_1_1__leaf_net70),
    .S0(clknet_1_1__leaf_net69),
    .S1(net879),
    .X(net88));
 sky130_fd_sc_hd__mux4_1 c101 (.A0(net71),
    .A1(net83),
    .A2(net76),
    .A3(net86),
    .S0(net73),
    .S1(net879),
    .X(net89));
 sky130_fd_sc_hd__mux4_1 c102 (.A0(net81),
    .A1(net89),
    .A2(net72),
    .A3(net86),
    .S0(net82),
    .S1(net879),
    .X(net90));
 sky130_fd_sc_hd__mux4_1 c103 (.A0(net79),
    .A1(net90),
    .A2(net89),
    .A3(clknet_1_1__leaf_net68),
    .S0(net879),
    .S1(net881),
    .X(net91));
 sky130_fd_sc_hd__mux4_1 c104 (.A0(net91),
    .A1(net89),
    .A2(net90),
    .A3(net85),
    .S0(net82),
    .S1(net880),
    .X(net92));
 sky130_fd_sc_hd__buf_1 c105 (.A(net882),
    .X(net93));
 sky130_fd_sc_hd__clkbuf_2 c106 (.A(net93),
    .X(net94));
 sky130_fd_sc_hd__and2_1 c107 (.A(net94),
    .B(net93),
    .X(net95));
 sky130_fd_sc_hd__and2_1 c108 (.A(net93),
    .B(net94),
    .X(net96));
 sky130_fd_sc_hd__dfbbn_1 c109 (.CLK_N(clknet_leaf_21_clk),
    .D(net95),
    .RESET_B(net96),
    .SET_B(net94),
    .Q(net97));
 sky130_fd_sc_hd__clkbuf_1 c110 (.A(net806),
    .X(net98));
 sky130_fd_sc_hd__dfbbp_1 c111 (.CLK(clknet_leaf_22_clk),
    .D(net95),
    .RESET_B(net96),
    .SET_B(net1170),
    .Q(net100),
    .Q_N(net99));
 sky130_fd_sc_hd__clkbuf_1 c112 (.A(net806),
    .X(net101));
 sky130_fd_sc_hd__buf_1 c113 (.A(net840),
    .X(net102));
 sky130_fd_sc_hd__buf_1 c114 (.A(net848),
    .X(net103));
 sky130_fd_sc_hd__and3_1 c115 (.A(net101),
    .B(net103),
    .C(net93),
    .X(net104));
 sky130_fd_sc_hd__a2111o_1 c116 (.A1(net100),
    .A2(net94),
    .B1(net102),
    .C1(net93),
    .D1(net103),
    .X(net105));
 sky130_fd_sc_hd__and2_1 c117 (.A(net103),
    .B(net102),
    .X(net106));
 sky130_fd_sc_hd__and3_2 c118 (.A(net98),
    .B(net101),
    .C(net106),
    .X(net107));
 sky130_fd_sc_hd__and3_1 c119 (.A(net107),
    .B(net103),
    .C(net102),
    .X(net108));
 sky130_fd_sc_hd__and2_0 c120 (.A(net103),
    .B(net107),
    .X(net109));
 sky130_fd_sc_hd__mux4_1 c121 (.A0(net105),
    .A1(net107),
    .A2(net106),
    .A3(net103),
    .S0(net94),
    .S1(net99),
    .X(net110));
 sky130_fd_sc_hd__and3_1 c122 (.A(net106),
    .B(net107),
    .C(net884),
    .X(net111));
 sky130_fd_sc_hd__mux4_1 c123 (.A0(net108),
    .A1(net94),
    .A2(net106),
    .A3(net102),
    .S0(net107),
    .S1(net883),
    .X(net112));
 sky130_fd_sc_hd__mux4_1 c124 (.A0(net109),
    .A1(net111),
    .A2(net95),
    .A3(net94),
    .S0(net107),
    .S1(net883),
    .X(net113));
 sky130_fd_sc_hd__mux4_1 c125 (.A0(net107),
    .A1(net103),
    .A2(net95),
    .A3(net884),
    .S0(net885),
    .S1(net1155),
    .X(net114));
 sky130_fd_sc_hd__and2_1 c126 (.A(net1038),
    .B(net773),
    .X(net115));
 sky130_fd_sc_hd__and2_2 c127 (.A(net115),
    .B(net1038),
    .X(net116));
 sky130_fd_sc_hd__and2_0 c128 (.A(net116),
    .B(net777),
    .X(net117));
 sky130_fd_sc_hd__and2_0 c129 (.A(net115),
    .B(net116),
    .X(net118));
 sky130_fd_sc_hd__and2_2 c130 (.A(net116),
    .B(net1038),
    .X(net119));
 sky130_fd_sc_hd__and2_1 c131 (.A(net116),
    .B(net1050),
    .X(net120));
 sky130_fd_sc_hd__clkbuf_2 c132 (.A(net781),
    .X(net121));
 sky130_fd_sc_hd__and2_0 c133 (.A(net121),
    .B(net1038),
    .X(net122));
 sky130_fd_sc_hd__clkbuf_2 c134 (.A(net1009),
    .X(net123));
 sky130_fd_sc_hd__clkbuf_1 c135 (.A(net1008),
    .X(net124));
 sky130_fd_sc_hd__or4bb_1 c136 (.A(net123),
    .B(net124),
    .C_N(net116),
    .D_N(net121),
    .X(net125));
 sky130_fd_sc_hd__and2_0 c137 (.A(net121),
    .B(net123),
    .X(net126));
 sky130_fd_sc_hd__sdfxbp_1 c138 (.CLK(clknet_leaf_1_clk),
    .D(net120),
    .SCD(net121),
    .SCE(net123),
    .Q(net127));
 sky130_fd_sc_hd__clkbuf_1 c139 (.A(net782),
    .X(net128));
 sky130_fd_sc_hd__mux4_1 c140 (.A0(net124),
    .A1(net125),
    .A2(net121),
    .A3(net115),
    .S0(net123),
    .S1(net126),
    .X(net129));
 sky130_fd_sc_hd__and3_1 c141 (.A(net122),
    .B(net116),
    .C(net121),
    .X(net130));
 sky130_fd_sc_hd__mux4_1 c142 (.A0(net128),
    .A1(net1051),
    .A2(net115),
    .A3(net130),
    .S0(net119),
    .S1(net121),
    .X(net131));
 sky130_fd_sc_hd__sdfxbp_1 c143 (.CLK(clknet_leaf_1_clk),
    .D(net130),
    .SCD(net126),
    .SCE(net121),
    .Q(net133),
    .Q_N(net132));
 sky130_fd_sc_hd__mux4_1 c144 (.A0(net1189),
    .A1(net132),
    .A2(net119),
    .A3(net130),
    .S0(net123),
    .S1(net116),
    .X(net134));
 sky130_fd_sc_hd__mux4_1 c145 (.A0(net1037),
    .A1(net130),
    .A2(net123),
    .A3(net121),
    .S0(net119),
    .S1(clknet_1_1__leaf_net890),
    .X(net135));
 sky130_fd_sc_hd__mux4_1 c146 (.A0(net133),
    .A1(net128),
    .A2(net123),
    .A3(net121),
    .S0(net888),
    .S1(clknet_1_0__leaf_net890),
    .X(net136));
 sky130_fd_sc_hd__and2_0 c147 (.A(net1080),
    .B(net889),
    .X(net137));
 sky130_fd_sc_hd__and2_0 c148 (.A(clknet_1_0__leaf_net137),
    .B(net1109),
    .X(net138));
 sky130_fd_sc_hd__and3_1 c149 (.A(net1080),
    .B(net1035),
    .C(clknet_1_0__leaf_net137),
    .X(net139));
 sky130_fd_sc_hd__clkbuf_2 c150 (.X(net140));
 sky130_fd_sc_hd__and2_0 c151 (.A(net140),
    .B(net891),
    .X(net141));
 sky130_fd_sc_hd__clkbuf_1 c152 (.A(net800),
    .X(net142));
 sky130_fd_sc_hd__dlymetal6s2s_1 c153 (.A(net1014),
    .X(net143));
 sky130_fd_sc_hd__clkbuf_1 c154 (.A(net1016),
    .X(net144));
 sky130_fd_sc_hd__and2_0 c155 (.A(net144),
    .B(net143),
    .X(net145));
 sky130_fd_sc_hd__sdfrtp_1 c156 (.CLK(clknet_leaf_7_clk),
    .D(net140),
    .RESET_B(clknet_1_0__leaf_net138),
    .SCD(clknet_1_0__leaf_net141),
    .SCE(clknet_1_0__leaf_net139),
    .Q(net146));
 sky130_fd_sc_hd__and2_0 c157 (.A(net142),
    .B(clknet_1_1__leaf_net137),
    .X(net147));
 sky130_fd_sc_hd__and2_0 c158 (.A(net145),
    .B(clknet_1_1__leaf_net137),
    .X(net148));
 sky130_fd_sc_hd__sdfbbn_1 c159 (.CLK_N(clknet_leaf_7_clk),
    .D(net118),
    .RESET_B(net143),
    .SCD(clknet_1_1__leaf_net141),
    .SCE(clknet_1_1__leaf_net139),
    .SET_B(clknet_1_0__leaf_net137),
    .Q(net150),
    .Q_N(net149));
 sky130_fd_sc_hd__sdfbbp_1 c160 (.CLK(clknet_leaf_7_clk),
    .D(clknet_1_0__leaf_net137),
    .RESET_B(net150),
    .SCD(net143),
    .SCE(clknet_1_1__leaf_net139),
    .SET_B(net140),
    .Q(net151));
 sky130_fd_sc_hd__buf_1 c161 (.A(clknet_1_0__leaf_net1027),
    .X(net152));
 sky130_fd_sc_hd__sdfxtp_1 c162 (.CLK(clknet_leaf_7_clk),
    .D(net147),
    .SCD(net1152),
    .SCE(net143),
    .Q(net153));
 sky130_fd_sc_hd__and3_1 c163 (.A(net146),
    .B(net153),
    .C(net149),
    .X(net154));
 sky130_fd_sc_hd__sdfrtp_1 c164 (.CLK(clknet_leaf_6_clk),
    .D(net148),
    .RESET_B(clknet_1_1__leaf_net139),
    .SCD(clknet_1_1__leaf_net137),
    .SCE(net146),
    .Q(net155));
 sky130_fd_sc_hd__and3_1 c165 (.A(net155),
    .B(net154),
    .C(net8),
    .X(net156));
 sky130_fd_sc_hd__mux4_1 c166 (.A0(net151),
    .A1(net156),
    .A2(net150),
    .A3(net155),
    .S0(net143),
    .S1(clknet_1_1__leaf_net137),
    .X(net157));
 sky130_fd_sc_hd__mux4_1 c167 (.A0(net152),
    .A1(net157),
    .A2(net140),
    .A3(net156),
    .S0(net146),
    .S1(net155),
    .X(net158));
 sky130_fd_sc_hd__and2_0 c168 (.A(clknet_1_0__leaf_net872),
    .B(net893),
    .X(net159));
 sky130_fd_sc_hd__and2_0 c169 (.A(clknet_1_0__leaf_net159),
    .B(net892),
    .X(net160));
 sky130_fd_sc_hd__and2_0 c170 (.A(clknet_1_0__leaf_net159),
    .B(clknet_1_0__leaf_net160),
    .X(net161));
 sky130_fd_sc_hd__buf_1 c171 (.A(net787),
    .X(net162));
 sky130_fd_sc_hd__clkbuf_2 c172 (.A(net787),
    .X(net163));
 sky130_fd_sc_hd__sdfxtp_1 c173 (.CLK(clknet_leaf_5_clk),
    .D(clknet_1_0__leaf_net160),
    .SCD(clknet_1_0__leaf_net161),
    .SCE(net893),
    .Q(net164));
 sky130_fd_sc_hd__and2_0 c174 (.A(net163),
    .B(clknet_1_0__leaf_net872),
    .X(net165));
 sky130_fd_sc_hd__and2_0 c175 (.A(net153),
    .B(clknet_1_0__leaf_net872),
    .X(net166));
 sky130_fd_sc_hd__and2_0 c176 (.A(net162),
    .B(clknet_1_0__leaf_net159),
    .X(net167));
 sky130_fd_sc_hd__and3_1 c177 (.A(clknet_1_0__leaf_net167),
    .B(clknet_1_1__leaf_net159),
    .C(clknet_1_0__leaf_net872),
    .X(net168));
 sky130_fd_sc_hd__and3_1 c178 (.A(net163),
    .B(net162),
    .C(net164),
    .X(net169));
 sky130_fd_sc_hd__and3_1 c179 (.A(net166),
    .B(net163),
    .C(net169),
    .X(net170));
 sky130_fd_sc_hd__or4bb_1 c180 (.A(clknet_1_0__leaf_net160),
    .B(net162),
    .C_N(net163),
    .D_N(net169),
    .X(net171));
 sky130_fd_sc_hd__or4bb_1 c181 (.A(net164),
    .B(net169),
    .C_N(net153),
    .D_N(clknet_1_0__leaf_net167),
    .X(net172));
 sky130_fd_sc_hd__buf_1 c182 (.A(net1024),
    .X(net173));
 sky130_fd_sc_hd__mux4_1 c183 (.A0(net172),
    .A1(net173),
    .A2(net169),
    .A3(clknet_1_1__leaf_net159),
    .S0(net163),
    .S1(net162),
    .X(net174));
 sky130_fd_sc_hd__or4bb_1 c184 (.A(net165),
    .B(clknet_1_1__leaf_net167),
    .C_N(net153),
    .D_N(net894),
    .X(net175));
 sky130_fd_sc_hd__or4bb_1 c185 (.A(net162),
    .B(net163),
    .C_N(net173),
    .D_N(net895),
    .X(net176));
 sky130_fd_sc_hd__sdfrtp_1 c186 (.CLK(clknet_leaf_16_clk),
    .D(net170),
    .RESET_B(net175),
    .SCD(net173),
    .SCE(net894),
    .Q(net177));
 sky130_fd_sc_hd__mux4_1 c187 (.A0(net177),
    .A1(net171),
    .A2(net176),
    .A3(net173),
    .S0(net163),
    .S1(net162),
    .X(net178));
 sky130_fd_sc_hd__sdfsbp_1 c188 (.CLK(clknet_leaf_16_clk),
    .D(clknet_1_1__leaf_net161),
    .SCD(clknet_1_1__leaf_net160),
    .SCE(net895),
    .SET_B(net1087),
    .Q(net180),
    .Q_N(net179));
 sky130_fd_sc_hd__and2_1 c189 (.A(net180),
    .B(net51),
    .X(net181));
 sky130_fd_sc_hd__and2_0 c190 (.A(net181),
    .B(net66),
    .X(net182));
 sky130_fd_sc_hd__and2_0 c191 (.A(net181),
    .B(net179),
    .X(net183));
 sky130_fd_sc_hd__and2_2 c192 (.A(net182),
    .B(net66),
    .X(net184));
 sky130_fd_sc_hd__buf_1 c193 (.A(net778),
    .X(net185));
 sky130_fd_sc_hd__and2_1 c194 (.A(net185),
    .B(net1074),
    .X(net186));
 sky130_fd_sc_hd__clkbuf_4 c195 (.A(net1020),
    .X(net187));
 sky130_fd_sc_hd__clkbuf_1 c196 (.A(net778),
    .X(net188));
 sky130_fd_sc_hd__and2_1 c197 (.A(net51),
    .B(net1074),
    .X(net189));
 sky130_fd_sc_hd__clkbuf_2 c198 (.A(net1017),
    .X(net190));
 sky130_fd_sc_hd__sdfsbp_1 c199 (.CLK(clknet_leaf_15_clk),
    .D(net1074),
    .SCD(net190),
    .SCE(net189),
    .SET_B(net1108),
    .Q(net192),
    .Q_N(net191));
 sky130_fd_sc_hd__sdfstp_1 c200 (.CLK(clknet_leaf_12_clk),
    .D(net189),
    .SCD(net187),
    .SCE(net190),
    .SET_B(net1074),
    .Q(net193));
 sky130_fd_sc_hd__sdfstp_1 c201 (.CLK(clknet_leaf_15_clk),
    .D(net188),
    .SCD(net1074),
    .SCE(net184),
    .SET_B(net1100),
    .Q(net194));
 sky130_fd_sc_hd__a2111o_1 c202 (.A1(net194),
    .A2(net187),
    .B1(net51),
    .C1(net193),
    .D1(net1074),
    .X(net195));
 sky130_fd_sc_hd__mux4_1 c203 (.A0(net190),
    .A1(net189),
    .A2(net193),
    .A3(net1074),
    .S0(net187),
    .S1(net194),
    .X(net196));
 sky130_fd_sc_hd__mux4_1 c204 (.A0(net192),
    .A1(net194),
    .A2(net193),
    .A3(net181),
    .S0(net1074),
    .S1(net897),
    .X(net197));
 sky130_fd_sc_hd__mux4_1 c205 (.A0(net197),
    .A1(net193),
    .A2(net182),
    .A3(net195),
    .S0(net190),
    .S1(net897),
    .X(net198));
 sky130_fd_sc_hd__mux4_1 c206 (.A0(net191),
    .A1(net197),
    .A2(net50),
    .A3(net187),
    .S0(net897),
    .S1(net898),
    .X(net199));
 sky130_fd_sc_hd__mux4_1 c207 (.A0(net193),
    .A1(net190),
    .A2(net185),
    .A3(net179),
    .S0(net898),
    .S1(net899),
    .X(net200));
 sky130_fd_sc_hd__mux4_1 c208 (.A0(net195),
    .A1(net197),
    .A2(net1074),
    .A3(net193),
    .S0(net897),
    .S1(net1173),
    .X(net201));
 sky130_fd_sc_hd__mux4_1 c209 (.A0(net200),
    .A1(net197),
    .A2(net1074),
    .A3(net187),
    .S0(net898),
    .S1(net899),
    .X(net202));
 sky130_fd_sc_hd__buf_1 c210 (.A(net802),
    .X(net203));
 sky130_fd_sc_hd__and2_1 c211 (.A(net187),
    .B(net203),
    .X(net204));
 sky130_fd_sc_hd__and2_0 c212 (.A(net204),
    .B(net901),
    .X(net205));
 sky130_fd_sc_hd__and2_1 c213 (.A(net205),
    .B(net203),
    .X(net206));
 sky130_fd_sc_hd__and2_2 c214 (.A(net205),
    .B(net203),
    .X(net207));
 sky130_fd_sc_hd__clkbuf_1 c215 (.A(net802),
    .X(net208));
 sky130_fd_sc_hd__buf_1 c216 (.A(net831),
    .X(net209));
 sky130_fd_sc_hd__clkbuf_2 c217 (.A(net821),
    .X(net210));
 sky130_fd_sc_hd__and2_1 c218 (.A(net203),
    .B(net209),
    .X(net211));
 sky130_fd_sc_hd__clkbuf_1 c219 (.A(net1019),
    .X(net212));
 sky130_fd_sc_hd__and2_1 c220 (.A(net210),
    .B(net211),
    .X(net213));
 sky130_fd_sc_hd__sdfbbn_1 c221 (.CLK_N(clknet_leaf_19_clk),
    .D(net212),
    .RESET_B(net204),
    .SCD(net207),
    .SCE(net210),
    .SET_B(net209),
    .Q(net215),
    .Q_N(net214));
 sky130_fd_sc_hd__and2_0 c222 (.A(net215),
    .B(net208),
    .X(net216));
 sky130_fd_sc_hd__sdfstp_1 c223 (.CLK(clknet_leaf_20_clk),
    .D(net211),
    .SCD(net209),
    .SCE(net213),
    .SET_B(net1122),
    .Q(net217));
 sky130_fd_sc_hd__sedfxbp_1 c224 (.CLK(clknet_leaf_20_clk),
    .D(net195),
    .DE(net213),
    .SCD(net210),
    .SCE(net207),
    .Q(net219),
    .Q_N(net218));
 sky130_fd_sc_hd__and2_0 c225 (.A(net210),
    .B(net219),
    .X(net220));
 sky130_fd_sc_hd__sedfxbp_1 c226 (.CLK(clknet_leaf_19_clk),
    .D(net1175),
    .DE(net206),
    .SCD(net214),
    .SCE(net218),
    .Q(net222),
    .Q_N(net221));
 sky130_fd_sc_hd__mux4_1 c227 (.A0(net216),
    .A1(net212),
    .A2(net221),
    .A3(net220),
    .S0(net211),
    .S1(net210),
    .X(net223));
 sky130_fd_sc_hd__mux4_1 c228 (.A0(net206),
    .A1(net216),
    .A2(net223),
    .A3(net217),
    .S0(net211),
    .S1(net210),
    .X(net224));
 sky130_fd_sc_hd__sdfbbn_1 c229 (.CLK_N(clknet_leaf_19_clk),
    .D(net204),
    .RESET_B(net223),
    .SCD(net219),
    .SCE(net207),
    .SET_B(net903),
    .Q(net226),
    .Q_N(net225));
 sky130_fd_sc_hd__mux4_2 c230 (.A0(net223),
    .A1(net220),
    .A2(net210),
    .A3(net225),
    .S0(net218),
    .S1(net902),
    .X(net227));
 sky130_fd_sc_hd__buf_2 c231 (.X(net228));
 sky130_fd_sc_hd__and2_2 c232 (.A(net1078),
    .B(net225),
    .X(net229));
 sky130_fd_sc_hd__and2_2 c233 (.A(net229),
    .B(net228),
    .X(net230));
 sky130_fd_sc_hd__and3_1 c234 (.A(net230),
    .B(net229),
    .C(net1078),
    .X(net231));
 sky130_fd_sc_hd__buf_1 c235 (.A(net776),
    .X(net232));
 sky130_fd_sc_hd__sdfxtp_1 c236 (.CLK(clknet_leaf_23_clk),
    .D(net231),
    .SCD(net232),
    .SCE(net1078),
    .Q(net233));
 sky130_fd_sc_hd__and3_1 c237 (.A(net233),
    .B(net230),
    .C(net1078),
    .X(net234));
 sky130_fd_sc_hd__a2111o_1 c238 (.A1(net232),
    .A2(net233),
    .B1(net230),
    .C1(net1078),
    .D1(net229),
    .X(net235));
 sky130_fd_sc_hd__dfbbn_1 c239 (.CLK_N(clknet_leaf_23_clk),
    .D(net234),
    .RESET_B(net229),
    .SET_B(net233),
    .Q(net237),
    .Q_N(net236));
 sky130_fd_sc_hd__or4bb_4 c240 (.A(net1078),
    .B(net233),
    .C_N(net236),
    .D_N(net887),
    .X(net1058));
 sky130_fd_sc_hd__dfbbn_1 c241 (.CLK_N(clknet_leaf_22_clk),
    .D(net231),
    .RESET_B(net230),
    .SET_B(net232),
    .Q(net239),
    .Q_N(net238));
 sky130_fd_sc_hd__a2111o_1 c242 (.A1(net239),
    .A2(net229),
    .B1(net1078),
    .C1(net1058),
    .D1(net233),
    .X(net240));
 sky130_fd_sc_hd__sdfbbp_1 c243 (.CLK(clknet_leaf_22_clk),
    .D(net240),
    .RESET_B(net235),
    .SCD(net230),
    .SCE(net238),
    .SET_B(net1078),
    .Q(net241));
 sky130_fd_sc_hd__and3_1 c244 (.A(net229),
    .B(net230),
    .C(net232),
    .X(net242));
 sky130_fd_sc_hd__sedfxtp_1 c245 (.CLK(clknet_leaf_22_clk),
    .D(net242),
    .DE(net239),
    .SCD(net231),
    .SCE(net232),
    .Q(net243));
 sky130_fd_sc_hd__sedfxtp_1 c246 (.CLK(clknet_leaf_23_clk),
    .D(net243),
    .DE(net242),
    .SCD(net237),
    .SCE(net1147),
    .Q(net244));
 sky130_fd_sc_hd__buf_1 c247 (.A(net847),
    .X(net245));
 sky130_fd_sc_hd__mux4_1 c248 (.A0(net245),
    .A1(net243),
    .A2(net235),
    .A3(net242),
    .S0(net1078),
    .S1(net229),
    .X(net246));
 sky130_fd_sc_hd__mux4_1 c249 (.A0(net244),
    .A1(net241),
    .A2(net1078),
    .A3(net243),
    .S0(net245),
    .S1(net229),
    .X(net247));
 sky130_fd_sc_hd__and2_0 c25 (.A(net1044),
    .B(net8),
    .X(net0));
 sky130_fd_sc_hd__mux4_1 c250 (.A0(net247),
    .A1(net1058),
    .A2(net245),
    .A3(net229),
    .S0(net228),
    .S1(net905),
    .X(net248));
 sky130_fd_sc_hd__mux4_1 c251 (.A0(net237),
    .A1(net248),
    .A2(net1058),
    .A3(net242),
    .S0(net230),
    .S1(net1185),
    .X(net249));
 sky130_fd_sc_hd__clkbuf_2 c252 (.A(in19),
    .X(net250));
 sky130_fd_sc_hd__and2_1 c253 (.A(net1042),
    .B(net250),
    .X(net251));
 sky130_fd_sc_hd__and2_0 c254 (.A(net251),
    .B(net250),
    .X(net252));
 sky130_fd_sc_hd__and2_1 c255 (.A(net250),
    .B(net251),
    .X(net253));
 sky130_fd_sc_hd__clkbuf_1 c256 (.A(net815),
    .X(net254));
 sky130_fd_sc_hd__buf_1 c257 (.A(net814),
    .X(net255));
 sky130_fd_sc_hd__and2_2 c258 (.A(net254),
    .B(net250),
    .X(net256));
 sky130_fd_sc_hd__dfbbp_1 c259 (.CLK(clknet_leaf_1_clk),
    .D(net252),
    .RESET_B(net254),
    .SET_B(net256),
    .Q(net258),
    .Q_N(net257));
 sky130_fd_sc_hd__and3_1 c26 (.A(net1045),
    .B(net804),
    .C(net8),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 c260 (.A(net1101),
    .X(net259));
 sky130_fd_sc_hd__and3_1 c261 (.A(net255),
    .B(net259),
    .C(net256),
    .X(net260));
 sky130_fd_sc_hd__buf_1 c262 (.A(net837),
    .X(net261));
 sky130_fd_sc_hd__a2111o_1 c263 (.A1(net136),
    .A2(net255),
    .B1(net261),
    .C1(net251),
    .D1(net250),
    .X(net262));
 sky130_fd_sc_hd__dlymetal6s2s_1 c264 (.A(net1021),
    .X(net263));
 sky130_fd_sc_hd__a2111o_1 c265 (.A1(net259),
    .A2(net263),
    .B1(net251),
    .C1(net255),
    .D1(net250),
    .X(net264));
 sky130_fd_sc_hd__mux4_1 c266 (.A0(net264),
    .A1(net261),
    .A2(clknet_1_0__leaf_net262),
    .A3(net251),
    .S0(net253),
    .S1(net250),
    .X(net265));
 sky130_fd_sc_hd__and2_0 c267 (.A(net263),
    .B(net907),
    .X(net266));
 sky130_fd_sc_hd__mux4_1 c268 (.A0(net250),
    .A1(net254),
    .A2(net261),
    .A3(net256),
    .S0(net263),
    .S1(net255),
    .X(net267));
 sky130_fd_sc_hd__sedfxtp_1 c269 (.CLK(clknet_leaf_2_clk),
    .D(net253),
    .DE(net263),
    .SCD(clknet_1_0__leaf_net262),
    .SCE(net1151),
    .Q(net268));
 sky130_fd_sc_hd__and3_1 c27 (.A(net1),
    .B(net1044),
    .C(net1046),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 c270 (.A(net825),
    .X(net269));
 sky130_fd_sc_hd__mux4_1 c271 (.A0(net261),
    .A1(net269),
    .A2(net263),
    .A3(net255),
    .S0(net250),
    .S1(net258),
    .X(net270));
 sky130_fd_sc_hd__or4bb_1 c272 (.A(net266),
    .B(net270),
    .C_N(net269),
    .D_N(net256),
    .X(net271));
 sky130_fd_sc_hd__buf_1 c273 (.A(net893),
    .X(net272));
 sky130_fd_sc_hd__and2_2 c274 (.A(net272),
    .B(net892),
    .X(net273));
 sky130_fd_sc_hd__and3_1 c275 (.A(net272),
    .B(net273),
    .C(net892),
    .X(net274));
 sky130_fd_sc_hd__clkbuf_2 c276 (.A(net796),
    .X(net275));
 sky130_fd_sc_hd__and2_0 c277 (.A(net275),
    .B(net893),
    .X(net276));
 sky130_fd_sc_hd__and2_1 c278 (.A(net276),
    .B(net275),
    .X(net277));
 sky130_fd_sc_hd__sdfrbp_1 c279 (.CLK(clknet_leaf_7_clk),
    .D(net274),
    .RESET_B(net1093),
    .SCD(net273),
    .SCE(net893),
    .Q(net279),
    .Q_N(net278));
 sky130_fd_sc_hd__and3_1 c28 (.A(net792),
    .B(net801),
    .C(net1046),
    .X(net3));
 sky130_fd_sc_hd__and2_1 c280 (.A(net273),
    .B(net277),
    .X(net280));
 sky130_fd_sc_hd__or4bb_1 c281 (.A(net279),
    .B(net273),
    .C_N(net277),
    .D_N(net275),
    .X(net281));
 sky130_fd_sc_hd__sdfrbp_1 c282 (.CLK(clknet_leaf_5_clk),
    .D(net277),
    .RESET_B(net280),
    .SCD(net275),
    .SCE(net892),
    .Q(net283),
    .Q_N(net282));
 sky130_fd_sc_hd__buf_1 c283 (.A(net796),
    .X(net284));
 sky130_fd_sc_hd__clkbuf_1 c284 (.A(net825),
    .X(net285));
 sky130_fd_sc_hd__sdfrtn_1 c285 (.CLK_N(clknet_leaf_5_clk),
    .D(net283),
    .RESET_B(net275),
    .SCD(net280),
    .SCE(net273),
    .Q(net286));
 sky130_fd_sc_hd__and2_0 c286 (.A(net285),
    .B(net284),
    .X(net287));
 sky130_fd_sc_hd__or4bb_1 c287 (.A(net287),
    .B(net277),
    .C_N(net282),
    .D_N(net273),
    .X(net288));
 sky130_fd_sc_hd__and2_1 c288 (.A(net275),
    .B(net284),
    .X(net289));
 sky130_fd_sc_hd__sdfbbn_1 c289 (.CLK_N(clknet_leaf_5_clk),
    .D(net281),
    .RESET_B(net283),
    .SCD(net289),
    .SCE(net275),
    .SET_B(net1117),
    .Q(net291),
    .Q_N(net290));
 sky130_fd_sc_hd__and2_1 c29 (.A(net0),
    .B(net1039),
    .X(net4));
 sky130_fd_sc_hd__and3_1 c290 (.A(net1181),
    .B(net273),
    .C(net290),
    .X(net292));
 sky130_fd_sc_hd__sdfrtp_1 c291 (.CLK(clknet_leaf_5_clk),
    .D(net288),
    .RESET_B(net292),
    .SCD(net291),
    .SCE(net289),
    .Q(net293));
 sky130_fd_sc_hd__sdfbbn_1 c292 (.CLK_N(clknet_leaf_5_clk),
    .D(net1103),
    .RESET_B(net1118),
    .SCD(net287),
    .SCE(net288),
    .SET_B(net282),
    .Q(net295),
    .Q_N(net294));
 sky130_fd_sc_hd__a2111o_2 c293 (.A1(net284),
    .A2(net293),
    .B1(net294),
    .C1(net289),
    .D1(net290),
    .X(net296));
 sky130_fd_sc_hd__and2_1 c294 (.A(net295),
    .B(net180),
    .X(net297));
 sky130_fd_sc_hd__and2_1 c295 (.A(net297),
    .B(net180),
    .X(net298));
 sky130_fd_sc_hd__and2_2 c296 (.A(net297),
    .B(net298),
    .X(net299));
 sky130_fd_sc_hd__and2_1 c297 (.A(net298),
    .B(net297),
    .X(net300));
 sky130_fd_sc_hd__clkbuf_2 c298 (.A(net1094),
    .X(net301));
 sky130_fd_sc_hd__buf_1 c299 (.A(net779),
    .X(net302));
 sky130_fd_sc_hd__and3_1 c30 (.A(net1044),
    .B(net1052),
    .C(net3),
    .X(net5));
 sky130_fd_sc_hd__sdfxbp_1 c300 (.CLK(clknet_leaf_9_clk),
    .D(net301),
    .SCD(net299),
    .SCE(net300),
    .Q(net304),
    .Q_N(net303));
 sky130_fd_sc_hd__sdfxbp_1 c301 (.CLK(clknet_leaf_10_clk),
    .D(net302),
    .SCD(net300),
    .SCE(net1132),
    .Q(net306),
    .Q_N(net305));
 sky130_fd_sc_hd__sdfrtp_1 c302 (.CLK(clknet_leaf_9_clk),
    .D(net1132),
    .RESET_B(net301),
    .SCD(net299),
    .SCE(net305),
    .Q(net307));
 sky130_fd_sc_hd__and3_1 c303 (.A(net307),
    .B(net304),
    .C(net306),
    .X(net308));
 sky130_fd_sc_hd__mux4_1 c304 (.A0(net308),
    .A1(net300),
    .A2(net305),
    .A3(net303),
    .S0(net301),
    .S1(net299),
    .X(net309));
 sky130_fd_sc_hd__sdfrtp_1 c305 (.CLK(clknet_leaf_10_clk),
    .D(net1125),
    .RESET_B(net299),
    .SCD(net301),
    .SCE(net303),
    .Q(net310));
 sky130_fd_sc_hd__sdfxtp_1 c306 (.CLK(clknet_leaf_6_clk),
    .D(net300),
    .SCD(net1114),
    .SCE(net1158),
    .Q(net311));
 sky130_fd_sc_hd__and3_1 c307 (.A(net310),
    .B(net298),
    .C(net908),
    .X(net312));
 sky130_fd_sc_hd__buf_1 c308 (.A(clknet_1_1__leaf_net1027),
    .X(net313));
 sky130_fd_sc_hd__mux4_1 c309 (.A0(net311),
    .A1(net298),
    .A2(net312),
    .A3(net306),
    .S0(net301),
    .S1(clknet_1_0__leaf_net313),
    .X(net314));
 sky130_fd_sc_hd__dlymetal6s2s_1 c31 (.X(net6));
 sky130_fd_sc_hd__sdfbbp_1 c310 (.CLK(clknet_leaf_6_clk),
    .D(net312),
    .RESET_B(net311),
    .SCD(clknet_1_0__leaf_net313),
    .SCE(net1158),
    .SET_B(clknet_1_0__leaf_net909),
    .Q(net316),
    .Q_N(net315));
 sky130_fd_sc_hd__mux4_1 c311 (.A0(net312),
    .A1(net315),
    .A2(clknet_1_0__leaf_net313),
    .A3(net299),
    .S0(net302),
    .S1(clknet_1_0__leaf_net909),
    .X(net317));
 sky130_fd_sc_hd__sdfbbn_1 c312 (.CLK_N(clknet_leaf_6_clk),
    .D(net316),
    .RESET_B(clknet_1_1__leaf_net313),
    .SCD(net299),
    .SCE(clknet_1_0__leaf_net909),
    .SET_B(clknet_1_0__leaf_net910),
    .Q(net319),
    .Q_N(net318));
 sky130_fd_sc_hd__mux4_1 c313 (.A0(clknet_1_1__leaf_net313),
    .A1(net312),
    .A2(net318),
    .A3(net908),
    .S0(clknet_1_1__leaf_net909),
    .S1(clknet_1_1__leaf_net910),
    .X(net320));
 sky130_fd_sc_hd__sdfbbn_1 c314 (.CLK_N(clknet_leaf_15_clk),
    .D(net1126),
    .RESET_B(clknet_1_1__leaf_net313),
    .SCD(net299),
    .SCE(clknet_1_1__leaf_net909),
    .SET_B(clknet_1_0__leaf_net911),
    .Q(net322),
    .Q_N(net321));
 sky130_fd_sc_hd__and2_1 c315 (.A(net296),
    .B(net180),
    .X(net323));
 sky130_fd_sc_hd__buf_1 c316 (.A(net789),
    .X(net324));
 sky130_fd_sc_hd__buf_1 c317 (.A(net789),
    .X(net325));
 sky130_fd_sc_hd__clkbuf_1 c318 (.A(net1015),
    .X(net326));
 sky130_fd_sc_hd__clkbuf_2 c319 (.A(net821),
    .X(net327));
 sky130_fd_sc_hd__clkbuf_1 c32 (.A(net803),
    .X(net7));
 sky130_fd_sc_hd__and2_1 c320 (.A(net326),
    .B(net327),
    .X(net328));
 sky130_fd_sc_hd__and3_1 c321 (.A(net325),
    .B(net1073),
    .C(net327),
    .X(net329));
 sky130_fd_sc_hd__and2_1 c322 (.A(net329),
    .B(net324),
    .X(net330));
 sky130_fd_sc_hd__buf_1 c323 (.A(net1015),
    .X(net331));
 sky130_fd_sc_hd__buf_2 c324 (.A(net1023),
    .X(net332));
 sky130_fd_sc_hd__sdfbbp_1 c325 (.CLK(clknet_leaf_16_clk),
    .D(net1073),
    .RESET_B(net326),
    .SCD(net329),
    .SCE(net330),
    .SET_B(net1172),
    .Q(net334),
    .Q_N(net333));
 sky130_fd_sc_hd__sdfbbn_1 c326 (.CLK_N(clknet_leaf_16_clk),
    .D(net1160),
    .RESET_B(net1073),
    .SCD(net332),
    .SCE(net330),
    .SET_B(net324),
    .Q(net336),
    .Q_N(net335));
 sky130_fd_sc_hd__mux4_1 c327 (.A0(net334),
    .A1(net336),
    .A2(net322),
    .A3(net332),
    .S0(net327),
    .S1(net1073),
    .X(net337));
 sky130_fd_sc_hd__mux4_2 c328 (.A0(net297),
    .A1(net334),
    .A2(net335),
    .A3(net327),
    .S0(net331),
    .S1(net1073),
    .X(net338));
 sky130_fd_sc_hd__mux4_1 c329 (.A0(net337),
    .A1(net330),
    .A2(net338),
    .A3(net332),
    .S0(net329),
    .S1(net1073),
    .X(net339));
 sky130_fd_sc_hd__and2_2 c33 (.A(net1041),
    .B(net1036),
    .X(net8));
 sky130_fd_sc_hd__mux4_1 c330 (.A0(net323),
    .A1(net336),
    .A2(net338),
    .A3(net324),
    .S0(net328),
    .S1(net912),
    .X(net340));
 sky130_fd_sc_hd__or4bb_1 c331 (.A(net325),
    .B(net1073),
    .C_N(net338),
    .D_N(net329),
    .X(net341));
 sky130_fd_sc_hd__sdfbbn_1 c332 (.CLK_N(clknet_leaf_16_clk),
    .D(net1177),
    .RESET_B(net341),
    .SCD(net332),
    .SCE(net1073),
    .SET_B(net184),
    .Q(net343),
    .Q_N(net342));
 sky130_fd_sc_hd__mux4_1 c333 (.A0(net338),
    .A1(net343),
    .A2(net337),
    .A3(net1073),
    .S0(net327),
    .S1(net341),
    .X(net344));
 sky130_fd_sc_hd__mux4_1 c334 (.A0(net341),
    .A1(net338),
    .A2(net328),
    .A3(net333),
    .S0(net915),
    .S1(net917),
    .X(net345));
 sky130_fd_sc_hd__mux4_1 c335 (.A0(net342),
    .A1(net341),
    .A2(net328),
    .A3(net913),
    .S0(net916),
    .S1(net918),
    .X(net346));
 sky130_fd_sc_hd__buf_1 c336 (.A(net813),
    .X(net347));
 sky130_fd_sc_hd__and2_1 c337 (.A(net226),
    .B(net915),
    .X(net348));
 sky130_fd_sc_hd__and2_2 c338 (.A(net348),
    .B(net226),
    .X(net349));
 sky130_fd_sc_hd__and3_2 c339 (.A(net332),
    .B(net349),
    .C(net348),
    .X(net350));
 sky130_fd_sc_hd__and2_1 c34 (.A(net1046),
    .B(net1040),
    .X(net9));
 sky130_fd_sc_hd__sdfsbp_1 c340 (.CLK(clknet_leaf_29_clk),
    .D(net348),
    .SCD(net347),
    .SCE(net350),
    .SET_B(net915),
    .Q(net352),
    .Q_N(net351));
 sky130_fd_sc_hd__and3_1 c341 (.A(net348),
    .B(net352),
    .C(net919),
    .X(net353));
 sky130_fd_sc_hd__buf_1 c342 (.A(net812),
    .X(net354));
 sky130_fd_sc_hd__clkbuf_2 c343 (.A(net857),
    .X(net355));
 sky130_fd_sc_hd__a2111o_1 c344 (.A1(net347),
    .A2(net355),
    .B1(net354),
    .C1(net351),
    .D1(net1096),
    .X(net356));
 sky130_fd_sc_hd__and3_1 c345 (.A(net349),
    .B(net1187),
    .C(net355),
    .X(net357));
 sky130_fd_sc_hd__buf_1 c346 (.A(net856),
    .X(net358));
 sky130_fd_sc_hd__sdfbbp_1 c347 (.CLK(clknet_leaf_18_clk),
    .D(net354),
    .RESET_B(net355),
    .SCD(net350),
    .SCE(net349),
    .SET_B(net1105),
    .Q(net360),
    .Q_N(net359));
 sky130_fd_sc_hd__sdfbbn_1 c348 (.CLK_N(clknet_leaf_18_clk),
    .D(net348),
    .RESET_B(net1188),
    .SCD(net357),
    .SCE(net359),
    .SET_B(net354),
    .Q(net361));
 sky130_fd_sc_hd__sdfbbn_1 c349 (.CLK_N(clknet_leaf_19_clk),
    .D(net222),
    .RESET_B(net360),
    .SCD(net227),
    .SCE(net349),
    .SET_B(net350),
    .Q(net363),
    .Q_N(net362));
 sky130_fd_sc_hd__mux4_1 c35 (.A0(net2),
    .A1(net5),
    .A2(net1038),
    .A3(net1080),
    .S0(net4),
    .S1(net6),
    .X(net10));
 sky130_fd_sc_hd__mux4_1 c350 (.A0(net357),
    .A1(net355),
    .A2(net350),
    .A3(net354),
    .S0(net349),
    .S1(net351),
    .X(net364));
 sky130_fd_sc_hd__a2111o_1 c351 (.A1(net360),
    .A2(net347),
    .B1(net358),
    .C1(net355),
    .D1(net352),
    .X(net365));
 sky130_fd_sc_hd__sdfbbp_1 c352 (.CLK(clknet_leaf_19_clk),
    .D(net361),
    .RESET_B(net365),
    .SCD(net350),
    .SCE(net362),
    .SET_B(net357),
    .Q(net367),
    .Q_N(net366));
 sky130_fd_sc_hd__mux4_2 c353 (.A0(net352),
    .A1(net358),
    .A2(net355),
    .A3(net365),
    .S0(net353),
    .S1(net366),
    .X(net368));
 sky130_fd_sc_hd__mux4_1 c354 (.A0(net353),
    .A1(net363),
    .A2(net367),
    .A3(net368),
    .S0(net332),
    .S1(net355),
    .X(net369));
 sky130_fd_sc_hd__sdfbbn_1 c355 (.CLK_N(clknet_leaf_28_clk),
    .D(net367),
    .RESET_B(net368),
    .SCD(net355),
    .SCE(net1163),
    .SET_B(net921),
    .Q(net370));
 sky130_fd_sc_hd__mux4_1 c356 (.A0(net365),
    .A1(net370),
    .A2(net353),
    .A3(net366),
    .S0(net368),
    .S1(net921),
    .X(net371));
 sky130_fd_sc_hd__and2_1 c357 (.A(net886),
    .B(net906),
    .X(net372));
 sky130_fd_sc_hd__and3_1 c358 (.A(net372),
    .B(net225),
    .C(net906),
    .X(net373));
 sky130_fd_sc_hd__and2_2 c359 (.A(net1058),
    .B(net906),
    .X(net374));
 sky130_fd_sc_hd__sdfbbn_1 c36 (.CLK_N(clknet_leaf_9_clk),
    .D(net5),
    .RESET_B(net4),
    .SCD(net3),
    .SCE(net6),
    .SET_B(net1080),
    .Q(net12),
    .Q_N(net11));
 sky130_fd_sc_hd__and2_1 c360 (.A(net1112),
    .B(net922),
    .X(net375));
 sky130_fd_sc_hd__buf_1 c361 (.A(clknet_1_0__leaf_net1007),
    .X(net376));
 sky130_fd_sc_hd__and2_0 c362 (.A(net374),
    .B(clknet_1_0__leaf_net376),
    .X(net377));
 sky130_fd_sc_hd__and3_1 c363 (.A(net375),
    .B(net372),
    .C(net905),
    .X(net378));
 sky130_fd_sc_hd__buf_1 c364 (.A(clknet_1_1__leaf_net1007),
    .X(net379));
 sky130_fd_sc_hd__clkbuf_1 c365 (.X(net861));
 sky130_fd_sc_hd__clkbuf_2 c366 (.A(net861),
    .X(net381));
 sky130_fd_sc_hd__sdfbbn_1 c367 (.CLK_N(clknet_leaf_28_clk),
    .D(net380),
    .RESET_B(net375),
    .SCD(net374),
    .SCE(clknet_1_0__leaf_net377),
    .SET_B(net368),
    .Q(net383),
    .Q_N(net382));
 sky130_fd_sc_hd__sdfbbp_1 c368 (.CLK(clknet_leaf_25_clk),
    .D(net383),
    .RESET_B(net368),
    .SCD(net372),
    .SCE(net380),
    .SET_B(net1097),
    .Q(net385),
    .Q_N(net384));
 sky130_fd_sc_hd__sdfbbn_1 c369 (.CLK_N(clknet_leaf_25_clk),
    .D(net374),
    .RESET_B(net381),
    .SCD(clknet_1_1__leaf_net376),
    .SCE(clknet_1_1__leaf_net377),
    .SET_B(net380),
    .Q(net387),
    .Q_N(net386));
 sky130_fd_sc_hd__mux4_1 c37 (.A0(net7),
    .A1(net2),
    .A2(net6),
    .A3(net8),
    .S0(net11),
    .S1(net1142),
    .X(net13));
 sky130_fd_sc_hd__mux4_2 c370 (.A0(net387),
    .A1(net385),
    .A2(net381),
    .A3(net380),
    .S0(net374),
    .S1(net906),
    .X(net388));
 sky130_fd_sc_hd__mux4_1 c371 (.A0(net378),
    .A1(net388),
    .A2(net383),
    .A3(net380),
    .S0(net381),
    .S1(clknet_1_1__leaf_net379),
    .X(net389));
 sky130_fd_sc_hd__sdfbbn_1 c372 (.CLK_N(clknet_leaf_25_clk),
    .D(net1143),
    .RESET_B(net1133),
    .SCD(net388),
    .SCE(net384),
    .SET_B(net924),
    .Q(net391),
    .Q_N(net390));
 sky130_fd_sc_hd__mux4_1 c373 (.A0(net385),
    .A1(net388),
    .A2(net391),
    .A3(net386),
    .S0(net1058),
    .S1(net1180),
    .X(net392));
 sky130_fd_sc_hd__mux4_1 c374 (.A0(clknet_1_0__leaf_net379),
    .A1(net391),
    .A2(clknet_1_1__leaf_net377),
    .A3(net382),
    .S0(net374),
    .S1(net381),
    .X(net393));
 sky130_fd_sc_hd__mux4_1 c375 (.A0(net388),
    .A1(net374),
    .A2(net384),
    .A3(net390),
    .S0(net924),
    .S1(net1144),
    .X(net394));
 sky130_fd_sc_hd__mux4_1 c376 (.A0(net391),
    .A1(net382),
    .A2(net388),
    .A3(net923),
    .S0(net1176),
    .S1(net927),
    .X(net395));
 sky130_fd_sc_hd__mux4_1 c377 (.A0(net372),
    .A1(net387),
    .A2(net390),
    .A3(net924),
    .S0(net927),
    .S1(net928),
    .X(net396));
 sky130_fd_sc_hd__clkbuf_2 c378 (.A(net1098),
    .X(net397));
 sky130_fd_sc_hd__dlymetal6s2s_1 c379 (.A(net1098),
    .X(net398));
 sky130_fd_sc_hd__sdfbbn_1 c38 (.CLK_N(clknet_leaf_9_clk),
    .D(net1123),
    .RESET_B(net1080),
    .SCD(net4),
    .SCE(net1046),
    .SET_B(net867),
    .Q(net14));
 sky130_fd_sc_hd__sdfxtp_1 c380 (.CLK(clknet_leaf_42_clk),
    .D(net271),
    .SCD(net398),
    .SCE(net397),
    .Q(net399));
 sky130_fd_sc_hd__and2_1 c381 (.A(net1083),
    .B(net398),
    .X(net400));
 sky130_fd_sc_hd__and2_1 c382 (.A(net400),
    .B(net399),
    .X(net401));
 sky130_fd_sc_hd__and2_0 c383 (.A(net401),
    .B(net397),
    .X(net402));
 sky130_fd_sc_hd__clkbuf_1 c384 (.A(net859),
    .X(net403));
 sky130_fd_sc_hd__sdfbbp_1 c385 (.CLK(clknet_leaf_0_clk),
    .D(net400),
    .RESET_B(net1116),
    .SCD(net1083),
    .SCE(net1067),
    .SET_B(net398),
    .Q(net405),
    .Q_N(net404));
 sky130_fd_sc_hd__clkbuf_1 c386 (.A(net826),
    .X(net406));
 sky130_fd_sc_hd__buf_1 c387 (.A(net858),
    .X(net407));
 sky130_fd_sc_hd__and3_1 c388 (.A(net403),
    .B(net400),
    .C(net407),
    .X(net408));
 sky130_fd_sc_hd__sdfbbn_1 c389 (.CLK_N(clknet_leaf_0_clk),
    .D(net406),
    .RESET_B(net400),
    .SCD(net408),
    .SCE(net399),
    .SET_B(net1067),
    .Q(net410),
    .Q_N(net409));
 sky130_fd_sc_hd__mux4_1 c39 (.A0(net6),
    .A1(net14),
    .A2(net3),
    .A3(net1044),
    .S0(net4),
    .S1(net866),
    .X(net15));
 sky130_fd_sc_hd__or4bb_1 c390 (.A(net410),
    .B(net1083),
    .C_N(net408),
    .D_N(net398),
    .X(net411));
 sky130_fd_sc_hd__sdfbbn_1 c391 (.CLK_N(clknet_leaf_0_clk),
    .D(net1067),
    .RESET_B(net1084),
    .SCD(net1159),
    .SCE(net397),
    .SET_B(net398),
    .Q(net412));
 sky130_fd_sc_hd__mux4_1 c392 (.A0(net398),
    .A1(net410),
    .A2(net411),
    .A3(net1067),
    .S0(net397),
    .S1(net404),
    .X(net413));
 sky130_fd_sc_hd__buf_1 c393 (.A(net836),
    .X(net414));
 sky130_fd_sc_hd__sdfbbp_1 c394 (.CLK(clknet_leaf_0_clk),
    .D(net412),
    .RESET_B(net1084),
    .SCD(net402),
    .SCE(net405),
    .SET_B(clknet_1_0__leaf_net929),
    .Q(net416),
    .Q_N(net415));
 sky130_fd_sc_hd__sdfbbn_1 c395 (.CLK_N(clknet_leaf_0_clk),
    .D(net414),
    .RESET_B(net416),
    .SCD(net1067),
    .SCE(net404),
    .SET_B(clknet_1_0__leaf_net929),
    .Q(net418),
    .Q_N(net417));
 sky130_fd_sc_hd__mux4_1 c396 (.A0(net408),
    .A1(net416),
    .A2(net418),
    .A3(net399),
    .S0(net401),
    .S1(net1067),
    .X(net419));
 sky130_fd_sc_hd__mux4_1 c397 (.A0(net397),
    .A1(net414),
    .A2(net415),
    .A3(net417),
    .S0(net407),
    .S1(clknet_1_0__leaf_net930),
    .X(net420));
 sky130_fd_sc_hd__mux4_1 c398 (.A0(net418),
    .A1(net420),
    .A2(net415),
    .A3(net1067),
    .S0(clknet_1_1__leaf_net929),
    .S1(clknet_1_1__leaf_net930),
    .X(net421));
 sky130_fd_sc_hd__and2_2 c399 (.A(net272),
    .B(net405),
    .X(net422));
 sky130_fd_sc_hd__mux4_1 c40 (.A0(net3),
    .A1(net6),
    .A2(net8),
    .A3(net1),
    .S0(net867),
    .S1(net868),
    .X(net16));
 sky130_fd_sc_hd__and2_1 c400 (.A(net422),
    .B(net405),
    .X(net423));
 sky130_fd_sc_hd__clkbuf_2 c401 (.A(net790),
    .X(net424));
 sky130_fd_sc_hd__buf_2 c402 (.A(net790),
    .X(net425));
 sky130_fd_sc_hd__sdfsbp_1 c403 (.CLK(clknet_leaf_2_clk),
    .D(net424),
    .SCD(net422),
    .SCE(net1069),
    .SET_B(net425),
    .Q(net427),
    .Q_N(net426));
 sky130_fd_sc_hd__and2_1 c404 (.A(net425),
    .B(net426),
    .X(net428));
 sky130_fd_sc_hd__and2_1 c405 (.A(net424),
    .B(net425),
    .X(net429));
 sky130_fd_sc_hd__and3_2 c406 (.A(net427),
    .B(net424),
    .C(net422),
    .X(net430));
 sky130_fd_sc_hd__sdfbbn_1 c407 (.CLK_N(clknet_leaf_2_clk),
    .D(net422),
    .RESET_B(net428),
    .SCD(net1069),
    .SCE(net425),
    .SET_B(net404),
    .Q(net432),
    .Q_N(net431));
 sky130_fd_sc_hd__sdfbbp_1 c408 (.CLK(clknet_leaf_3_clk),
    .D(net429),
    .RESET_B(net431),
    .SCD(net428),
    .SCE(net430),
    .SET_B(net1069),
    .Q(net434),
    .Q_N(net433));
 sky130_fd_sc_hd__and3_1 c409 (.A(net428),
    .B(net424),
    .C(net422),
    .X(net435));
 sky130_fd_sc_hd__mux4_1 c41 (.A0(net16),
    .A1(net6),
    .A2(net1080),
    .A3(net1046),
    .S0(net866),
    .S1(net1149),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 c410 (.A(net1022),
    .X(net436));
 sky130_fd_sc_hd__sdfbbn_1 c411 (.CLK_N(clknet_leaf_3_clk),
    .D(net1131),
    .RESET_B(net296),
    .SCD(net425),
    .SCE(net424),
    .SET_B(net1069),
    .Q(net438),
    .Q_N(net437));
 sky130_fd_sc_hd__sdfxtp_1 c412 (.CLK(clknet_leaf_3_clk),
    .D(net435),
    .SCD(net430),
    .SCE(net425),
    .Q(net439));
 sky130_fd_sc_hd__dfbbn_1 c413 (.CLK_N(clknet_leaf_4_clk),
    .D(net436),
    .RESET_B(net439),
    .SET_B(net430),
    .Q(net441),
    .Q_N(net440));
 sky130_fd_sc_hd__a2111o_4 c414 (.A1(net425),
    .A2(net437),
    .B1(net429),
    .C1(net424),
    .D1(net428),
    .X(net442));
 sky130_fd_sc_hd__mux4_1 c415 (.A0(net434),
    .A1(net429),
    .A2(net442),
    .A3(net422),
    .S0(net424),
    .S1(net430),
    .X(net443));
 sky130_fd_sc_hd__dfbbn_1 c416 (.CLK_N(clknet_leaf_3_clk),
    .D(net280),
    .RESET_B(net425),
    .SET_B(net1115),
    .Q(net445),
    .Q_N(net444));
 sky130_fd_sc_hd__mux4_1 c417 (.A0(net445),
    .A1(net438),
    .A2(net442),
    .A3(net430),
    .S0(net422),
    .S1(net933),
    .X(net446));
 sky130_fd_sc_hd__mux4_1 c418 (.A0(net438),
    .A1(net439),
    .A2(net445),
    .A3(net430),
    .S0(net442),
    .S1(net1182),
    .X(net447));
 sky130_fd_sc_hd__mux4_1 c419 (.A0(net430),
    .A1(net432),
    .A2(net444),
    .A3(net422),
    .S0(net934),
    .S1(net935),
    .X(net448));
 sky130_fd_sc_hd__and2_1 c42 (.A(net1080),
    .B(net1109),
    .X(net18));
 sky130_fd_sc_hd__and2_1 c420 (.A(net322),
    .B(net936),
    .X(net449));
 sky130_fd_sc_hd__and2_0 c421 (.A(net449),
    .B(clknet_1_1__leaf_net911),
    .X(net450));
 sky130_fd_sc_hd__and2_0 c422 (.A(clknet_1_0__leaf_net450),
    .B(net442),
    .X(net451));
 sky130_fd_sc_hd__dfbbp_1 c423 (.CLK(clknet_leaf_40_clk),
    .D(net441),
    .RESET_B(clknet_1_1__leaf_net451),
    .SET_B(net936),
    .Q(net452));
 sky130_fd_sc_hd__clkbuf_1 c424 (.A(net807),
    .X(net453));
 sky130_fd_sc_hd__and2_0 c425 (.A(net442),
    .B(clknet_1_0__leaf_net450),
    .X(net454));
 sky130_fd_sc_hd__buf_1 c426 (.A(net1025),
    .X(net455));
 sky130_fd_sc_hd__and2_1 c427 (.A(net453),
    .B(net322),
    .X(net456));
 sky130_fd_sc_hd__and3_1 c428 (.A(net449),
    .B(net1068),
    .C(net453),
    .X(net457));
 sky130_fd_sc_hd__and2_0 c429 (.A(net457),
    .B(net449),
    .X(net458));
 sky130_fd_sc_hd__and2_1 c43 (.A(net18),
    .B(net1080),
    .X(net19));
 sky130_fd_sc_hd__buf_1 c430 (.A(net807),
    .X(net459));
 sky130_fd_sc_hd__and3_1 c431 (.A(net459),
    .B(net455),
    .C(net936),
    .X(net460));
 sky130_fd_sc_hd__and2_1 c432 (.A(net459),
    .B(net441),
    .X(net461));
 sky130_fd_sc_hd__or4bb_1 c433 (.A(clknet_1_1__leaf_net450),
    .B(net461),
    .C_N(net459),
    .D_N(net1068),
    .X(net462));
 sky130_fd_sc_hd__or4bb_1 c434 (.A(net455),
    .B(net1068),
    .C_N(net461),
    .D_N(net457),
    .X(net463));
 sky130_fd_sc_hd__mux4_1 c435 (.A0(net460),
    .A1(net461),
    .A2(clknet_1_1__leaf_net462),
    .A3(net459),
    .S0(net1068),
    .S1(net463),
    .X(net464));
 sky130_fd_sc_hd__sdfbbn_1 c436 (.CLK_N(clknet_leaf_4_clk),
    .D(clknet_1_0__leaf_net462),
    .RESET_B(net459),
    .SCD(net1068),
    .SCE(net455),
    .SET_B(net1119),
    .Q(net465));
 sky130_fd_sc_hd__mux4_1 c437 (.A0(net461),
    .A1(net465),
    .A2(clknet_1_1__leaf_net462),
    .A3(net460),
    .S0(net1068),
    .S1(net937),
    .X(net466));
 sky130_fd_sc_hd__mux4_1 c438 (.A0(net458),
    .A1(net440),
    .A2(net459),
    .A3(net463),
    .S0(net1068),
    .S1(net1134),
    .X(net467));
 sky130_fd_sc_hd__mux4_1 c439 (.A0(net463),
    .A1(net459),
    .A2(clknet_1_0__leaf_net462),
    .A3(clknet_1_1__leaf_net450),
    .S0(net455),
    .S1(net1119),
    .X(net468));
 sky130_fd_sc_hd__buf_1 c44 (.A(net808),
    .X(net20));
 sky130_fd_sc_hd__mux4_1 c440 (.A0(net463),
    .A1(clknet_1_0__leaf_net451),
    .A2(net936),
    .A3(net937),
    .S0(net939),
    .S1(net940),
    .X(net469));
 sky130_fd_sc_hd__buf_2 c441 (.X(net470));
 sky130_fd_sc_hd__and2_0 c442 (.A(net1079),
    .B(net941),
    .X(net471));
 sky130_fd_sc_hd__dlymetal6s2s_1 c443 (.A(net772),
    .X(net472));
 sky130_fd_sc_hd__and2_1 c444 (.A(net1079),
    .B(net472),
    .X(net473));
 sky130_fd_sc_hd__and2_1 c445 (.A(net1079),
    .B(net472),
    .X(net474));
 sky130_fd_sc_hd__and3_1 c446 (.A(net474),
    .B(net473),
    .C(net1079),
    .X(net475));
 sky130_fd_sc_hd__and2_1 c447 (.A(net475),
    .B(net1079),
    .X(net476));
 sky130_fd_sc_hd__sdfxbp_1 c448 (.CLK(clknet_leaf_30_clk),
    .D(net476),
    .SCD(net472),
    .SCE(net471),
    .Q(net478),
    .Q_N(net477));
 sky130_fd_sc_hd__and3_1 c449 (.A(net471),
    .B(net187),
    .C(net472),
    .X(net479));
 sky130_fd_sc_hd__clkbuf_1 c45 (.A(net808),
    .X(net21));
 sky130_fd_sc_hd__and2_0 c450 (.A(net472),
    .B(net1079),
    .X(net480));
 sky130_fd_sc_hd__sdfstp_1 c451 (.CLK(clknet_leaf_30_clk),
    .D(clknet_1_1__leaf_net454),
    .SCD(net479),
    .SCE(net476),
    .SET_B(net1079),
    .Q(net481));
 sky130_fd_sc_hd__and3_1 c452 (.A(net470),
    .B(net472),
    .C(net942),
    .X(net482));
 sky130_fd_sc_hd__buf_1 c453 (.A(net1031),
    .X(net483));
 sky130_fd_sc_hd__and3_1 c454 (.A(net479),
    .B(net474),
    .C(net483),
    .X(net484));
 sky130_fd_sc_hd__sdfxbp_1 c455 (.CLK(clknet_leaf_17_clk),
    .D(net483),
    .SCD(net1129),
    .SCE(net484),
    .Q(net486),
    .Q_N(net485));
 sky130_fd_sc_hd__mux4_1 c456 (.A0(net1153),
    .A1(net482),
    .A2(net483),
    .A3(net484),
    .S0(net1079),
    .S1(net479),
    .X(net487));
 sky130_fd_sc_hd__mux4_1 c457 (.A0(net484),
    .A1(net1169),
    .A2(net472),
    .A3(net483),
    .S0(net1079),
    .S1(net943),
    .X(net488));
 sky130_fd_sc_hd__mux4_1 c458 (.A0(net478),
    .A1(net482),
    .A2(net485),
    .A3(net483),
    .S0(net1079),
    .S1(net943),
    .X(net489));
 sky130_fd_sc_hd__mux4_1 c459 (.A0(net480),
    .A1(net483),
    .A2(net489),
    .A3(net486),
    .S0(net474),
    .S1(net470),
    .X(net490));
 sky130_fd_sc_hd__buf_1 c46 (.A(net827),
    .X(net22));
 sky130_fd_sc_hd__mux4_1 c460 (.A0(net479),
    .A1(net484),
    .A2(net490),
    .A3(net485),
    .S0(net489),
    .S1(net1135),
    .X(net491));
 sky130_fd_sc_hd__mux4_1 c461 (.A0(net490),
    .A1(net489),
    .A2(net473),
    .A3(net483),
    .S0(net1179),
    .S1(net946),
    .X(net492));
 sky130_fd_sc_hd__buf_1 c462 (.A(net774),
    .X(net493));
 sky130_fd_sc_hd__buf_1 c463 (.A(net774),
    .X(net494));
 sky130_fd_sc_hd__and2_0 c464 (.A(net494),
    .B(net946),
    .X(net495));
 sky130_fd_sc_hd__and2_1 c465 (.A(net493),
    .B(net494),
    .X(net496));
 sky130_fd_sc_hd__and2_1 c466 (.A(net496),
    .B(net495),
    .X(net497));
 sky130_fd_sc_hd__and3_1 c467 (.A(net497),
    .B(net494),
    .C(net496),
    .X(net498));
 sky130_fd_sc_hd__buf_1 c468 (.X(net852));
 sky130_fd_sc_hd__a2111o_1 c469 (.A1(net495),
    .A2(net497),
    .B1(net499),
    .C1(net922),
    .D1(net946),
    .X(net500));
 sky130_fd_sc_hd__clkbuf_1 c47 (.A(net829),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_1 c470 (.A(net851),
    .X(net501));
 sky130_fd_sc_hd__clkbuf_1 c471 (.A(net1029),
    .X(net502));
 sky130_fd_sc_hd__and3_1 c472 (.A(net502),
    .B(net496),
    .C(net494),
    .X(net503));
 sky130_fd_sc_hd__sdfxtp_1 c473 (.CLK(clknet_leaf_29_clk),
    .D(net495),
    .SCD(net500),
    .SCE(net496),
    .Q(net504));
 sky130_fd_sc_hd__and3_1 c474 (.A(net493),
    .B(net502),
    .C(net494),
    .X(net505));
 sky130_fd_sc_hd__and3_1 c475 (.A(net499),
    .B(net503),
    .C(net505),
    .X(net506));
 sky130_fd_sc_hd__sdfbbp_1 c476 (.CLK(clknet_leaf_29_clk),
    .D(net498),
    .RESET_B(net505),
    .SCD(net506),
    .SCE(net499),
    .SET_B(net1095),
    .Q(net508),
    .Q_N(net507));
 sky130_fd_sc_hd__and2_0 c477 (.A(net505),
    .B(net501),
    .X(net509));
 sky130_fd_sc_hd__sdfbbn_1 c478 (.CLK_N(clknet_leaf_29_clk),
    .D(net504),
    .RESET_B(net493),
    .SCD(net506),
    .SCE(net499),
    .SET_B(net1186),
    .Q(net511),
    .Q_N(net510));
 sky130_fd_sc_hd__sdfbbn_1 c479 (.CLK_N(clknet_leaf_29_clk),
    .D(net503),
    .RESET_B(net504),
    .SCD(net506),
    .SCE(net510),
    .SET_B(net499),
    .Q(net513),
    .Q_N(net512));
 sky130_fd_sc_hd__and2_2 c48 (.A(net23),
    .B(net22),
    .X(net24));
 sky130_fd_sc_hd__sdfbbp_1 c480 (.CLK(clknet_leaf_28_clk),
    .D(net500),
    .RESET_B(net499),
    .SCD(net511),
    .SCE(net512),
    .SET_B(net506),
    .Q(net515),
    .Q_N(net514));
 sky130_fd_sc_hd__mux4_1 c481 (.A0(net511),
    .A1(net506),
    .A2(net513),
    .A3(net497),
    .S0(net514),
    .S1(net499),
    .X(net516));
 sky130_fd_sc_hd__mux4_1 c482 (.A0(net513),
    .A1(net515),
    .A2(net507),
    .A3(net506),
    .S0(net499),
    .S1(clknet_1_1__leaf_net948),
    .X(net517));
 sky130_fd_sc_hd__and2_0 c483 (.A(net509),
    .B(clknet_1_0__leaf_net948),
    .X(net518));
 sky130_fd_sc_hd__clkbuf_1 c484 (.A(net811),
    .X(net519));
 sky130_fd_sc_hd__sdfxtp_1 c485 (.CLK(clknet_leaf_27_clk),
    .D(net519),
    .SCD(net509),
    .SCE(clknet_1_0__leaf_net518),
    .Q(net1064));
 sky130_fd_sc_hd__buf_8 c486 (.A(net811),
    .X(net1059));
 sky130_fd_sc_hd__and3_1 c487 (.A(net1064),
    .B(net1072),
    .C(net949),
    .X(net520));
 sky130_fd_sc_hd__sdfbbn_1 c488 (.CLK_N(clknet_leaf_28_clk),
    .D(net381),
    .RESET_B(net519),
    .SCD(net1064),
    .SCE(net1081),
    .SET_B(clknet_1_0__leaf_net518),
    .Q(net522),
    .Q_N(net521));
 sky130_fd_sc_hd__and3_1 c489 (.A(clknet_1_0__leaf_net520),
    .B(net522),
    .C(net1072),
    .X(net523));
 sky130_fd_sc_hd__and2_1 c49 (.A(net22),
    .B(net21),
    .X(net25));
 sky130_fd_sc_hd__sdfxtp_1 c490 (.CLK(clknet_leaf_27_clk),
    .D(clknet_1_1__leaf_net518),
    .SCD(net1081),
    .SCE(net521),
    .Q(net524));
 sky130_fd_sc_hd__mux4_1 c491 (.A0(net519),
    .A1(clknet_1_1__leaf_net523),
    .A2(clknet_1_1__leaf_net518),
    .A3(net1072),
    .S0(net521),
    .S1(net927),
    .X(net525));
 sky130_fd_sc_hd__a2111o_1 c492 (.A1(clknet_1_0__leaf_net523),
    .A2(net1064),
    .B1(net524),
    .C1(net521),
    .D1(clknet_1_0__leaf_net950),
    .X(net526));
 sky130_fd_sc_hd__sdfstp_1 c493 (.CLK(clknet_leaf_27_clk),
    .D(net522),
    .SCD(net1081),
    .SCE(clknet_1_0__leaf_net526),
    .SET_B(net1089),
    .Q(net527));
 sky130_fd_sc_hd__sdfbbn_1 c494 (.CLK_N(clknet_leaf_26_clk),
    .D(clknet_1_0__leaf_net520),
    .RESET_B(net1064),
    .SCD(clknet_1_1__leaf_net518),
    .SCE(clknet_1_0__leaf_net526),
    .SET_B(clknet_1_0__leaf_net950),
    .Q(net529),
    .Q_N(net528));
 sky130_fd_sc_hd__sdfbbp_1 c495 (.CLK(clknet_leaf_27_clk),
    .D(clknet_1_1__leaf_net526),
    .RESET_B(net521),
    .SCD(net528),
    .SCE(net1157),
    .SET_B(clknet_1_0__leaf_net950),
    .Q(net531),
    .Q_N(net530));
 sky130_fd_sc_hd__mux4_1 c496 (.A0(clknet_1_0__leaf_net523),
    .A1(clknet_1_0__leaf_net526),
    .A2(net527),
    .A3(net522),
    .S0(net528),
    .S1(net1081),
    .X(net532));
 sky130_fd_sc_hd__a2111o_1 c497 (.A1(net524),
    .A2(net528),
    .B1(clknet_1_1__leaf_net950),
    .C1(clknet_1_0__leaf_net948),
    .D1(net1072),
    .X(net533));
 sky130_fd_sc_hd__sdfbbn_1 c498 (.CLK_N(clknet_leaf_27_clk),
    .D(net531),
    .RESET_B(net1130),
    .SCD(clknet_1_1__leaf_net526),
    .SCE(net1081),
    .SET_B(net1107),
    .Q(net1065),
    .Q_N(net534));
 sky130_fd_sc_hd__sdfbbn_1 c499 (.CLK_N(clknet_leaf_26_clk),
    .D(clknet_1_0__leaf_net533),
    .RESET_B(clknet_1_1__leaf_net526),
    .SCD(net524),
    .SCE(net534),
    .SET_B(net1064),
    .Q(net1060),
    .Q_N(net535));
 sky130_fd_sc_hd__buf_1 c50 (.A(net1017),
    .X(net26));
 sky130_fd_sc_hd__a2111o_1 c500 (.A1(net527),
    .A2(net535),
    .B1(net951),
    .C1(clknet_1_1__leaf_net950),
    .D1(net1072),
    .X(net1057));
 sky130_fd_sc_hd__mux4_2 c501 (.A0(net1065),
    .A1(clknet_1_1__leaf_net533),
    .A2(net529),
    .A3(clknet_1_0__leaf_net1057),
    .S0(net1059),
    .S1(clknet_1_1__leaf_net950),
    .X(net536));
 sky130_fd_sc_hd__mux4_1 c502 (.A0(clknet_1_0__leaf_net536),
    .A1(net530),
    .A2(net529),
    .A3(clknet_1_1__leaf_net1057),
    .S0(clknet_1_1__leaf_net518),
    .S1(clknet_1_1__leaf_net520),
    .X(net537));
 sky130_fd_sc_hd__mux4_2 c503 (.A0(net529),
    .A1(net1059),
    .A2(clknet_1_1__leaf_net536),
    .A3(net381),
    .S0(clknet_1_1__leaf_net1057),
    .S1(net1063),
    .X(net1055));
 sky130_fd_sc_hd__and2_0 c504 (.A(net414),
    .B(clknet_1_0__leaf_net931),
    .X(net538));
 sky130_fd_sc_hd__and3_1 c505 (.A(net405),
    .B(net414),
    .C(clknet_1_1__leaf_net538),
    .X(net539));
 sky130_fd_sc_hd__and2_0 c506 (.A(clknet_1_0__leaf_net538),
    .B(clknet_1_0__leaf_net539),
    .X(net540));
 sky130_fd_sc_hd__and2_0 c507 (.A(net407),
    .B(clknet_1_1__leaf_net931),
    .X(net541));
 sky130_fd_sc_hd__clkbuf_1 c508 (.A(net795),
    .X(net542));
 sky130_fd_sc_hd__and2_0 c509 (.A(net542),
    .B(clknet_1_1__leaf_net541),
    .X(net543));
 sky130_fd_sc_hd__and2_1 c51 (.A(net26),
    .B(net24),
    .X(net27));
 sky130_fd_sc_hd__and2_0 c510 (.A(clknet_1_0__leaf_net541),
    .B(clknet_1_1__leaf_net543),
    .X(net544));
 sky130_fd_sc_hd__and2_0 c511 (.A(clknet_1_1__leaf_net543),
    .B(clknet_1_1__leaf_net931),
    .X(net545));
 sky130_fd_sc_hd__clkbuf_2 c512 (.A(net795),
    .X(net546));
 sky130_fd_sc_hd__sdfbbp_1 c513 (.CLK(clknet_leaf_45_clk),
    .D(clknet_1_1__leaf_net543),
    .RESET_B(clknet_1_0__leaf_net539),
    .SCD(clknet_1_1__leaf_net545),
    .SCE(clknet_1_1__leaf_net538),
    .SET_B(net546),
    .Q(net548),
    .Q_N(net547));
 sky130_fd_sc_hd__and2_0 c514 (.A(net546),
    .B(clknet_1_0__leaf_net931),
    .X(net549));
 sky130_fd_sc_hd__and2_0 c515 (.A(net546),
    .B(clknet_1_0__leaf_net549),
    .X(net550));
 sky130_fd_sc_hd__sdfbbn_1 c516 (.CLK_N(clknet_leaf_45_clk),
    .D(clknet_1_0__leaf_net538),
    .RESET_B(clknet_1_0__leaf_net544),
    .SCD(clknet_1_0__leaf_net549),
    .SCE(clknet_1_0__leaf_net550),
    .SET_B(clknet_1_0__leaf_net543),
    .Q(net552),
    .Q_N(net551));
 sky130_fd_sc_hd__a2111o_1 c517 (.A1(clknet_1_1__leaf_net539),
    .A2(net552),
    .B1(net548),
    .C1(clknet_1_0__leaf_net550),
    .D1(net546),
    .X(net553));
 sky130_fd_sc_hd__sdfbbn_1 c518 (.CLK_N(clknet_leaf_45_clk),
    .D(net1136),
    .RESET_B(clknet_1_0__leaf_net550),
    .SCD(clknet_1_0__leaf_net540),
    .SCE(net546),
    .SET_B(clknet_1_0__leaf_net543),
    .Q(net555),
    .Q_N(net554));
 sky130_fd_sc_hd__and3_1 c519 (.A(clknet_1_0__leaf_net550),
    .B(net554),
    .C(clknet_1_1__leaf_net549),
    .X(net556));
 sky130_fd_sc_hd__and3_1 c52 (.A(net24),
    .B(net25),
    .C(net27),
    .X(net28));
 sky130_fd_sc_hd__mux4_1 c520 (.A0(clknet_1_1__leaf_net549),
    .A1(clknet_1_1__leaf_net544),
    .A2(net546),
    .A3(clknet_1_1__leaf_net550),
    .S0(net547),
    .S1(clknet_1_0__leaf_net556),
    .X(net557));
 sky130_fd_sc_hd__sdfbbp_1 c521 (.CLK(clknet_leaf_45_clk),
    .D(clknet_1_0__leaf_net553),
    .RESET_B(net548),
    .SCD(net551),
    .SCE(clknet_1_0__leaf_net550),
    .SET_B(clknet_1_1__leaf_net539),
    .Q(net559),
    .Q_N(net558));
 sky130_fd_sc_hd__mux4_1 c522 (.A0(net555),
    .A1(net558),
    .A2(clknet_1_1__leaf_net550),
    .A3(clknet_1_1__leaf_net539),
    .S0(net546),
    .S1(net954),
    .X(net560));
 sky130_fd_sc_hd__mux4_1 c523 (.A0(net559),
    .A1(net546),
    .A2(clknet_1_1__leaf_net560),
    .A3(clknet_1_1__leaf_net550),
    .S0(clknet_1_1__leaf_net931),
    .S1(net955),
    .X(net561));
 sky130_fd_sc_hd__mux4_1 c524 (.A0(clknet_1_0__leaf_net560),
    .A1(clknet_1_1__leaf_net556),
    .A2(clknet_1_1__leaf_net553),
    .A3(net546),
    .S0(clknet_1_1__leaf_net550),
    .S1(net956),
    .X(net562));
 sky130_fd_sc_hd__and2_2 c525 (.A(net442),
    .B(net405),
    .X(net563));
 sky130_fd_sc_hd__clkbuf_2 c526 (.A(net775),
    .X(net564));
 sky130_fd_sc_hd__dfbbn_1 c527 (.CLK_N(clknet_leaf_42_clk),
    .D(net563),
    .RESET_B(net442),
    .SET_B(net1127),
    .Q(net566),
    .Q_N(net565));
 sky130_fd_sc_hd__and3_2 c528 (.A(net564),
    .B(net565),
    .C(net442),
    .X(net567));
 sky130_fd_sc_hd__and2_1 c529 (.A(net566),
    .B(net564),
    .X(net568));
 sky130_fd_sc_hd__or4bb_4 c53 (.A(net18),
    .B(net1080),
    .C_N(net26),
    .D_N(net24),
    .X(net29));
 sky130_fd_sc_hd__buf_1 c530 (.A(net1018),
    .X(net569));
 sky130_fd_sc_hd__and2_1 c531 (.A(net569),
    .B(net568),
    .X(net570));
 sky130_fd_sc_hd__mux4_1 c532 (.A0(net566),
    .A1(net296),
    .A2(net563),
    .A3(net564),
    .S0(net1069),
    .S1(net568),
    .X(net571));
 sky130_fd_sc_hd__clkbuf_1 c533 (.A(net775),
    .X(net572));
 sky130_fd_sc_hd__and3_1 c534 (.A(net564),
    .B(net569),
    .C(net957),
    .X(net573));
 sky130_fd_sc_hd__sdfstp_1 c535 (.CLK(clknet_leaf_42_clk),
    .D(net573),
    .SCD(net570),
    .SCE(net567),
    .SET_B(net1099),
    .Q(net574));
 sky130_fd_sc_hd__sedfxbp_1 c536 (.CLK(clknet_leaf_42_clk),
    .D(net569),
    .DE(net564),
    .SCD(net567),
    .SCE(net563),
    .Q(net576),
    .Q_N(net575));
 sky130_fd_sc_hd__sdfbbn_1 c537 (.CLK_N(clknet_leaf_41_clk),
    .D(net572),
    .RESET_B(net563),
    .SCD(net576),
    .SCE(net564),
    .SET_B(net442),
    .Q(net577));
 sky130_fd_sc_hd__mux4_1 c538 (.A0(net568),
    .A1(net575),
    .A2(net570),
    .A3(net1069),
    .S0(net563),
    .S1(net1148),
    .X(net578));
 sky130_fd_sc_hd__and2_1 c539 (.A(net576),
    .B(net565),
    .X(net579));
 sky130_fd_sc_hd__sdfbbp_1 c54 (.CLK(clknet_leaf_11_clk),
    .D(net27),
    .RESET_B(net25),
    .SCD(net29),
    .SCE(net24),
    .SET_B(net9),
    .Q(net31),
    .Q_N(net30));
 sky130_fd_sc_hd__or4bb_1 c540 (.A(net579),
    .B(net569),
    .C_N(net570),
    .D_N(net575),
    .X(net580));
 sky130_fd_sc_hd__mux4_1 c541 (.A0(net574),
    .A1(net564),
    .A2(net580),
    .A3(net579),
    .S0(net568),
    .S1(net563),
    .X(net581));
 sky130_fd_sc_hd__mux4_1 c542 (.A0(net577),
    .A1(net580),
    .A2(net579),
    .A3(net564),
    .S0(net575),
    .S1(net960),
    .X(net582));
 sky130_fd_sc_hd__sdfbbn_1 c543 (.CLK_N(clknet_leaf_42_clk),
    .D(net576),
    .RESET_B(net580),
    .SCD(net579),
    .SCE(net1148),
    .SET_B(net962),
    .Q(net584),
    .Q_N(net583));
 sky130_fd_sc_hd__mux4_1 c544 (.A0(net580),
    .A1(net583),
    .A2(net564),
    .A3(net563),
    .S0(net579),
    .S1(net1140),
    .X(net585));
 sky130_fd_sc_hd__mux4_1 c545 (.A0(net584),
    .A1(net567),
    .A2(net580),
    .A3(net579),
    .S0(net961),
    .S1(net1146),
    .X(net586));
 sky130_fd_sc_hd__buf_4 c546 (.X(net587));
 sky130_fd_sc_hd__clkbuf_1 c547 (.A(net791),
    .X(net588));
 sky130_fd_sc_hd__and3_2 c548 (.A(net570),
    .B(net1075),
    .C(net964),
    .X(net589));
 sky130_fd_sc_hd__dfbbn_1 c549 (.CLK_N(clknet_leaf_41_clk),
    .D(net567),
    .RESET_B(net1075),
    .SET_B(net960),
    .Q(net591),
    .Q_N(net590));
 sky130_fd_sc_hd__sdfrbp_1 c55 (.CLK(clknet_leaf_11_clk),
    .D(net31),
    .RESET_B(net1110),
    .SCD(net28),
    .SCE(net24),
    .Q(net33),
    .Q_N(net32));
 sky130_fd_sc_hd__sedfxbp_1 c550 (.CLK(clknet_leaf_40_clk),
    .D(net589),
    .DE(net456),
    .SCD(net590),
    .SCE(net1076),
    .Q(net592));
 sky130_fd_sc_hd__sdfbbp_1 c551 (.CLK(clknet_leaf_39_clk),
    .D(net1120),
    .RESET_B(net589),
    .SCD(clknet_1_0__leaf_net454),
    .SCE(net590),
    .SET_B(net1076),
    .Q(net593));
 sky130_fd_sc_hd__and2_0 c552 (.A(net591),
    .B(net941),
    .X(net594));
 sky130_fd_sc_hd__clkbuf_1 c553 (.A(net817),
    .X(net595));
 sky130_fd_sc_hd__and2_0 c554 (.A(net591),
    .B(net1075),
    .X(net596));
 sky130_fd_sc_hd__and2_1 c555 (.A(net588),
    .B(net591),
    .X(net597));
 sky130_fd_sc_hd__and2_0 c556 (.A(net597),
    .B(net1068),
    .X(net598));
 sky130_fd_sc_hd__mux4_1 c557 (.A0(net596),
    .A1(net591),
    .A2(net589),
    .A3(net595),
    .S0(net597),
    .S1(net1075),
    .X(net599));
 sky130_fd_sc_hd__and2_2 c558 (.A(net596),
    .B(net590),
    .X(net600));
 sky130_fd_sc_hd__and3_1 c559 (.A(net594),
    .B(net600),
    .C(net1075),
    .X(net601));
 sky130_fd_sc_hd__sdfbbn_1 c56 (.CLK_N(clknet_leaf_11_clk),
    .D(net21),
    .RESET_B(net24),
    .SCD(net26),
    .SCE(net27),
    .SET_B(net29),
    .Q(net35),
    .Q_N(net34));
 sky130_fd_sc_hd__mux4_1 c560 (.A0(net595),
    .A1(net600),
    .A2(net589),
    .A3(net590),
    .S0(net1075),
    .S1(net1137),
    .X(net602));
 sky130_fd_sc_hd__sedfxtp_1 c561 (.CLK(clknet_leaf_41_clk),
    .D(net1069),
    .DE(net1075),
    .SCD(net600),
    .SCE(net589),
    .Q(net603));
 sky130_fd_sc_hd__sedfxtp_1 c562 (.CLK(clknet_leaf_39_clk),
    .D(net601),
    .DE(net591),
    .SCD(net600),
    .SCE(net1075),
    .Q(net604));
 sky130_fd_sc_hd__sedfxtp_1 c563 (.CLK(clknet_leaf_43_clk),
    .D(net595),
    .DE(net589),
    .SCD(net600),
    .SCE(net1075),
    .Q(net605));
 sky130_fd_sc_hd__a2111o_1 c564 (.A1(net604),
    .A2(net605),
    .B1(net600),
    .C1(net1076),
    .D1(net966),
    .X(net606));
 sky130_fd_sc_hd__mux4_1 c565 (.A0(net1183),
    .A1(net604),
    .A2(net605),
    .A3(net606),
    .S0(net1076),
    .S1(net600),
    .X(net607));
 sky130_fd_sc_hd__sdfbbn_1 c566 (.CLK_N(clknet_leaf_37_clk),
    .D(net605),
    .RESET_B(net606),
    .SCD(net600),
    .SCE(net589),
    .SET_B(net1076),
    .Q(net608));
 sky130_fd_sc_hd__and2_0 c567 (.A(net1075),
    .B(net967),
    .X(net609));
 sky130_fd_sc_hd__and2_0 c568 (.A(clknet_1_1__leaf_net609),
    .B(net1076),
    .X(net610));
 sky130_fd_sc_hd__and2_0 c569 (.A(net600),
    .B(clknet_1_0__leaf_net610),
    .X(net611));
 sky130_fd_sc_hd__sdfbbn_1 c57 (.CLK_N(clknet_leaf_11_clk),
    .D(net1138),
    .RESET_B(net28),
    .SCD(net30),
    .SCE(net29),
    .SET_B(net24),
    .Q(net37),
    .Q_N(net36));
 sky130_fd_sc_hd__clkbuf_1 c570 (.A(net786),
    .X(net612));
 sky130_fd_sc_hd__and2_0 c571 (.A(clknet_1_1__leaf_net609),
    .B(net946),
    .X(net613));
 sky130_fd_sc_hd__buf_1 c572 (.A(net786),
    .X(net614));
 sky130_fd_sc_hd__and3_1 c573 (.A(clknet_1_0__leaf_net610),
    .B(net614),
    .C(clknet_1_0__leaf_net613),
    .X(net615));
 sky130_fd_sc_hd__sdfrbp_1 c574 (.CLK(clknet_leaf_39_clk),
    .D(net614),
    .RESET_B(clknet_1_1__leaf_net615),
    .SCD(clknet_1_1__leaf_net613),
    .SCE(clknet_1_0__leaf_net609),
    .Q(net616));
 sky130_fd_sc_hd__and2_0 c575 (.A(net612),
    .B(net614),
    .X(net617));
 sky130_fd_sc_hd__sdfrbp_1 c576 (.CLK(clknet_leaf_39_clk),
    .D(clknet_1_1__leaf_net611),
    .RESET_B(net614),
    .SCD(clknet_1_0__leaf_net615),
    .SCE(clknet_1_0__leaf_net613),
    .Q(net619),
    .Q_N(net618));
 sky130_fd_sc_hd__a2111o_1 c577 (.A1(clknet_1_0__leaf_net609),
    .A2(clknet_1_0__leaf_net613),
    .B1(net614),
    .C1(clknet_1_1__leaf_net610),
    .D1(net619),
    .X(net620));
 sky130_fd_sc_hd__clkbuf_1 c578 (.A(net824),
    .X(net621));
 sky130_fd_sc_hd__and2_0 c579 (.A(net617),
    .B(clknet_1_0__leaf_net613),
    .X(net622));
 sky130_fd_sc_hd__mux4_1 c58 (.A0(net28),
    .A1(net29),
    .A2(net35),
    .A3(net36),
    .S0(net22),
    .S1(net32),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_1 c580 (.A(net824),
    .X(net623));
 sky130_fd_sc_hd__sdfbbn_1 c581 (.CLK_N(clknet_leaf_39_clk),
    .D(net620),
    .RESET_B(net621),
    .SCD(clknet_1_1__leaf_net615),
    .SCE(clknet_1_0__leaf_net622),
    .SET_B(clknet_1_1__leaf_net613),
    .Q(net625),
    .Q_N(net624));
 sky130_fd_sc_hd__and3_1 c582 (.A(net625),
    .B(clknet_1_1__leaf_net610),
    .C(net947),
    .X(net626));
 sky130_fd_sc_hd__and2_1 c583 (.A(net598),
    .B(net625),
    .X(net627));
 sky130_fd_sc_hd__buf_1 c584 (.A(clknet_1_0__leaf_net1026),
    .X(net628));
 sky130_fd_sc_hd__sdfrtn_1 c585 (.CLK_N(clknet_leaf_30_clk),
    .D(clknet_1_0__leaf_net622),
    .RESET_B(clknet_1_1__leaf_net628),
    .SCD(net627),
    .SCE(clknet_1_1__leaf_net613),
    .Q(net629));
 sky130_fd_sc_hd__mux4_1 c586 (.A0(net616),
    .A1(net623),
    .A2(net627),
    .A3(net624),
    .S0(clknet_1_0__leaf_net622),
    .S1(clknet_1_0__leaf_net628),
    .X(net630));
 sky130_fd_sc_hd__mux4_1 c587 (.A0(net629),
    .A1(clknet_1_1__leaf_net628),
    .A2(net627),
    .A3(clknet_1_1__leaf_net613),
    .S0(clknet_1_0__leaf_net626),
    .S1(net968),
    .X(net631));
 sky130_fd_sc_hd__clkbuf_2 c588 (.A(net784),
    .X(net632));
 sky130_fd_sc_hd__and2_0 c589 (.A(net632),
    .B(clknet_1_1__leaf_net948),
    .X(net633));
 sky130_fd_sc_hd__mux4_1 c59 (.A0(net37),
    .A1(net1053),
    .A2(net31),
    .A3(net19),
    .S0(net24),
    .S1(net29),
    .X(net39));
 sky130_fd_sc_hd__and2_0 c590 (.A(net632),
    .B(net1077),
    .X(net634));
 sky130_fd_sc_hd__and2_0 c591 (.A(net634),
    .B(net632),
    .X(net635));
 sky130_fd_sc_hd__and2_0 c592 (.A(net632),
    .B(net634),
    .X(net636));
 sky130_fd_sc_hd__and2_0 c593 (.A(net635),
    .B(net226),
    .X(net637));
 sky130_fd_sc_hd__and3_1 c594 (.A(clknet_1_1__leaf_net633),
    .B(net635),
    .C(net944),
    .X(net638));
 sky130_fd_sc_hd__and2_0 c595 (.A(clknet_1_0__leaf_net633),
    .B(net635),
    .X(net639));
 sky130_fd_sc_hd__buf_1 c596 (.A(net783),
    .X(net640));
 sky130_fd_sc_hd__clkbuf_2 c597 (.A(net1013),
    .X(net641));
 sky130_fd_sc_hd__sdfbbp_1 c598 (.CLK(clknet_leaf_31_clk),
    .D(clknet_1_1__leaf_net626),
    .RESET_B(net636),
    .SCD(net641),
    .SCE(net632),
    .SET_B(clknet_1_0__leaf_net639),
    .Q(net642));
 sky130_fd_sc_hd__dfbbp_1 c599 (.CLK(clknet_leaf_31_clk),
    .D(net637),
    .RESET_B(clknet_1_0__leaf_net639),
    .SET_B(net641),
    .Q(net644),
    .Q_N(net643));
 sky130_fd_sc_hd__sdfbbp_1 c60 (.CLK(clknet_leaf_10_clk),
    .D(net24),
    .RESET_B(net18),
    .SCD(net37),
    .SCE(net20),
    .SET_B(net19),
    .Q(net40));
 sky130_fd_sc_hd__clkbuf_1 c600 (.A(net1012),
    .X(net645));
 sky130_fd_sc_hd__sdfxbp_1 c601 (.CLK(clknet_leaf_33_clk),
    .D(net642),
    .SCD(net644),
    .SCE(clknet_1_0__leaf_net639),
    .Q(net647),
    .Q_N(net646));
 sky130_fd_sc_hd__sdfbbn_1 c602 (.CLK_N(clknet_leaf_27_clk),
    .D(net647),
    .RESET_B(net645),
    .SCD(clknet_1_1__leaf_net639),
    .SCE(net641),
    .SET_B(clknet_1_1__leaf_net948),
    .Q(net648));
 sky130_fd_sc_hd__mux4_1 c603 (.A0(net638),
    .A1(clknet_1_1__leaf_net639),
    .A2(net643),
    .A3(net646),
    .S0(net640),
    .S1(net641),
    .X(net649));
 sky130_fd_sc_hd__mux4_1 c604 (.A0(net645),
    .A1(net1077),
    .A2(net641),
    .A3(net647),
    .S0(clknet_1_1__leaf_net626),
    .S1(net971),
    .X(net650));
 sky130_fd_sc_hd__mux4_1 c605 (.A0(net636),
    .A1(net647),
    .A2(clknet_1_1__leaf_net639),
    .A3(net641),
    .S0(net640),
    .S1(net973),
    .X(net651));
 sky130_fd_sc_hd__mux4_1 c606 (.A0(net640),
    .A1(net647),
    .A2(net645),
    .A3(net632),
    .S0(clknet_1_1__leaf_net639),
    .S1(net974),
    .X(net652));
 sky130_fd_sc_hd__mux4_2 c607 (.A0(net648),
    .A1(net641),
    .A2(net646),
    .A3(net970),
    .S0(net972),
    .S1(net975),
    .X(net1066));
 sky130_fd_sc_hd__mux4_1 c608 (.A0(net508),
    .A1(net646),
    .A2(net1066),
    .A3(net641),
    .S0(net971),
    .S1(net973),
    .X(net653));
 sky130_fd_sc_hd__a2111o_1 c61 (.A1(net40),
    .A2(net37),
    .B1(net34),
    .C1(net24),
    .D1(clknet_1_0__leaf_net871),
    .X(net41));
 sky130_fd_sc_hd__mux4_1 c62 (.A0(net41),
    .A1(net33),
    .A2(net20),
    .A3(net29),
    .S0(net36),
    .S1(clknet_1_1__leaf_net871),
    .X(net42));
 sky130_fd_sc_hd__mux4_1 c629 (.A0(net396),
    .A1(net381),
    .A2(net1066),
    .A3(clknet_1_0__leaf_net1055),
    .S0(clknet_1_1__leaf_net1057),
    .S1(net953),
    .X(net654));
 sky130_fd_sc_hd__and2_1 c63 (.A(net45),
    .B(net25),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_2 c630 (.A(net957),
    .X(net655));
 sky130_fd_sc_hd__and2_1 c631 (.A(net655),
    .B(net957),
    .X(net656));
 sky130_fd_sc_hd__and2_1 c632 (.A(net1071),
    .B(net957),
    .X(net657));
 sky130_fd_sc_hd__clkbuf_1 c633 (.A(net785),
    .X(net658));
 sky130_fd_sc_hd__and2_0 c634 (.A(net658),
    .B(net655),
    .X(net659));
 sky130_fd_sc_hd__dlymetal6s2s_1 c635 (.A(net785),
    .X(net660));
 sky130_fd_sc_hd__and3_1 c636 (.A(net659),
    .B(net1071),
    .C(net660),
    .X(net661));
 sky130_fd_sc_hd__sdfxbp_1 c637 (.CLK(clknet_leaf_44_clk),
    .D(net661),
    .SCD(net655),
    .SCE(net957),
    .Q(net663),
    .Q_N(net662));
 sky130_fd_sc_hd__sdfxtp_1 c638 (.CLK(clknet_leaf_44_clk),
    .D(net657),
    .SCD(net660),
    .SCE(net662),
    .Q(net664));
 sky130_fd_sc_hd__mux4_1 c639 (.A0(net663),
    .A1(net664),
    .A2(net655),
    .A3(net660),
    .S0(net1071),
    .S1(net661),
    .X(net665));
 sky130_fd_sc_hd__and2_1 c64 (.A(net45),
    .B(net25),
    .X(net44));
 sky130_fd_sc_hd__and3_1 c640 (.A(net1071),
    .B(net660),
    .C(net976),
    .X(net666));
 sky130_fd_sc_hd__sdfrtp_1 c641 (.CLK(clknet_leaf_44_clk),
    .D(net655),
    .RESET_B(net1086),
    .SCD(net657),
    .SCE(net1164),
    .Q(net667));
 sky130_fd_sc_hd__a2111o_2 c642 (.A1(net667),
    .A2(net664),
    .B1(net1071),
    .C1(net662),
    .D1(net957),
    .X(net668));
 sky130_fd_sc_hd__mux4_1 c643 (.A0(net668),
    .A1(net666),
    .A2(net663),
    .A3(net660),
    .S0(net1071),
    .S1(net655),
    .X(net669));
 sky130_fd_sc_hd__mux4_1 c644 (.A0(net666),
    .A1(net659),
    .A2(net663),
    .A3(net668),
    .S0(net656),
    .S1(net657),
    .X(net670));
 sky130_fd_sc_hd__clkbuf_1 c645 (.A(net819),
    .X(net671));
 sky130_fd_sc_hd__sdfxtp_1 c646 (.CLK(clknet_leaf_44_clk),
    .D(net671),
    .SCD(net660),
    .SCE(net668),
    .Q(net672));
 sky130_fd_sc_hd__mux4_1 c647 (.A0(net660),
    .A1(net672),
    .A2(net668),
    .A3(net657),
    .S0(net957),
    .S1(net1167),
    .X(net673));
 sky130_fd_sc_hd__mux4_1 c648 (.A0(net671),
    .A1(net668),
    .A2(net672),
    .A3(net1071),
    .S0(net662),
    .S1(net1165),
    .X(net674));
 sky130_fd_sc_hd__mux4_1 c649 (.A0(net1191),
    .A1(net1190),
    .A2(net1071),
    .A3(net976),
    .S0(net1192),
    .S1(net1091),
    .X(net675));
 sky130_fd_sc_hd__and2_1 c65 (.A(net1048),
    .B(net25),
    .X(net45));
 sky130_fd_sc_hd__mux4_1 c650 (.A0(net672),
    .A1(net1071),
    .A2(net405),
    .A3(net978),
    .S0(net980),
    .S1(net981),
    .X(net676));
 sky130_fd_sc_hd__buf_2 c651 (.A(net810),
    .X(net677));
 sky130_fd_sc_hd__and2_1 c652 (.A(net677),
    .B(net570),
    .X(net678));
 sky130_fd_sc_hd__and2_0 c653 (.A(net677),
    .B(net977),
    .X(net679));
 sky130_fd_sc_hd__buf_2 c654 (.A(net1018),
    .X(net680));
 sky130_fd_sc_hd__buf_1 c655 (.A(clknet_1_0__leaf_net1028),
    .X(net681));
 sky130_fd_sc_hd__and2_1 c656 (.A(net680),
    .B(net960),
    .X(net682));
 sky130_fd_sc_hd__and2_1 c657 (.A(net680),
    .B(net682),
    .X(net683));
 sky130_fd_sc_hd__and2_2 c658 (.A(net683),
    .B(net1150),
    .X(net684));
 sky130_fd_sc_hd__clkbuf_1 c659 (.A(net1168),
    .X(net685));
 sky130_fd_sc_hd__and2_0 c66 (.A(net45),
    .B(clknet_1_1__leaf_net872),
    .X(net46));
 sky130_fd_sc_hd__sdfxtp_1 c660 (.CLK(clknet_leaf_37_clk),
    .D(net685),
    .SCD(net684),
    .SCE(net680),
    .Q(net686));
 sky130_fd_sc_hd__buf_1 c661 (.A(net809),
    .X(net687));
 sky130_fd_sc_hd__or4bb_1 c662 (.A(net679),
    .B(net683),
    .C_N(net682),
    .D_N(net687),
    .X(net688));
 sky130_fd_sc_hd__clkbuf_1 c663 (.A(net820),
    .X(net689));
 sky130_fd_sc_hd__sdfbbn_1 c664 (.CLK_N(clknet_leaf_43_clk),
    .D(net688),
    .RESET_B(net682),
    .SCD(net683),
    .SCE(net677),
    .SET_B(net687),
    .Q(net690));
 sky130_fd_sc_hd__sdfrtp_1 c665 (.CLK(clknet_leaf_43_clk),
    .D(net677),
    .RESET_B(net1088),
    .SCD(net684),
    .SCE(net683),
    .Q(net691));
 sky130_fd_sc_hd__mux4_1 c666 (.A0(net681),
    .A1(net691),
    .A2(net686),
    .A3(net680),
    .S0(net677),
    .S1(net684),
    .X(net692));
 sky130_fd_sc_hd__mux4_1 c667 (.A0(net690),
    .A1(net684),
    .A2(net682),
    .A3(net680),
    .S0(net960),
    .S1(net983),
    .X(net693));
 sky130_fd_sc_hd__mux4_1 c668 (.A0(net689),
    .A1(net688),
    .A2(net691),
    .A3(net684),
    .S0(net677),
    .S1(net983),
    .X(net694));
 sky130_fd_sc_hd__sdfrtp_1 c669 (.CLK(clknet_leaf_37_clk),
    .D(net677),
    .RESET_B(net684),
    .SCD(net983),
    .SCE(net1174),
    .Q(net695));
 sky130_fd_sc_hd__buf_1 c67 (.A(net798),
    .X(net47));
 sky130_fd_sc_hd__mux4_1 c670 (.A0(net686),
    .A1(net695),
    .A2(net680),
    .A3(net960),
    .S0(net984),
    .S1(net985),
    .X(net696));
 sky130_fd_sc_hd__mux4_1 c671 (.A0(net675),
    .A1(net696),
    .A2(net1178),
    .A3(net684),
    .S0(net983),
    .S1(net1174),
    .X(net697));
 sky130_fd_sc_hd__buf_2 c672 (.A(net608),
    .X(net698));
 sky130_fd_sc_hd__clkbuf_1 c673 (.A(net698),
    .X(net699));
 sky130_fd_sc_hd__and2_0 c674 (.A(net698),
    .B(net986),
    .X(net700));
 sky130_fd_sc_hd__and2_0 c675 (.A(clknet_1_0__leaf_net700),
    .B(net960),
    .X(net701));
 sky130_fd_sc_hd__and2_0 c676 (.A(net699),
    .B(clknet_1_1__leaf_net700),
    .X(net702));
 sky130_fd_sc_hd__clkbuf_1 c677 (.A(net793),
    .X(net703));
 sky130_fd_sc_hd__clkbuf_1 c678 (.A(net793),
    .X(net704));
 sky130_fd_sc_hd__and2_0 c679 (.A(clknet_1_1__leaf_net700),
    .B(net698),
    .X(net705));
 sky130_fd_sc_hd__and3_1 c68 (.A(net45),
    .B(net1070),
    .C(clknet_1_1__leaf_net872),
    .X(net48));
 sky130_fd_sc_hd__and2_0 c680 (.A(net704),
    .B(net703),
    .X(net706));
 sky130_fd_sc_hd__dfbbn_1 c681 (.CLK_N(clknet_leaf_36_clk),
    .D(net706),
    .RESET_B(clknet_1_0__leaf_net702),
    .SET_B(clknet_1_0__leaf_net700),
    .Q(net708),
    .Q_N(net707));
 sky130_fd_sc_hd__and2_0 c682 (.A(net708),
    .B(net704),
    .X(net709));
 sky130_fd_sc_hd__mux4_1 c683 (.A0(clknet_1_0__leaf_net701),
    .A1(net706),
    .A2(net707),
    .A3(net698),
    .S0(clknet_1_0__leaf_net700),
    .S1(clknet_1_0__leaf_net702),
    .X(net710));
 sky130_fd_sc_hd__sdfbbp_1 c684 (.CLK(clknet_leaf_36_clk),
    .D(net703),
    .RESET_B(net709),
    .SCD(clknet_1_1__leaf_net701),
    .SCE(clknet_1_0__leaf_net702),
    .SET_B(clknet_1_0__leaf_net987),
    .Q(net712),
    .Q_N(net711));
 sky130_fd_sc_hd__sdfsbp_1 c685 (.CLK(clknet_leaf_36_clk),
    .D(net712),
    .SCD(net706),
    .SCE(clknet_1_1__leaf_net702),
    .SET_B(clknet_1_0__leaf_net987),
    .Q(net714),
    .Q_N(net713));
 sky130_fd_sc_hd__mux4_1 c686 (.A0(net709),
    .A1(net713),
    .A2(net708),
    .A3(net698),
    .S0(clknet_1_1__leaf_net702),
    .S1(clknet_1_1__leaf_net987),
    .X(net715));
 sky130_fd_sc_hd__mux4_1 c687 (.A0(net714),
    .A1(net712),
    .A2(clknet_1_1__leaf_net702),
    .A3(net707),
    .S0(net698),
    .S1(clknet_1_1__leaf_net987),
    .X(net716));
 sky130_fd_sc_hd__mux4_1 c688 (.A0(clknet_1_0__leaf_net705),
    .A1(net699),
    .A2(net707),
    .A3(net698),
    .S0(clknet_1_1__leaf_net987),
    .S1(net990),
    .X(net717));
 sky130_fd_sc_hd__mux4_1 c689 (.A0(net708),
    .A1(clknet_1_1__leaf_net700),
    .A2(net711),
    .A3(clknet_1_1__leaf_net702),
    .S0(clknet_1_0__leaf_net987),
    .S1(net992),
    .X(net718));
 sky130_fd_sc_hd__clkbuf_1 c69 (.A(net798),
    .X(net49));
 sky130_fd_sc_hd__mux4_1 c690 (.A0(clknet_1_1__leaf_net705),
    .A1(clknet_1_1__leaf_net702),
    .A2(clknet_1_1__leaf_net987),
    .A3(net988),
    .S0(net989),
    .S1(net991),
    .X(net719));
 sky130_fd_sc_hd__mux4_1 c691 (.A0(clknet_1_1__leaf_net700),
    .A1(net1068),
    .A2(net711),
    .A3(net992),
    .S0(net993),
    .S1(net995),
    .X(net720));
 sky130_fd_sc_hd__mux4_1 c692 (.A0(net712),
    .A1(clknet_1_1__leaf_net720),
    .A2(net1077),
    .A3(net990),
    .S0(net994),
    .S1(net995),
    .X(net721));
 sky130_fd_sc_hd__buf_1 c693 (.A(clknet_1_0__leaf_net805),
    .X(net722));
 sky130_fd_sc_hd__buf_1 c694 (.A(clknet_1_1__leaf_net805),
    .X(net723));
 sky130_fd_sc_hd__buf_1 c695 (.A(net835),
    .X(net724));
 sky130_fd_sc_hd__and2_0 c696 (.A(clknet_1_0__leaf_net722),
    .B(net1076),
    .X(net725));
 sky130_fd_sc_hd__clkbuf_1 c697 (.A(net834),
    .X(net726));
 sky130_fd_sc_hd__and2_0 c698 (.A(clknet_1_1__leaf_net723),
    .B(clknet_1_0__leaf_net725),
    .X(net727));
 sky130_fd_sc_hd__and3_1 c699 (.A(net726),
    .B(net698),
    .C(clknet_1_0__leaf_net725),
    .X(net728));
 sky130_fd_sc_hd__dfbbn_2 c70 (.CLK_N(clknet_leaf_12_clk),
    .D(clknet_1_0__leaf_net48),
    .RESET_B(net45),
    .SET_B(net1070),
    .Q(net51),
    .Q_N(net50));
 sky130_fd_sc_hd__or4bb_1 c700 (.A(net724),
    .B(clknet_1_0__leaf_net628),
    .C_N(clknet_1_0__leaf_net727),
    .D_N(clknet_1_0__leaf_net725),
    .X(net729));
 sky130_fd_sc_hd__sdfsbp_1 c701 (.CLK(clknet_leaf_38_clk),
    .D(clknet_1_1__leaf_net722),
    .SCD(clknet_1_0__leaf_net728),
    .SCE(clknet_1_0__leaf_net729),
    .SET_B(clknet_1_0__leaf_net727),
    .Q(net731),
    .Q_N(net730));
 sky130_fd_sc_hd__sdfbbn_1 c702 (.CLK_N(clknet_leaf_38_clk),
    .D(clknet_1_0__leaf_net720),
    .RESET_B(clknet_1_1__leaf_net729),
    .SCD(clknet_1_0__leaf_net727),
    .SCE(net724),
    .SET_B(clknet_1_0__leaf_net725),
    .Q(net733),
    .Q_N(net732));
 sky130_fd_sc_hd__mux4_1 c703 (.A0(net733),
    .A1(net731),
    .A2(clknet_1_0__leaf_net729),
    .A3(clknet_1_1__leaf_net727),
    .S0(clknet_1_0__leaf_net725),
    .S1(clknet_1_1__leaf_net720),
    .X(net734));
 sky130_fd_sc_hd__sdfbbn_1 c704 (.CLK_N(clknet_leaf_38_clk),
    .D(clknet_1_0__leaf_net727),
    .RESET_B(net733),
    .SCD(net726),
    .SCE(clknet_1_0__leaf_net729),
    .SET_B(clknet_1_0__leaf_net725),
    .Q(net736),
    .Q_N(net735));
 sky130_fd_sc_hd__sdfstp_1 c705 (.CLK(clknet_leaf_31_clk),
    .D(clknet_1_0__leaf_net723),
    .SCD(clknet_1_0__leaf_net727),
    .SCE(clknet_1_0__leaf_net626),
    .SET_B(clknet_1_0__leaf_net725),
    .Q(net737));
 sky130_fd_sc_hd__sdfbbp_1 c706 (.CLK(clknet_leaf_31_clk),
    .D(net1139),
    .RESET_B(net724),
    .SCD(net736),
    .SCE(clknet_1_1__leaf_net729),
    .SET_B(clknet_1_0__leaf_net725),
    .Q(net738));
 sky130_fd_sc_hd__sdfbbn_1 c707 (.CLK_N(clknet_leaf_38_clk),
    .D(clknet_1_0__leaf_net729),
    .RESET_B(clknet_1_0__leaf_net728),
    .SCD(net1162),
    .SCE(clknet_1_0__leaf_net727),
    .SET_B(clknet_1_0__leaf_net725),
    .Q(net740),
    .Q_N(net739));
 sky130_fd_sc_hd__clkbuf_1 c708 (.A(net1032),
    .X(net741));
 sky130_fd_sc_hd__mux4_1 c709 (.A0(net741),
    .A1(net737),
    .A2(clknet_1_1__leaf_net729),
    .A3(clknet_1_1__leaf_net727),
    .S0(clknet_1_0__leaf_net725),
    .S1(net997),
    .X(net742));
 sky130_fd_sc_hd__clkbuf_1 c71 (.A(net1023),
    .X(net52));
 sky130_fd_sc_hd__mux4_1 c710 (.A0(net737),
    .A1(clknet_1_0__leaf_net723),
    .A2(clknet_1_0__leaf_net626),
    .A3(clknet_1_1__leaf_net628),
    .S0(clknet_1_1__leaf_net727),
    .S1(net998),
    .X(net743));
 sky130_fd_sc_hd__mux4_1 c711 (.A0(net698),
    .A1(clknet_1_1__leaf_net727),
    .A2(clknet_1_1__leaf_net728),
    .A3(clknet_1_0__leaf_net729),
    .S0(net998),
    .S1(net999),
    .X(net744));
 sky130_fd_sc_hd__mux4_1 c712 (.A0(net736),
    .A1(clknet_1_0__leaf_net729),
    .A2(clknet_1_1__leaf_net727),
    .A3(clknet_1_1__leaf_net725),
    .S0(net999),
    .S1(net1001),
    .X(net745));
 sky130_fd_sc_hd__mux4_1 c713 (.A0(net740),
    .A1(clknet_1_1__leaf_net725),
    .A2(clknet_1_0__leaf_net729),
    .A3(net999),
    .S0(net1000),
    .S1(net1002),
    .X(net746));
 sky130_fd_sc_hd__and2_0 c714 (.A(net653),
    .B(clknet_1_1__leaf_net725),
    .X(net747));
 sky130_fd_sc_hd__clkbuf_1 c715 (.A(net794),
    .X(net748));
 sky130_fd_sc_hd__clkbuf_2 c716 (.A(net794),
    .X(net1061));
 sky130_fd_sc_hd__dfbbn_1 c717 (.CLK_N(clknet_leaf_32_clk),
    .D(net1128),
    .RESET_B(clknet_1_1__leaf_net747),
    .SET_B(net1003),
    .Q(net750),
    .Q_N(net749));
 sky130_fd_sc_hd__dfbbp_1 c718 (.CLK(clknet_leaf_32_clk),
    .D(net1061),
    .RESET_B(clknet_1_1__leaf_net725),
    .SET_B(clknet_1_0__leaf_net747),
    .Q(net752),
    .Q_N(net751));
 sky130_fd_sc_hd__sdfxbp_1 c719 (.CLK(clknet_leaf_32_clk),
    .D(net1184),
    .SCD(net748),
    .SCE(clknet_1_0__leaf_net747),
    .Q(net754),
    .Q_N(net753));
 sky130_fd_sc_hd__buf_1 c72 (.A(net1033),
    .X(net53));
 sky130_fd_sc_hd__and3_1 c720 (.A(net754),
    .B(net749),
    .C(clknet_1_1__leaf_net725),
    .X(net755));
 sky130_fd_sc_hd__or4bb_1 c721 (.A(net731),
    .B(clknet_1_0__leaf_net755),
    .C_N(net750),
    .D_N(net753),
    .X(net756));
 sky130_fd_sc_hd__sdfstp_1 c722 (.CLK(clknet_leaf_32_clk),
    .D(clknet_1_1__leaf_net747),
    .SCD(net754),
    .SCE(net1061),
    .SET_B(clknet_1_1__leaf_net725),
    .Q(net757));
 sky130_fd_sc_hd__mux4_1 c723 (.A0(net757),
    .A1(net752),
    .A2(clknet_1_0__leaf_net756),
    .A3(clknet_1_0__leaf_net747),
    .S0(net754),
    .S1(clknet_1_1__leaf_net725),
    .X(net758));
 sky130_fd_sc_hd__buf_1 c724 (.A(clknet_1_1__leaf_net1026),
    .X(net759));
 sky130_fd_sc_hd__sdfbbn_1 c725 (.CLK_N(clknet_leaf_34_clk),
    .D(net754),
    .RESET_B(clknet_1_1__leaf_net756),
    .SCD(clknet_1_1__leaf_net626),
    .SCE(net1061),
    .SET_B(net1082),
    .Q(net761),
    .Q_N(net760));
 sky130_fd_sc_hd__sdfbbp_1 c726 (.CLK(clknet_leaf_32_clk),
    .D(clknet_1_1__leaf_net725),
    .RESET_B(net1161),
    .SCD(clknet_1_1__leaf_net747),
    .SCE(net1061),
    .SET_B(net1082),
    .Q(net763),
    .Q_N(net762));
 sky130_fd_sc_hd__mux4_1 c727 (.A0(clknet_1_1__leaf_net725),
    .A1(clknet_1_0__leaf_net759),
    .A2(net763),
    .A3(clknet_1_0__leaf_net747),
    .S0(net753),
    .S1(net751),
    .X(net764));
 sky130_fd_sc_hd__sdfbbn_1 c728 (.CLK_N(clknet_leaf_34_clk),
    .D(net748),
    .RESET_B(net1111),
    .SCD(net762),
    .SCE(clknet_1_1__leaf_net747),
    .SET_B(net753),
    .Q(net766),
    .Q_N(net765));
 sky130_fd_sc_hd__or4bb_1 c729 (.A(net763),
    .B(net760),
    .C_N(net765),
    .D_N(net753),
    .X(net767));
 sky130_fd_sc_hd__sdfbbn_1 c73 (.CLK_N(clknet_leaf_12_clk),
    .D(net25),
    .RESET_B(clknet_1_1__leaf_net48),
    .SCD(net45),
    .SCE(net50),
    .SET_B(net44),
    .Q(net55),
    .Q_N(net54));
 sky130_fd_sc_hd__and3_1 c730 (.A(net766),
    .B(net767),
    .C(net1005),
    .X(net1062));
 sky130_fd_sc_hd__or4bb_1 c731 (.A(clknet_1_1__leaf_net759),
    .B(net653),
    .C_N(clknet_1_1__leaf_net725),
    .D_N(net1005),
    .X(net768));
 sky130_fd_sc_hd__and3_1 c732 (.A(net750),
    .B(net767),
    .C(net1062),
    .X(net769));
 sky130_fd_sc_hd__mux4_1 c733 (.A0(clknet_1_1__leaf_net755),
    .A1(net769),
    .A2(clknet_1_1__leaf_net768),
    .A3(clknet_1_1__leaf_net747),
    .S0(net1004),
    .S1(net1005),
    .X(net770));
 sky130_fd_sc_hd__mux4_1 c734 (.A0(clknet_1_0__leaf_net768),
    .A1(net769),
    .A2(net1062),
    .A3(clknet_1_1__leaf_net747),
    .S0(net754),
    .S1(net1006),
    .X(net771));
 sky130_fd_sc_hd__and3_1 c74 (.A(net55),
    .B(net53),
    .C(net1085),
    .X(net56));
 sky130_fd_sc_hd__and3_1 c75 (.A(net56),
    .B(net55),
    .C(net51),
    .X(net57));
 sky130_fd_sc_hd__or4bb_1 c76 (.A(net53),
    .B(net55),
    .C_N(net56),
    .D_N(net1070),
    .X(net58));
 sky130_fd_sc_hd__mux4_1 c77 (.A0(net46),
    .A1(net51),
    .A2(net53),
    .A3(net56),
    .S0(net1070),
    .S1(net54),
    .X(net59));
 sky130_fd_sc_hd__mux4_1 c78 (.A0(net57),
    .A1(net54),
    .A2(net56),
    .A3(net50),
    .S0(net1070),
    .S1(clknet_1_0__leaf_net873),
    .X(net60));
 sky130_fd_sc_hd__mux4_1 c79 (.A0(net58),
    .A1(net55),
    .A2(clknet_1_0__leaf_net60),
    .A3(net45),
    .S0(net1070),
    .S1(clknet_1_0__leaf_net873),
    .X(net61));
 sky130_fd_sc_hd__sdfbbn_1 c80 (.CLK_N(clknet_leaf_13_clk),
    .D(net1070),
    .RESET_B(net56),
    .SCD(clknet_1_0__leaf_net60),
    .SCE(net54),
    .SET_B(clknet_1_0__leaf_net873),
    .Q(net62));
 sky130_fd_sc_hd__mux4_1 c81 (.A0(net49),
    .A1(clknet_1_0__leaf_net60),
    .A2(net53),
    .A3(net1070),
    .S0(clknet_1_1__leaf_net873),
    .S1(net875),
    .X(net63));
 sky130_fd_sc_hd__mux4_1 c82 (.A0(net52),
    .A1(net62),
    .A2(clknet_1_1__leaf_net60),
    .A3(clknet_1_1__leaf_net872),
    .S0(clknet_1_1__leaf_net873),
    .S1(net874),
    .X(net64));
 sky130_fd_sc_hd__sdfbbp_1 c83 (.CLK(clknet_leaf_13_clk),
    .D(clknet_1_1__leaf_net60),
    .RESET_B(net54),
    .SCD(clknet_1_1__leaf_net873),
    .SCE(net876),
    .SET_B(net1090),
    .Q(net66),
    .Q_N(net65));
 sky130_fd_sc_hd__and2_0 c84 (.A(net66),
    .B(clknet_1_1__leaf_net872),
    .X(net67));
 sky130_fd_sc_hd__and2_0 c85 (.A(clknet_1_0__leaf_net67),
    .B(net65),
    .X(net68));
 sky130_fd_sc_hd__and2_0 c86 (.A(clknet_1_0__leaf_net68),
    .B(net65),
    .X(net69));
 sky130_fd_sc_hd__and2_0 c87 (.A(clknet_1_0__leaf_net67),
    .B(clknet_1_0__leaf_net68),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_1 c88 (.A(net799),
    .X(net71));
 sky130_fd_sc_hd__dlymetal6s2s_1 c89 (.A(net799),
    .X(net72));
 sky130_fd_sc_hd__sdfrbp_1 c90 (.CLK(clknet_leaf_20_clk),
    .D(clknet_1_0__leaf_net69),
    .RESET_B(net1092),
    .SCD(clknet_1_0__leaf_net70),
    .SCE(clknet_1_0__leaf_net68),
    .Q(net74),
    .Q_N(net73));
 sky130_fd_sc_hd__and2_0 c91 (.A(clknet_1_0__leaf_net68),
    .B(net65),
    .X(net75));
 sky130_fd_sc_hd__sdfrtn_1 c92 (.CLK_N(clknet_leaf_21_clk),
    .D(net74),
    .RESET_B(net72),
    .SCD(clknet_1_1__leaf_net75),
    .SCE(clknet_1_1__leaf_net68),
    .Q(net76));
 sky130_fd_sc_hd__mux4_1 c93 (.A0(net76),
    .A1(net71),
    .A2(net66),
    .A3(clknet_1_0__leaf_net68),
    .S0(net72),
    .S1(clknet_1_1__leaf_net70),
    .X(net77));
 sky130_fd_sc_hd__sdfbbn_1 c94 (.CLK_N(clknet_leaf_20_clk),
    .D(clknet_1_0__leaf_net70),
    .RESET_B(net1106),
    .SCD(clknet_1_0__leaf_net68),
    .SCE(clknet_1_0__leaf_net69),
    .SET_B(net65),
    .Q(net79),
    .Q_N(net78));
 sky130_fd_sc_hd__sdfbbn_1 c95 (.CLK_N(clknet_leaf_20_clk),
    .D(net66),
    .RESET_B(clknet_1_0__leaf_net70),
    .SCD(clknet_1_0__leaf_net69),
    .SCE(net78),
    .SET_B(clknet_1_0__leaf_net68),
    .Q(net81),
    .Q_N(net80));
 sky130_fd_sc_hd__sdfbbp_1 c96 (.CLK(clknet_leaf_20_clk),
    .D(net72),
    .RESET_B(clknet_1_1__leaf_net67),
    .SCD(clknet_1_1__leaf_net69),
    .SCE(clknet_1_1__leaf_net68),
    .SET_B(net878),
    .Q(net83),
    .Q_N(net82));
 sky130_fd_sc_hd__mux4_1 c97 (.A0(net83),
    .A1(net80),
    .A2(net76),
    .A3(clknet_1_1__leaf_net69),
    .S0(clknet_1_1__leaf_net68),
    .S1(net878),
    .X(net84));
 sky130_fd_sc_hd__sdfbbn_1 c98 (.CLK_N(clknet_leaf_21_clk),
    .D(clknet_1_0__leaf_net75),
    .RESET_B(net1121),
    .SCD(clknet_1_1__leaf_net68),
    .SCE(net878),
    .SET_B(net1141),
    .Q(net86),
    .Q_N(net85));
 sky130_fd_sc_hd__mux4_1 c99 (.A0(net71),
    .A1(clknet_1_1__leaf_net68),
    .A2(net83),
    .A3(clknet_1_1__leaf_net70),
    .S0(net85),
    .S1(net879),
    .X(net87));
 sky130_fd_sc_hd__sdfbbn_2 merge740 (.CLK_N(clknet_leaf_17_clk),
    .D(clknet_1_1__leaf_net454),
    .RESET_B(net187),
    .SCD(net1068),
    .SCE(net1069),
    .Q(net470),
    .Q_N(net772));
 sky130_fd_sc_hd__buf_1 merge741 (.A(net1024),
    .X(net774));
 sky130_fd_sc_hd__clkbuf_1 merge742 (.A(net1011),
    .X(net775));
 sky130_fd_sc_hd__sdfbbp_1 merge743 (.CLK(clknet_leaf_22_clk),
    .D(net104),
    .RESET_B(net227),
    .SCD(net230),
    .SCE(net231),
    .Q(net228),
    .Q_N(net776));
 sky130_fd_sc_hd__sdfstp_1 merge744 (.CLK(clknet_leaf_15_clk),
    .D(net184),
    .SCD(net50),
    .SCE(net186),
    .SET_B(clknet_1_0__leaf_net872),
    .Q(net778));
 sky130_fd_sc_hd__sedfxbp_1 merge745 (.CLK(clknet_leaf_6_clk),
    .D(net299),
    .DE(net179),
    .SCD(net300),
    .SCE(net298),
    .Q(net780),
    .Q_N(net779));
 sky130_fd_sc_hd__sdfbbn_1 merge746 (.CLK_N(clknet_leaf_8_clk),
    .D(net125),
    .RESET_B(net1049),
    .SCD(net118),
    .SCE(net119),
    .SET_B(net116),
    .Q(net782),
    .Q_N(net781));
 sky130_fd_sc_hd__sdfxbp_1 merge747 (.CLK(clknet_leaf_31_clk),
    .D(clknet_1_1__leaf_net626),
    .SCD(clknet_1_0__leaf_net639),
    .SCE(net969),
    .Q(net784),
    .Q_N(net783));
 sky130_fd_sc_hd__sdfxtp_1 merge748 (.CLK(clknet_leaf_44_clk),
    .D(net657),
    .SCD(net1071),
    .SCE(net655),
    .Q(net785));
 sky130_fd_sc_hd__clkbuf_1 merge749 (.A(net1010),
    .X(net786));
 sky130_fd_sc_hd__sdfxtp_1 merge750 (.CLK(clknet_leaf_15_clk),
    .D(clknet_1_0__leaf_net161),
    .SCD(clknet_1_1__leaf_net160),
    .SCE(net1085),
    .Q(net787));
 sky130_fd_sc_hd__clkbuf_1 merge751 (.A(net818),
    .X(net788));
 sky130_fd_sc_hd__clkbuf_1 merge752 (.A(net1034),
    .X(net789));
 sky130_fd_sc_hd__clkbuf_1 merge753 (.A(net1014),
    .X(net790));
 sky130_fd_sc_hd__sedfxbp_2 merge754 (.CLK(clknet_leaf_41_clk),
    .D(net423),
    .SCD(net567),
    .SCE(net957),
    .Q(net587),
    .Q_N(net791));
 sky130_fd_sc_hd__clkbuf_1 merge755 (.A(net823),
    .X(net793));
 sky130_fd_sc_hd__clkbuf_1 merge756 (.A(net1025),
    .X(net794));
 sky130_fd_sc_hd__sedfxtp_1 merge757 (.CLK(clknet_leaf_45_clk),
    .D(clknet_1_1__leaf_net540),
    .DE(clknet_1_1__leaf_net538),
    .SCD(clknet_1_0__leaf_net545),
    .SCE(clknet_1_0__leaf_net931),
    .Q(net795));
 sky130_fd_sc_hd__sedfxtp_1 merge758 (.CLK(clknet_leaf_5_clk),
    .D(net274),
    .DE(net272),
    .SCD(net280),
    .SCE(net278),
    .Q(net796));
 sky130_fd_sc_hd__mux4_1 merge759 (.A0(net373),
    .A1(net374),
    .A2(net227),
    .A3(net368),
    .S0(net375),
    .S1(net904),
    .X(net797));
 sky130_fd_sc_hd__clkbuf_1 merge760 (.A(net830),
    .X(net798));
 sky130_fd_sc_hd__sdfxtp_1 merge761 (.CLK(clknet_leaf_20_clk),
    .D(clknet_1_0__leaf_net70),
    .SCD(clknet_1_0__leaf_net69),
    .SCE(clknet_1_0__leaf_net68),
    .Q(net799));
 sky130_fd_sc_hd__sdfbbn_2 merge762 (.CLK_N(clknet_leaf_7_clk),
    .D(clknet_1_0__leaf_net138),
    .RESET_B(net1080),
    .SCD(clknet_1_1__leaf_net141),
    .SCE(clknet_1_0__leaf_net139),
    .Q(net140),
    .Q_N(net800));
 sky130_fd_sc_hd__sedfxtp_1 merge763 (.CLK(clknet_leaf_20_clk),
    .D(net195),
    .DE(net65),
    .SCD(net207),
    .SCE(net1124),
    .Q(net802));
 sky130_fd_sc_hd__sdfbbp_1 merge764 (.CLK(clknet_leaf_8_clk),
    .D(net1043),
    .RESET_B(net4),
    .SCD(net1038),
    .SCE(net1046),
    .Q(net6),
    .Q_N(net803));
 sky130_fd_sc_hd__buf_1 merge765 (.A(clknet_1_1__leaf_net1028),
    .X(net805));
 sky130_fd_sc_hd__clkbuf_1 merge766 (.A(net841),
    .X(net806));
 sky130_fd_sc_hd__clkbuf_1 merge767 (.A(net1016),
    .X(net807));
 sky130_fd_sc_hd__clkbuf_1 merge768 (.A(net827),
    .X(net808));
 sky130_fd_sc_hd__sdfrbp_1 merge769 (.CLK(clknet_leaf_43_clk),
    .D(net570),
    .RESET_B(net675),
    .SCD(net684),
    .SCE(net683),
    .Q(net810),
    .Q_N(net809));
 sky130_fd_sc_hd__buf_6 merge770 (.A(net1030),
    .X(net811));
 sky130_fd_sc_hd__sdfbbn_1 merge771 (.CLK_N(clknet_leaf_18_clk),
    .D(net330),
    .RESET_B(net332),
    .SCD(net350),
    .SCE(net351),
    .SET_B(net349),
    .Q(net813),
    .Q_N(net812));
 sky130_fd_sc_hd__dfbbn_1 merge772 (.CLK_N(clknet_leaf_1_clk),
    .D(net253),
    .RESET_B(net250),
    .SET_B(net251),
    .Q(net815),
    .Q_N(net814));
 sky130_fd_sc_hd__mux4_1 merge773 (.A0(net119),
    .A1(net1047),
    .A2(net115),
    .A3(net117),
    .S0(net120),
    .S1(net123),
    .X(net816));
 sky130_fd_sc_hd__sdfrbp_1 merge774 (.CLK(clknet_leaf_3_clk),
    .D(net271),
    .RESET_B(net397),
    .SCD(net593),
    .SCE(net589),
    .Q(net818),
    .Q_N(net817));
 sky130_fd_sc_hd__sdfbbn_1 merge775 (.CLK_N(clknet_leaf_43_clk),
    .D(net687),
    .RESET_B(net684),
    .SCD(net662),
    .SCE(net668),
    .SET_B(net978),
    .Q(net820),
    .Q_N(net819));
 sky130_fd_sc_hd__sdfrtn_1 merge776 (.CLK_N(clknet_leaf_14_clk),
    .D(net184),
    .RESET_B(net187),
    .SCD(net207),
    .SCE(net203),
    .Q(net821));
 sky130_fd_sc_hd__sdfbbp_1 merge777 (.CLK(clknet_leaf_37_clk),
    .D(clknet_1_0__leaf_net702),
    .RESET_B(net698),
    .SCD(net682),
    .SCE(net684),
    .SET_B(net1088),
    .Q(net823),
    .Q_N(net822));
 sky130_fd_sc_hd__sdfrtp_1 merge778 (.CLK(clknet_leaf_39_clk),
    .D(clknet_1_0__leaf_net615),
    .RESET_B(clknet_1_1__leaf_net613),
    .SCD(net1171),
    .SCE(clknet_1_0__leaf_net622),
    .Q(net824));
 sky130_fd_sc_hd__sdfrtp_1 merge779 (.CLK(clknet_leaf_2_clk),
    .D(net267),
    .RESET_B(net1102),
    .SCD(net273),
    .SCE(net281),
    .Q(net825));
 sky130_fd_sc_hd__sdfrtp_1 merge780 (.CLK(clknet_leaf_0_clk),
    .D(net256),
    .RESET_B(net253),
    .SCD(net401),
    .SCE(net1067),
    .Q(net826));
 sky130_fd_sc_hd__clkbuf_1 merge781 (.A(net828),
    .X(net827));
 sky130_fd_sc_hd__dfbbn_1 merge782 (.CLK_N(clknet_leaf_10_clk),
    .D(net20),
    .RESET_B(net19),
    .SET_B(net8),
    .Q(net829),
    .Q_N(net828));
 sky130_fd_sc_hd__sdfbbn_1 merge783 (.CLK_N(clknet_leaf_13_clk),
    .D(net207),
    .RESET_B(net203),
    .SCD(net44),
    .SCE(net43),
    .SET_B(net47),
    .Q(net831),
    .Q_N(net830));
 sky130_fd_sc_hd__mux4_1 merge784 (.A0(net563),
    .A1(net404),
    .A2(net567),
    .A3(clknet_1_0__leaf_net611),
    .S0(clknet_1_0__leaf_net613),
    .S1(net946),
    .X(net832));
 sky130_fd_sc_hd__mux4_1 merge785 (.A0(net1077),
    .A1(net637),
    .A2(clknet_1_0__leaf_net633),
    .A3(net641),
    .S0(net632),
    .S1(clknet_1_0__leaf_net639),
    .X(net833));
 sky130_fd_sc_hd__sdfsbp_1 merge786 (.CLK(clknet_leaf_38_clk),
    .D(clknet_1_0__leaf_net628),
    .SCD(clknet_1_0__leaf_net626),
    .SCE(clknet_1_0__leaf_net725),
    .SET_B(clknet_1_0__leaf_net720),
    .Q(net835),
    .Q_N(net834));
 sky130_fd_sc_hd__sdfbbn_1 merge787 (.CLK_N(clknet_leaf_0_clk),
    .D(net257),
    .RESET_B(net260),
    .SCD(net411),
    .SCE(net408),
    .SET_B(net1067),
    .Q(net837),
    .Q_N(net836));
 sky130_fd_sc_hd__mux4_1 merge788 (.A0(clknet_1_1__leaf_net138),
    .A1(clknet_1_0__leaf_net141),
    .A2(net140),
    .A3(net1069),
    .S0(net404),
    .S1(net296),
    .X(net838));
 sky130_fd_sc_hd__mux4_1 merge789 (.A0(net324),
    .A1(net325),
    .A2(net184),
    .A3(net330),
    .S0(net321),
    .S1(net327),
    .X(net839));
 sky130_fd_sc_hd__sdfsbp_1 merge790 (.CLK(clknet_leaf_22_clk),
    .D(net96),
    .SCD(net94),
    .SCE(net97),
    .SET_B(net1145),
    .Q(net841),
    .Q_N(net840));
 sky130_fd_sc_hd__mux4_1 merge791 (.A0(clknet_1_0__leaf_net451),
    .A1(net449),
    .A2(clknet_1_0__leaf_net139),
    .A3(clknet_1_1__leaf_net138),
    .S0(net140),
    .S1(clknet_1_0__leaf_net911),
    .X(net842));
 sky130_fd_sc_hd__mux4_1 merge792 (.A0(net21),
    .A1(net25),
    .A2(net19),
    .A3(net185),
    .S0(net189),
    .S1(net188),
    .X(net843));
 sky130_fd_sc_hd__mux4_1 merge793 (.A0(net678),
    .A1(net676),
    .A2(net570),
    .A3(net568),
    .S0(net567),
    .S1(net1154),
    .X(net844));
 sky130_fd_sc_hd__mux4_1 merge794 (.A0(net183),
    .A1(net181),
    .A2(net186),
    .A3(net208),
    .S0(net207),
    .S1(net210),
    .X(net845));
 sky130_fd_sc_hd__mux4_1 merge795 (.A0(net430),
    .A1(net433),
    .A2(net1069),
    .A3(clknet_1_1__leaf_net262),
    .S0(net256),
    .S1(net261),
    .X(net846));
 sky130_fd_sc_hd__sdfbbp_1 merge796 (.CLK(clknet_leaf_22_clk),
    .D(net102),
    .RESET_B(net96),
    .SCD(net235),
    .SCE(net238),
    .SET_B(net1104),
    .Q(net848),
    .Q_N(net847));
 sky130_fd_sc_hd__mux4_1 merge797 (.A0(net331),
    .A1(net330),
    .A2(net1073),
    .A3(net49),
    .S0(net44),
    .S1(net1070),
    .X(net849));
 sky130_fd_sc_hd__mux4_1 merge798 (.A0(net227),
    .A1(net168),
    .A2(net169),
    .A3(clknet_1_1__leaf_net167),
    .S0(net922),
    .S1(net946),
    .X(net850));
 sky130_fd_sc_hd__sdfbbn_1 merge799 (.CLK_N(clknet_leaf_29_clk),
    .D(net494),
    .RESET_B(net498),
    .SCD(net496),
    .SET_B(net473),
    .Q(net852),
    .Q_N(net851));
 sky130_fd_sc_hd__mux4_1 merge800 (.A0(net739),
    .A1(clknet_1_0__leaf_net747),
    .A2(net730),
    .A3(net452),
    .S0(clknet_1_1__leaf_net451),
    .S1(clknet_1_0__leaf_net454),
    .X(net853));
 sky130_fd_sc_hd__mux4_1 merge801 (.A0(net627),
    .A1(net618),
    .A2(clknet_1_1__leaf_net622),
    .A3(clknet_1_0__leaf_net756),
    .S0(net757),
    .S1(net753),
    .X(net854));
 sky130_fd_sc_hd__mux4_1 merge802 (.A0(net149),
    .A1(clknet_1_1__leaf_net139),
    .A2(net145),
    .A3(net312),
    .S0(net299),
    .S1(net908),
    .X(net855));
 sky130_fd_sc_hd__sdfbbn_1 merge803 (.CLK_N(clknet_leaf_18_clk),
    .D(net209),
    .RESET_B(net350),
    .SCD(net356),
    .SCE(net348),
    .SET_B(net1096),
    .Q(net857),
    .Q_N(net856));
 sky130_fd_sc_hd__sdfbbp_1 merge804 (.CLK(clknet_leaf_0_clk),
    .D(net1067),
    .RESET_B(net397),
    .SCD(net401),
    .SCE(net1116),
    .SET_B(net1166),
    .Q(net859),
    .Q_N(net858));
 sky130_fd_sc_hd__mux4_1 merge805 (.A0(net678),
    .A1(net677),
    .A2(net680),
    .A3(clknet_1_0__leaf_net720),
    .S0(clknet_1_0__leaf_net722),
    .S1(net996),
    .X(net860));
 sky130_fd_sc_hd__sdfstp_1 merge806 (.CLK(clknet_leaf_28_clk),
    .D(clknet_1_0__leaf_net376),
    .SCE(clknet_1_0__leaf_net377),
    .SET_B(net1113),
    .Q(net861));
 sky130_fd_sc_hd__mux4_1 merge807 (.A0(clknet_1_0__leaf_net518),
    .A1(net473),
    .A2(net500),
    .A3(net499),
    .S0(net927),
    .S1(clknet_1_0__leaf_net948),
    .X(net862));
 sky130_fd_sc_hd__mux4_1 merge808 (.A0(net738),
    .A1(net735),
    .A2(clknet_1_1__leaf_net729),
    .A3(net482),
    .S0(net476),
    .S1(net470),
    .X(net863));
 sky130_fd_sc_hd__mux4_1 merge809 (.A0(net323),
    .A1(net321),
    .A2(net297),
    .A3(net1070),
    .S0(net50),
    .S1(net43),
    .X(net864));
 sky130_fd_sc_hd__dfxbp_1 s810 (.CLK(clknet_leaf_8_clk),
    .D(net10),
    .Q(net865));
 sky130_fd_sc_hd__dfxbp_1 s811 (.CLK(clknet_leaf_8_clk),
    .D(net13),
    .Q(net867),
    .Q_N(net866));
 sky130_fd_sc_hd__dfxtp_1 s812 (.CLK(clknet_leaf_9_clk),
    .D(net15),
    .Q(net868));
 sky130_fd_sc_hd__dfxtp_1 s813 (.CLK(clknet_leaf_9_clk),
    .D(net17),
    .Q(net869));
 sky130_fd_sc_hd__dfxtp_1 s814 (.CLK(clknet_leaf_12_clk),
    .D(net38),
    .Q(net870));
 sky130_fd_sc_hd__dlclkp_1 s815 (.CLK(clknet_leaf_11_clk),
    .GATE(net39),
    .GCLK(net871));
 sky130_fd_sc_hd__dlclkp_2 s816 (.CLK(clknet_leaf_12_clk),
    .GATE(net42),
    .GCLK(net872));
 sky130_fd_sc_hd__dlclkp_4 s817 (.CLK(clknet_leaf_13_clk),
    .GATE(net59),
    .GCLK(net873));
 sky130_fd_sc_hd__dlxbn_1 s818 (.D(net61),
    .GATE_N(clknet_leaf_13_clk),
    .Q(net875),
    .Q_N(net874));
 sky130_fd_sc_hd__dlxbn_1 s819 (.D(net63),
    .GATE_N(clknet_leaf_13_clk),
    .Q(net876));
 sky130_fd_sc_hd__dlxbp_1 s820 (.D(net64),
    .GATE(clknet_leaf_13_clk),
    .Q(net877));
 sky130_fd_sc_hd__dlxtn_1 s821 (.D(net77),
    .GATE_N(clknet_leaf_20_clk),
    .Q(net878));
 sky130_fd_sc_hd__dlxtn_1 s822 (.D(net84),
    .GATE_N(clknet_leaf_21_clk),
    .Q(net879));
 sky130_fd_sc_hd__dlxtn_1 s823 (.D(net87),
    .GATE_N(clknet_leaf_21_clk),
    .Q(net880));
 sky130_fd_sc_hd__dlxtp_1 s824 (.D(net88),
    .GATE(clknet_leaf_21_clk),
    .Q(net881));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s825 (.D(net92),
    .SLEEP_B(clknet_leaf_22_clk),
    .Q(net882));
 sky130_fd_sc_hd__dfxbp_1 s826 (.CLK(clknet_leaf_24_clk),
    .D(net110),
    .Q(net884),
    .Q_N(net883));
 sky130_fd_sc_hd__dfxbp_1 s827 (.CLK(clknet_leaf_24_clk),
    .D(net112),
    .Q(net885));
 sky130_fd_sc_hd__dfxtp_1 s828 (.CLK(clknet_leaf_24_clk),
    .D(net113),
    .Q(net886));
 sky130_fd_sc_hd__dfxtp_1 s829 (.CLK(clknet_leaf_24_clk),
    .D(net1156),
    .Q(net887));
 sky130_fd_sc_hd__dfxtp_1 s830 (.CLK(clknet_leaf_8_clk),
    .D(net129),
    .Q(net888));
 sky130_fd_sc_hd__dlclkp_1 s831 (.CLK(clknet_leaf_7_clk),
    .GATE(net131),
    .GCLK(net889));
 sky130_fd_sc_hd__dlclkp_2 s832 (.CLK(clknet_leaf_1_clk),
    .GATE(net134),
    .GCLK(net890));
 sky130_fd_sc_hd__dlclkp_4 s833 (.CLK(clknet_leaf_7_clk),
    .GATE(net135),
    .GCLK(net891));
 sky130_fd_sc_hd__dlxbn_1 s834 (.D(net158),
    .GATE_N(clknet_leaf_7_clk),
    .Q(net893),
    .Q_N(net892));
 sky130_fd_sc_hd__dlxbn_1 s835 (.D(net174),
    .GATE_N(clknet_leaf_16_clk),
    .Q(net895),
    .Q_N(net894));
 sky130_fd_sc_hd__dlxbp_1 s836 (.D(net178),
    .GATE(clknet_leaf_16_clk),
    .Q(net896));
 sky130_fd_sc_hd__dlxtn_1 s837 (.D(net196),
    .GATE_N(clknet_leaf_14_clk),
    .Q(net897));
 sky130_fd_sc_hd__dlxtn_1 s838 (.D(net198),
    .GATE_N(clknet_leaf_14_clk),
    .Q(net898));
 sky130_fd_sc_hd__dlxtn_1 s839 (.D(net199),
    .GATE_N(clknet_leaf_14_clk),
    .Q(net899));
 sky130_fd_sc_hd__dlxtp_1 s840 (.D(net201),
    .GATE(clknet_leaf_14_clk),
    .Q(net900));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s841 (.D(net202),
    .SLEEP_B(clknet_leaf_14_clk),
    .Q(net901));
 sky130_fd_sc_hd__dfxbp_1 s842 (.CLK(clknet_leaf_19_clk),
    .D(net224),
    .Q(net903),
    .Q_N(net902));
 sky130_fd_sc_hd__dfxbp_1 s843 (.CLK(clknet_leaf_23_clk),
    .D(net246),
    .Q(net905),
    .Q_N(net904));
 sky130_fd_sc_hd__dfxtp_1 s844 (.CLK(clknet_leaf_25_clk),
    .D(net249),
    .Q(net906));
 sky130_fd_sc_hd__dfxtp_1 s845 (.CLK(clknet_leaf_2_clk),
    .D(net265),
    .Q(net907));
 sky130_fd_sc_hd__dfxtp_1 s846 (.CLK(clknet_leaf_6_clk),
    .D(net309),
    .Q(net908));
 sky130_fd_sc_hd__dlclkp_1 s847 (.CLK(clknet_leaf_15_clk),
    .GATE(net314),
    .GCLK(net909));
 sky130_fd_sc_hd__dlclkp_2 s848 (.CLK(clknet_leaf_5_clk),
    .GATE(net317),
    .GCLK(net910));
 sky130_fd_sc_hd__dlclkp_4 s849 (.CLK(clknet_leaf_6_clk),
    .GATE(net320),
    .GCLK(net911));
 sky130_fd_sc_hd__dlxbn_1 s850 (.D(net339),
    .GATE_N(clknet_leaf_18_clk),
    .Q(net913),
    .Q_N(net912));
 sky130_fd_sc_hd__dlxbn_1 s851 (.D(net340),
    .GATE_N(clknet_leaf_18_clk),
    .Q(net915),
    .Q_N(net914));
 sky130_fd_sc_hd__dlxbp_1 s852 (.D(net344),
    .GATE(clknet_leaf_18_clk),
    .Q(net917),
    .Q_N(net916));
 sky130_fd_sc_hd__dlxtn_1 s853 (.D(net345),
    .GATE_N(clknet_leaf_18_clk),
    .Q(net918));
 sky130_fd_sc_hd__dlxtn_1 s854 (.D(net346),
    .GATE_N(clknet_leaf_18_clk),
    .Q(net919));
 sky130_fd_sc_hd__dlxtn_1 s855 (.D(net364),
    .GATE_N(clknet_leaf_28_clk),
    .Q(net920));
 sky130_fd_sc_hd__dlxtp_1 s856 (.D(net369),
    .GATE(clknet_leaf_23_clk),
    .Q(net921));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s857 (.D(net371),
    .SLEEP_B(clknet_leaf_28_clk),
    .Q(net922));
 sky130_fd_sc_hd__dfxbp_1 s858 (.CLK(clknet_leaf_25_clk),
    .D(net389),
    .Q(net924),
    .Q_N(net923));
 sky130_fd_sc_hd__dfxbp_1 s859 (.CLK(clknet_leaf_25_clk),
    .D(net392),
    .Q(net925));
 sky130_fd_sc_hd__dfxtp_1 s860 (.CLK(clknet_leaf_25_clk),
    .D(net393),
    .Q(net926));
 sky130_fd_sc_hd__dfxtp_1 s861 (.CLK(clknet_leaf_26_clk),
    .D(net394),
    .Q(net927));
 sky130_fd_sc_hd__dfxtp_1 s862 (.CLK(clknet_leaf_26_clk),
    .D(net395),
    .Q(net928));
 sky130_fd_sc_hd__dlclkp_1 s863 (.CLK(clknet_leaf_0_clk),
    .GATE(net413),
    .GCLK(net929));
 sky130_fd_sc_hd__dlclkp_2 s864 (.CLK(clknet_leaf_42_clk),
    .GATE(net419),
    .GCLK(net930));
 sky130_fd_sc_hd__dlclkp_4 s865 (.CLK(clknet_leaf_42_clk),
    .GATE(net421),
    .GCLK(net931));
 sky130_fd_sc_hd__dlxbn_1 s866 (.D(net443),
    .GATE_N(clknet_leaf_4_clk),
    .Q(net933),
    .Q_N(net932));
 sky130_fd_sc_hd__dlxbn_1 s867 (.D(net446),
    .GATE_N(clknet_leaf_3_clk),
    .Q(net934));
 sky130_fd_sc_hd__dlxbp_1 s868 (.D(net447),
    .GATE(clknet_leaf_4_clk),
    .Q(net935));
 sky130_fd_sc_hd__dlxtn_1 s869 (.D(net448),
    .GATE_N(clknet_leaf_4_clk),
    .Q(net936));
 sky130_fd_sc_hd__dlxtn_1 s870 (.D(net464),
    .GATE_N(clknet_leaf_4_clk),
    .Q(net937));
 sky130_fd_sc_hd__dlxtn_1 s871 (.D(net466),
    .GATE_N(clknet_leaf_30_clk),
    .Q(net938));
 sky130_fd_sc_hd__dlxtp_1 s872 (.D(net467),
    .GATE(clknet_leaf_40_clk),
    .Q(net939));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s873 (.D(net468),
    .SLEEP_B(clknet_leaf_40_clk),
    .Q(net940));
 sky130_fd_sc_hd__dfxbp_1 s874 (.CLK(clknet_leaf_40_clk),
    .D(net469),
    .Q(net942),
    .Q_N(net941));
 sky130_fd_sc_hd__dfxbp_1 s875 (.CLK(clknet_leaf_29_clk),
    .D(net487),
    .Q(net944),
    .Q_N(net943));
 sky130_fd_sc_hd__dfxtp_1 s876 (.CLK(clknet_leaf_29_clk),
    .D(net488),
    .Q(net945));
 sky130_fd_sc_hd__dfxtp_2 s877 (.CLK(clknet_leaf_29_clk),
    .D(net491),
    .Q(net946));
 sky130_fd_sc_hd__dfxtp_1 s878 (.CLK(clknet_leaf_29_clk),
    .D(net492),
    .Q(net947));
 sky130_fd_sc_hd__dlclkp_1 s879 (.CLK(clknet_leaf_28_clk),
    .GATE(net516),
    .GCLK(net948));
 sky130_fd_sc_hd__dlclkp_2 s880 (.CLK(clknet_leaf_27_clk),
    .GATE(net517),
    .GCLK(net949));
 sky130_fd_sc_hd__dlclkp_4 s881 (.CLK(clknet_leaf_26_clk),
    .GATE(net525),
    .GCLK(net950));
 sky130_fd_sc_hd__dlxbn_1 s882 (.D(net532),
    .GATE_N(clknet_leaf_27_clk),
    .Q(net952),
    .Q_N(net951));
 sky130_fd_sc_hd__dlxbn_1 s883 (.D(net537),
    .GATE_N(clknet_leaf_26_clk),
    .Q(net1063),
    .Q_N(net953));
 sky130_fd_sc_hd__dlxbp_1 s884 (.D(net557),
    .GATE(clknet_leaf_45_clk),
    .Q(net955),
    .Q_N(net954));
 sky130_fd_sc_hd__dlxtn_1 s885 (.D(net561),
    .GATE_N(clknet_leaf_45_clk),
    .Q(net956));
 sky130_fd_sc_hd__dlxtn_2 s886 (.D(net562),
    .GATE_N(clknet_leaf_45_clk),
    .Q(net957));
 sky130_fd_sc_hd__dlxtn_1 s887 (.D(net571),
    .GATE_N(clknet_leaf_42_clk),
    .Q(net958));
 sky130_fd_sc_hd__dlxtp_1 s888 (.D(net578),
    .GATE(clknet_leaf_42_clk),
    .Q(net959));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s889 (.D(net581),
    .SLEEP_B(clknet_leaf_43_clk),
    .Q(net960));
 sky130_fd_sc_hd__dfxbp_1 s890 (.CLK(clknet_leaf_41_clk),
    .D(net582),
    .Q(net962),
    .Q_N(net961));
 sky130_fd_sc_hd__dfxbp_1 s891 (.CLK(clknet_leaf_43_clk),
    .D(net585),
    .Q(net963));
 sky130_fd_sc_hd__dfxtp_1 s892 (.CLK(clknet_leaf_43_clk),
    .D(net586),
    .Q(net964));
 sky130_fd_sc_hd__dfxtp_1 s893 (.CLK(clknet_leaf_39_clk),
    .D(net599),
    .Q(net965));
 sky130_fd_sc_hd__dfxtp_1 s894 (.CLK(clknet_leaf_39_clk),
    .D(net602),
    .Q(net966));
 sky130_fd_sc_hd__dlclkp_1 s895 (.CLK(clknet_leaf_38_clk),
    .GATE(net607),
    .GCLK(net967));
 sky130_fd_sc_hd__dlclkp_2 s896 (.CLK(clknet_leaf_31_clk),
    .GATE(net630),
    .GCLK(net968));
 sky130_fd_sc_hd__dlclkp_4 s897 (.CLK(clknet_leaf_31_clk),
    .GATE(net631),
    .GCLK(net969));
 sky130_fd_sc_hd__dlxbn_1 s898 (.D(net649),
    .GATE_N(clknet_leaf_33_clk),
    .Q(net971),
    .Q_N(net970));
 sky130_fd_sc_hd__dlxbn_1 s899 (.D(net650),
    .GATE_N(clknet_leaf_33_clk),
    .Q(net973),
    .Q_N(net972));
 sky130_fd_sc_hd__dlxbp_1 s900 (.D(net651),
    .GATE(clknet_leaf_33_clk),
    .Q(net974));
 sky130_fd_sc_hd__dlxtn_1 s901 (.D(net652),
    .GATE_N(clknet_leaf_33_clk),
    .Q(net975));
 sky130_fd_sc_hd__dlxtn_1 s902 (.D(net654),
    .GATE_N(clknet_leaf_26_clk),
    .Q(net1056));
 sky130_fd_sc_hd__dlxtn_1 s903 (.D(net665),
    .GATE_N(clknet_leaf_44_clk),
    .Q(net976));
 sky130_fd_sc_hd__dlxtp_1 s904 (.D(net669),
    .GATE(clknet_leaf_44_clk),
    .Q(net977));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s905 (.D(net670),
    .SLEEP_B(clknet_leaf_43_clk),
    .Q(net978));
 sky130_fd_sc_hd__dfxbp_1 s906 (.CLK(clknet_leaf_44_clk),
    .D(net673),
    .Q(net980),
    .Q_N(net979));
 sky130_fd_sc_hd__dfxbp_1 s907 (.CLK(clknet_leaf_43_clk),
    .D(net674),
    .Q(net982),
    .Q_N(net981));
 sky130_fd_sc_hd__dfxtp_1 s908 (.CLK(clknet_leaf_37_clk),
    .D(net692),
    .Q(net983));
 sky130_fd_sc_hd__dfxtp_1 s909 (.CLK(clknet_leaf_37_clk),
    .D(net693),
    .Q(net984));
 sky130_fd_sc_hd__dfxtp_1 s910 (.CLK(clknet_leaf_37_clk),
    .D(net694),
    .Q(net985));
 sky130_fd_sc_hd__dlclkp_1 s911 (.CLK(clknet_leaf_36_clk),
    .GATE(net697),
    .GCLK(net986));
 sky130_fd_sc_hd__dlclkp_2 s912 (.CLK(clknet_leaf_36_clk),
    .GATE(net710),
    .GCLK(net987));
 sky130_fd_sc_hd__dlclkp_4 s913 (.CLK(clknet_leaf_36_clk),
    .GATE(net715),
    .GCLK(net988));
 sky130_fd_sc_hd__dlxbn_1 s914 (.D(net716),
    .GATE_N(clknet_leaf_36_clk),
    .Q(net990),
    .Q_N(net989));
 sky130_fd_sc_hd__dlxbn_1 s915 (.D(net717),
    .GATE_N(clknet_leaf_35_clk),
    .Q(net992),
    .Q_N(net991));
 sky130_fd_sc_hd__dlxbp_1 s916 (.D(net718),
    .GATE(clknet_leaf_38_clk),
    .Q(net994),
    .Q_N(net993));
 sky130_fd_sc_hd__dlxtn_1 s917 (.D(net719),
    .GATE_N(clknet_leaf_35_clk),
    .Q(net995));
 sky130_fd_sc_hd__dlxtn_1 s918 (.D(net721),
    .GATE_N(clknet_leaf_38_clk),
    .Q(net996));
 sky130_fd_sc_hd__dlxtn_1 s919 (.D(net734),
    .GATE_N(clknet_leaf_32_clk),
    .Q(net997));
 sky130_fd_sc_hd__dlxtp_1 s920 (.D(net742),
    .GATE(clknet_leaf_32_clk),
    .Q(net998));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s921 (.D(net743),
    .SLEEP_B(clknet_leaf_32_clk),
    .Q(net999));
 sky130_fd_sc_hd__dfxbp_1 s922 (.CLK(clknet_leaf_38_clk),
    .D(net744),
    .Q(net1001),
    .Q_N(net1000));
 sky130_fd_sc_hd__dfxbp_1 s923 (.CLK(clknet_leaf_35_clk),
    .D(net745),
    .Q(net1002));
 sky130_fd_sc_hd__dfxtp_1 s924 (.CLK(clknet_leaf_35_clk),
    .D(net746),
    .Q(net1003));
 sky130_fd_sc_hd__dfxtp_1 s925 (.CLK(clknet_leaf_34_clk),
    .D(net758),
    .Q(net1004));
 sky130_fd_sc_hd__dfxtp_1 s926 (.CLK(clknet_leaf_33_clk),
    .D(net764),
    .Q(net1005));
 sky130_fd_sc_hd__dlclkp_1 s927 (.CLK(clknet_leaf_34_clk),
    .GATE(net770),
    .GCLK(net1006));
 sky130_fd_sc_hd__dlclkp_2 s928 (.CLK(clknet_leaf_34_clk),
    .GATE(net771),
    .GCLK(net1054));
 sky130_fd_sc_hd__dlclkp_4 s929 (.CLK(clknet_leaf_25_clk),
    .GATE(net797),
    .GCLK(net1007));
 sky130_fd_sc_hd__dlxbn_1 s930 (.D(net816),
    .GATE_N(clknet_leaf_8_clk),
    .Q(net1009),
    .Q_N(net1008));
 sky130_fd_sc_hd__dlxbn_1 s931 (.D(net832),
    .GATE_N(clknet_leaf_40_clk),
    .Q(net1011),
    .Q_N(net1010));
 sky130_fd_sc_hd__dlxbp_1 s932 (.D(net833),
    .GATE(clknet_leaf_27_clk),
    .Q(net1013),
    .Q_N(net1012));
 sky130_fd_sc_hd__dlxtn_1 s933 (.D(net838),
    .GATE_N(clknet_leaf_7_clk),
    .Q(net1014));
 sky130_fd_sc_hd__dlxtn_1 s934 (.D(net839),
    .GATE_N(clknet_leaf_15_clk),
    .Q(net1015));
 sky130_fd_sc_hd__dlxtn_1 s935 (.D(net842),
    .GATE_N(clknet_leaf_7_clk),
    .Q(net1016));
 sky130_fd_sc_hd__dlxtp_1 s936 (.D(net843),
    .GATE(clknet_leaf_12_clk),
    .Q(net1017));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s937 (.D(net844),
    .SLEEP_B(clknet_leaf_43_clk),
    .Q(net1018));
 sky130_fd_sc_hd__dfxbp_1 s938 (.CLK(clknet_leaf_19_clk),
    .D(net845),
    .Q(net1020),
    .Q_N(net1019));
 sky130_fd_sc_hd__dfxbp_1 s939 (.CLK(clknet_leaf_1_clk),
    .D(net846),
    .Q(net1022),
    .Q_N(net1021));
 sky130_fd_sc_hd__dfxtp_1 s940 (.CLK(clknet_leaf_14_clk),
    .D(net849),
    .Q(net1023));
 sky130_fd_sc_hd__dfxtp_1 s941 (.CLK(clknet_leaf_17_clk),
    .D(net850),
    .Q(net1024));
 sky130_fd_sc_hd__dfxtp_1 s942 (.CLK(clknet_leaf_39_clk),
    .D(net853),
    .Q(net1025));
 sky130_fd_sc_hd__dlclkp_1 s943 (.CLK(clknet_leaf_32_clk),
    .GATE(net854),
    .GCLK(net1026));
 sky130_fd_sc_hd__dlclkp_2 s944 (.CLK(clknet_leaf_6_clk),
    .GATE(net855),
    .GCLK(net1027));
 sky130_fd_sc_hd__dlclkp_4 s945 (.CLK(clknet_leaf_38_clk),
    .GATE(net860),
    .GCLK(net1028));
 sky130_fd_sc_hd__dlxbn_1 s946 (.D(net862),
    .GATE_N(clknet_leaf_27_clk),
    .Q(net1030),
    .Q_N(net1029));
 sky130_fd_sc_hd__dlxbn_1 s947 (.D(net863),
    .GATE_N(clknet_leaf_31_clk),
    .Q(net1032),
    .Q_N(net1031));
 sky130_fd_sc_hd__dlxbp_1 s948 (.D(net864),
    .GATE(clknet_leaf_15_clk),
    .Q(net1034),
    .Q_N(net1033));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Right_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Right_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Right_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Right_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Right_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Right_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Right_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Right_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Right_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Right_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Right_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Right_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Right_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Right_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Right_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Right_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Right_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Right_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Right_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Right_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Right_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_161 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_162 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_163 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_164 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_165 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_166 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_167 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_168 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_169 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_170 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_171 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_172 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_173 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_174 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_175 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_176 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_177 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_178 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_179 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_180 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_181 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_182 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Left_183 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Left_184 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Left_185 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Left_186 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Left_187 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Left_188 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Left_189 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Left_190 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Left_191 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Left_192 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Left_193 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Left_194 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Left_195 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Left_196 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Left_197 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Left_198 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Left_199 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Left_200 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Left_201 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Left_202 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Left_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1347 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(in0),
    .X(net773));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(in1),
    .X(net777));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(in10),
    .X(net792));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(in11),
    .X(net801));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(in12),
    .X(net804));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(in13),
    .X(net1035));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(in14),
    .X(net1036));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(in15),
    .X(net1037));
 sky130_fd_sc_hd__buf_1 input9 (.A(in16),
    .X(net1038));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(in17),
    .X(net1039));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(in18),
    .X(net1040));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(in2),
    .X(net1041));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(in20),
    .X(net1042));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(in21),
    .X(net1043));
 sky130_fd_sc_hd__buf_1 input15 (.A(in22),
    .X(net1044));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(in23),
    .X(net1045));
 sky130_fd_sc_hd__dlymetal6s2s_1 input17 (.A(in24),
    .X(net1046));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(in3),
    .X(net1047));
 sky130_fd_sc_hd__clkbuf_1 input19 (.A(in4),
    .X(net1048));
 sky130_fd_sc_hd__clkbuf_1 input20 (.A(in5),
    .X(net1049));
 sky130_fd_sc_hd__clkbuf_1 input21 (.A(in6),
    .X(net1050));
 sky130_fd_sc_hd__clkbuf_1 input22 (.A(in7),
    .X(net1051));
 sky130_fd_sc_hd__clkbuf_1 input23 (.A(in8),
    .X(net1052));
 sky130_fd_sc_hd__clkbuf_1 input24 (.A(in9),
    .X(net1053));
 sky130_fd_sc_hd__clkbuf_1 output25 (.A(net1054),
    .X(out0));
 sky130_fd_sc_hd__buf_8 output26 (.A(clknet_1_1__leaf_net1055),
    .X(out12));
 sky130_fd_sc_hd__buf_2 output27 (.A(net1056),
    .X(out13));
 sky130_fd_sc_hd__clkbuf_1 output28 (.A(clknet_1_0__leaf_net1057),
    .X(out15));
 sky130_fd_sc_hd__buf_2 output29 (.A(net1058),
    .X(out17));
 sky130_fd_sc_hd__buf_2 output30 (.A(net1059),
    .X(out18));
 sky130_fd_sc_hd__buf_2 output31 (.A(net1060),
    .X(out19));
 sky130_fd_sc_hd__buf_2 output32 (.A(net1061),
    .X(out2));
 sky130_fd_sc_hd__buf_2 output33 (.A(net1062),
    .X(out3));
 sky130_fd_sc_hd__buf_2 output34 (.A(net1063),
    .X(out4));
 sky130_fd_sc_hd__buf_2 output35 (.A(net1064),
    .X(out6));
 sky130_fd_sc_hd__buf_2 output36 (.A(net1065),
    .X(out7));
 sky130_fd_sc_hd__buf_2 output37 (.A(net1066),
    .X(out9));
 sky130_fd_sc_hd__buf_2 fanout38 (.A(net402),
    .X(net1067));
 sky130_fd_sc_hd__clkbuf_4 fanout39 (.A(net456),
    .X(net1068));
 sky130_fd_sc_hd__clkbuf_4 fanout40 (.A(net423),
    .X(net1069));
 sky130_fd_sc_hd__buf_2 fanout41 (.A(net47),
    .X(net1070));
 sky130_fd_sc_hd__buf_2 fanout42 (.A(net656),
    .X(net1071));
 sky130_fd_sc_hd__buf_8 fanout43 (.A(net1059),
    .X(net1072));
 sky130_fd_sc_hd__buf_2 fanout44 (.A(net328),
    .X(net1073));
 sky130_fd_sc_hd__buf_2 fanout45 (.A(net183),
    .X(net1074));
 sky130_fd_sc_hd__buf_2 fanout46 (.A(net1076),
    .X(net1075));
 sky130_fd_sc_hd__buf_2 fanout47 (.A(net1077),
    .X(net1076));
 sky130_fd_sc_hd__clkbuf_2 fanout48 (.A(net587),
    .X(net1077));
 sky130_fd_sc_hd__buf_2 fanout49 (.A(net228),
    .X(net1078));
 sky130_fd_sc_hd__buf_2 fanout50 (.A(net470),
    .X(net1079));
 sky130_fd_sc_hd__buf_2 fanout51 (.A(net9),
    .X(net1080));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_0_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_1_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_2_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_3_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_4_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_5_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_6_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_7_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_8_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_9_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_9_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_10_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_11_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_12_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_13_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_14_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_15_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_16_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_17_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_18_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_19_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_20_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_21_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_22_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_22_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_23_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_24_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_24_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_25_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_25_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_26_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_26_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_27_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_27_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_28_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_28_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_29_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_29_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_30_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_30_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_31_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_31_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_32_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_32_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_33_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_33_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_34_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_34_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_35_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_35_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_36_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_36_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_37_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_37_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_38_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_38_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_39_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_39_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_40_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_40_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_41_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_41_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_42_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_42_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_43_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_43_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_44_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_44_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_45_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_45_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net1028 (.A(net1028),
    .X(clknet_0_net1028));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net1028 (.A(clknet_0_net1028),
    .X(clknet_1_0__leaf_net1028));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net1028 (.A(clknet_0_net1028),
    .X(clknet_1_1__leaf_net1028));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net805 (.A(net805),
    .X(clknet_0_net805));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net805 (.A(clknet_0_net805),
    .X(clknet_1_0__leaf_net805));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net805 (.A(clknet_0_net805),
    .X(clknet_1_1__leaf_net805));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net723 (.A(net723),
    .X(clknet_0_net723));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net723 (.A(clknet_0_net723),
    .X(clknet_1_0__leaf_net723));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net723 (.A(clknet_0_net723),
    .X(clknet_1_1__leaf_net723));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net727 (.A(net727),
    .X(clknet_0_net727));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net727 (.A(clknet_0_net727),
    .X(clknet_1_0__leaf_net727));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net727 (.A(clknet_0_net727),
    .X(clknet_1_1__leaf_net727));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net729 (.A(net729),
    .X(clknet_0_net729));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net729 (.A(clknet_0_net729),
    .X(clknet_1_0__leaf_net729));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net729 (.A(clknet_0_net729),
    .X(clknet_1_1__leaf_net729));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net722 (.A(net722),
    .X(clknet_0_net722));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net722 (.A(clknet_0_net722),
    .X(clknet_1_0__leaf_net722));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net722 (.A(clknet_0_net722),
    .X(clknet_1_1__leaf_net722));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net725 (.A(net725),
    .X(clknet_0_net725));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net725 (.A(clknet_0_net725),
    .X(clknet_1_0__leaf_net725));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net725 (.A(clknet_0_net725),
    .X(clknet_1_1__leaf_net725));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net768 (.A(net768),
    .X(clknet_0_net768));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net768 (.A(clknet_0_net768),
    .X(clknet_1_0__leaf_net768));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net768 (.A(clknet_0_net768),
    .X(clknet_1_1__leaf_net768));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net755 (.A(net755),
    .X(clknet_0_net755));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net755 (.A(clknet_0_net755),
    .X(clknet_1_0__leaf_net755));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net755 (.A(clknet_0_net755),
    .X(clknet_1_1__leaf_net755));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net756 (.A(net756),
    .X(clknet_0_net756));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net756 (.A(clknet_0_net756),
    .X(clknet_1_0__leaf_net756));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net756 (.A(clknet_0_net756),
    .X(clknet_1_1__leaf_net756));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net1026 (.A(net1026),
    .X(clknet_0_net1026));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net1026 (.A(clknet_0_net1026),
    .X(clknet_1_0__leaf_net1026));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net1026 (.A(clknet_0_net1026),
    .X(clknet_1_1__leaf_net1026));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net759 (.A(net759),
    .X(clknet_0_net759));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net759 (.A(clknet_0_net759),
    .X(clknet_1_0__leaf_net759));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net759 (.A(clknet_0_net759),
    .X(clknet_1_1__leaf_net759));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net628 (.A(net628),
    .X(clknet_0_net628));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net628 (.A(clknet_0_net628),
    .X(clknet_1_0__leaf_net628));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net628 (.A(clknet_0_net628),
    .X(clknet_1_1__leaf_net628));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net747 (.A(net747),
    .X(clknet_0_net747));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net747 (.A(clknet_0_net747),
    .X(clknet_1_0__leaf_net747));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net747 (.A(clknet_0_net747),
    .X(clknet_1_1__leaf_net747));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net728 (.A(net728),
    .X(clknet_0_net728));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net728 (.A(clknet_0_net728),
    .X(clknet_1_0__leaf_net728));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net728 (.A(clknet_0_net728),
    .X(clknet_1_1__leaf_net728));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net1027 (.A(net1027),
    .X(clknet_0_net1027));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net1027 (.A(clknet_0_net1027),
    .X(clknet_1_0__leaf_net1027));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net1027 (.A(clknet_0_net1027),
    .X(clknet_1_1__leaf_net1027));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net313 (.A(net313),
    .X(clknet_0_net313));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net313 (.A(clknet_0_net313),
    .X(clknet_1_0__leaf_net313));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net313 (.A(clknet_0_net313),
    .X(clknet_1_1__leaf_net313));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net911 (.A(net911),
    .X(clknet_0_net911));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net911 (.A(clknet_0_net911),
    .X(clknet_1_0__leaf_net911));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net911 (.A(clknet_0_net911),
    .X(clknet_1_1__leaf_net911));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net450 (.A(net450),
    .X(clknet_0_net450));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net450 (.A(clknet_0_net450),
    .X(clknet_1_0__leaf_net450));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net450 (.A(clknet_0_net450),
    .X(clknet_1_1__leaf_net450));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net462 (.A(net462),
    .X(clknet_0_net462));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net462 (.A(clknet_0_net462),
    .X(clknet_1_0__leaf_net462));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net462 (.A(clknet_0_net462),
    .X(clknet_1_1__leaf_net462));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net454 (.A(net454),
    .X(clknet_0_net454));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net454 (.A(clknet_0_net454),
    .X(clknet_1_0__leaf_net454));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net454 (.A(clknet_0_net454),
    .X(clknet_1_1__leaf_net454));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net451 (.A(net451),
    .X(clknet_0_net451));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net451 (.A(clknet_0_net451),
    .X(clknet_1_0__leaf_net451));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net451 (.A(clknet_0_net451),
    .X(clknet_1_1__leaf_net451));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net910 (.A(net910),
    .X(clknet_0_net910));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net910 (.A(clknet_0_net910),
    .X(clknet_1_0__leaf_net910));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net910 (.A(clknet_0_net910),
    .X(clknet_1_1__leaf_net910));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net909 (.A(net909),
    .X(clknet_0_net909));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net909 (.A(clknet_0_net909),
    .X(clknet_1_0__leaf_net909));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net909 (.A(clknet_0_net909),
    .X(clknet_1_1__leaf_net909));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net1007 (.A(net1007),
    .X(clknet_0_net1007));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net1007 (.A(clknet_0_net1007),
    .X(clknet_1_0__leaf_net1007));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net1007 (.A(clknet_0_net1007),
    .X(clknet_1_1__leaf_net1007));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net379 (.A(net379),
    .X(clknet_0_net379));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net379 (.A(clknet_0_net379),
    .X(clknet_1_0__leaf_net379));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net379 (.A(clknet_0_net379),
    .X(clknet_1_1__leaf_net379));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net376 (.A(net376),
    .X(clknet_0_net376));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net376 (.A(clknet_0_net376),
    .X(clknet_1_0__leaf_net376));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net376 (.A(clknet_0_net376),
    .X(clknet_1_1__leaf_net376));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net377 (.A(net377),
    .X(clknet_0_net377));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net377 (.A(clknet_0_net377),
    .X(clknet_1_0__leaf_net377));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net377 (.A(clknet_0_net377),
    .X(clknet_1_1__leaf_net377));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net987 (.A(net987),
    .X(clknet_0_net987));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net987 (.A(clknet_0_net987),
    .X(clknet_1_0__leaf_net987));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net987 (.A(clknet_0_net987),
    .X(clknet_1_1__leaf_net987));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net700 (.A(net700),
    .X(clknet_0_net700));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net700 (.A(clknet_0_net700),
    .X(clknet_1_0__leaf_net700));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net700 (.A(clknet_0_net700),
    .X(clknet_1_1__leaf_net700));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net720 (.A(net720),
    .X(clknet_0_net720));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net720 (.A(clknet_0_net720),
    .X(clknet_1_0__leaf_net720));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net720 (.A(clknet_0_net720),
    .X(clknet_1_1__leaf_net720));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net705 (.A(net705),
    .X(clknet_0_net705));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net705 (.A(clknet_0_net705),
    .X(clknet_1_0__leaf_net705));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net705 (.A(clknet_0_net705),
    .X(clknet_1_1__leaf_net705));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net702 (.A(net702),
    .X(clknet_0_net702));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net702 (.A(clknet_0_net702),
    .X(clknet_1_0__leaf_net702));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net702 (.A(clknet_0_net702),
    .X(clknet_1_1__leaf_net702));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net701 (.A(net701),
    .X(clknet_0_net701));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net701 (.A(clknet_0_net701),
    .X(clknet_1_0__leaf_net701));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net701 (.A(clknet_0_net701),
    .X(clknet_1_1__leaf_net701));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net609 (.A(net609),
    .X(clknet_0_net609));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net609 (.A(clknet_0_net609),
    .X(clknet_1_0__leaf_net609));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net609 (.A(clknet_0_net609),
    .X(clknet_1_1__leaf_net609));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net613 (.A(net613),
    .X(clknet_0_net613));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net613 (.A(clknet_0_net613),
    .X(clknet_1_0__leaf_net613));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net613 (.A(clknet_0_net613),
    .X(clknet_1_1__leaf_net613));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net622 (.A(net622),
    .X(clknet_0_net622));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net622 (.A(clknet_0_net622),
    .X(clknet_1_0__leaf_net622));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net622 (.A(clknet_0_net622),
    .X(clknet_1_1__leaf_net622));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net615 (.A(net615),
    .X(clknet_0_net615));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net615 (.A(clknet_0_net615),
    .X(clknet_1_0__leaf_net615));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net615 (.A(clknet_0_net615),
    .X(clknet_1_1__leaf_net615));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net610 (.A(net610),
    .X(clknet_0_net610));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net610 (.A(clknet_0_net610),
    .X(clknet_1_0__leaf_net610));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net610 (.A(clknet_0_net610),
    .X(clknet_1_1__leaf_net610));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net626 (.A(net626),
    .X(clknet_0_net626));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net626 (.A(clknet_0_net626),
    .X(clknet_1_0__leaf_net626));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net626 (.A(clknet_0_net626),
    .X(clknet_1_1__leaf_net626));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net611 (.A(net611),
    .X(clknet_0_net611));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net611 (.A(clknet_0_net611),
    .X(clknet_1_0__leaf_net611));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net611 (.A(clknet_0_net611),
    .X(clknet_1_1__leaf_net611));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net950 (.A(net950),
    .X(clknet_0_net950));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net950 (.A(clknet_0_net950),
    .X(clknet_1_0__leaf_net950));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net950 (.A(clknet_0_net950),
    .X(clknet_1_1__leaf_net950));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net536 (.A(net536),
    .X(clknet_0_net536));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net536 (.A(clknet_0_net536),
    .X(clknet_1_0__leaf_net536));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net536 (.A(clknet_0_net536),
    .X(clknet_1_1__leaf_net536));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net1055 (.A(net1055),
    .X(clknet_0_net1055));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net1055 (.A(clknet_0_net1055),
    .X(clknet_1_0__leaf_net1055));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net1055 (.A(clknet_0_net1055),
    .X(clknet_1_1__leaf_net1055));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net1057 (.A(net1057),
    .X(clknet_0_net1057));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net1057 (.A(clknet_0_net1057),
    .X(clknet_1_0__leaf_net1057));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net1057 (.A(clknet_0_net1057),
    .X(clknet_1_1__leaf_net1057));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net533 (.A(net533),
    .X(clknet_0_net533));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net533 (.A(clknet_0_net533),
    .X(clknet_1_0__leaf_net533));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net533 (.A(clknet_0_net533),
    .X(clknet_1_1__leaf_net533));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net526 (.A(net526),
    .X(clknet_0_net526));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net526 (.A(clknet_0_net526),
    .X(clknet_1_0__leaf_net526));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net526 (.A(clknet_0_net526),
    .X(clknet_1_1__leaf_net526));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net520 (.A(net520),
    .X(clknet_0_net520));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net520 (.A(clknet_0_net520),
    .X(clknet_1_0__leaf_net520));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net520 (.A(clknet_0_net520),
    .X(clknet_1_1__leaf_net520));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net523 (.A(net523),
    .X(clknet_0_net523));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net523 (.A(clknet_0_net523),
    .X(clknet_1_0__leaf_net523));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net523 (.A(clknet_0_net523),
    .X(clknet_1_1__leaf_net523));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net948 (.A(net948),
    .X(clknet_0_net948));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net948 (.A(clknet_0_net948),
    .X(clknet_1_0__leaf_net948));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net948 (.A(clknet_0_net948),
    .X(clknet_1_1__leaf_net948));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net633 (.A(net633),
    .X(clknet_0_net633));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net633 (.A(clknet_0_net633),
    .X(clknet_1_0__leaf_net633));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net633 (.A(clknet_0_net633),
    .X(clknet_1_1__leaf_net633));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net639 (.A(net639),
    .X(clknet_0_net639));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net639 (.A(clknet_0_net639),
    .X(clknet_1_0__leaf_net639));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net639 (.A(clknet_0_net639),
    .X(clknet_1_1__leaf_net639));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net518 (.A(net518),
    .X(clknet_0_net518));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net518 (.A(clknet_0_net518),
    .X(clknet_1_0__leaf_net518));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net518 (.A(clknet_0_net518),
    .X(clknet_1_1__leaf_net518));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net931 (.A(net931),
    .X(clknet_0_net931));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net931 (.A(clknet_0_net931),
    .X(clknet_1_0__leaf_net931));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net931 (.A(clknet_0_net931),
    .X(clknet_1_1__leaf_net931));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net549 (.A(net549),
    .X(clknet_0_net549));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net549 (.A(clknet_0_net549),
    .X(clknet_1_0__leaf_net549));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net549 (.A(clknet_0_net549),
    .X(clknet_1_1__leaf_net549));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net556 (.A(net556),
    .X(clknet_0_net556));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net556 (.A(clknet_0_net556),
    .X(clknet_1_0__leaf_net556));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net556 (.A(clknet_0_net556),
    .X(clknet_1_1__leaf_net556));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net550 (.A(net550),
    .X(clknet_0_net550));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net550 (.A(clknet_0_net550),
    .X(clknet_1_0__leaf_net550));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net550 (.A(clknet_0_net550),
    .X(clknet_1_1__leaf_net550));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net560 (.A(net560),
    .X(clknet_0_net560));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net560 (.A(clknet_0_net560),
    .X(clknet_1_0__leaf_net560));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net560 (.A(clknet_0_net560),
    .X(clknet_1_1__leaf_net560));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net553 (.A(net553),
    .X(clknet_0_net553));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net553 (.A(clknet_0_net553),
    .X(clknet_1_0__leaf_net553));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net553 (.A(clknet_0_net553),
    .X(clknet_1_1__leaf_net553));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net545 (.A(net545),
    .X(clknet_0_net545));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net545 (.A(clknet_0_net545),
    .X(clknet_1_0__leaf_net545));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net545 (.A(clknet_0_net545),
    .X(clknet_1_1__leaf_net545));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net541 (.A(net541),
    .X(clknet_0_net541));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net541 (.A(clknet_0_net541),
    .X(clknet_1_0__leaf_net541));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net541 (.A(clknet_0_net541),
    .X(clknet_1_1__leaf_net541));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net544 (.A(net544),
    .X(clknet_0_net544));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net544 (.A(clknet_0_net544),
    .X(clknet_1_0__leaf_net544));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net544 (.A(clknet_0_net544),
    .X(clknet_1_1__leaf_net544));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net543 (.A(net543),
    .X(clknet_0_net543));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net543 (.A(clknet_0_net543),
    .X(clknet_1_0__leaf_net543));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net543 (.A(clknet_0_net543),
    .X(clknet_1_1__leaf_net543));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net538 (.A(net538),
    .X(clknet_0_net538));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net538 (.A(clknet_0_net538),
    .X(clknet_1_0__leaf_net538));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net538 (.A(clknet_0_net538),
    .X(clknet_1_1__leaf_net538));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net540 (.A(net540),
    .X(clknet_0_net540));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net540 (.A(clknet_0_net540),
    .X(clknet_1_0__leaf_net540));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net540 (.A(clknet_0_net540),
    .X(clknet_1_1__leaf_net540));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net539 (.A(net539),
    .X(clknet_0_net539));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net539 (.A(clknet_0_net539),
    .X(clknet_1_0__leaf_net539));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net539 (.A(clknet_0_net539),
    .X(clknet_1_1__leaf_net539));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net930 (.A(net930),
    .X(clknet_0_net930));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net930 (.A(clknet_0_net930),
    .X(clknet_1_0__leaf_net930));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net930 (.A(clknet_0_net930),
    .X(clknet_1_1__leaf_net930));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net929 (.A(net929),
    .X(clknet_0_net929));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net929 (.A(clknet_0_net929),
    .X(clknet_1_0__leaf_net929));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net929 (.A(clknet_0_net929),
    .X(clknet_1_1__leaf_net929));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net141 (.A(net141),
    .X(clknet_0_net141));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net141 (.A(clknet_0_net141),
    .X(clknet_1_0__leaf_net141));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net141 (.A(clknet_0_net141),
    .X(clknet_1_1__leaf_net141));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net890 (.A(net890),
    .X(clknet_0_net890));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net890 (.A(clknet_0_net890),
    .X(clknet_1_0__leaf_net890));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net890 (.A(clknet_0_net890),
    .X(clknet_1_1__leaf_net890));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net262 (.A(net262),
    .X(clknet_0_net262));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net262 (.A(clknet_0_net262),
    .X(clknet_1_0__leaf_net262));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net262 (.A(clknet_0_net262),
    .X(clknet_1_1__leaf_net262));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net137 (.A(net137),
    .X(clknet_0_net137));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net137 (.A(clknet_0_net137),
    .X(clknet_1_0__leaf_net137));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net137 (.A(clknet_0_net137),
    .X(clknet_1_1__leaf_net137));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net139 (.A(net139),
    .X(clknet_0_net139));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net139 (.A(clknet_0_net139),
    .X(clknet_1_0__leaf_net139));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net139 (.A(clknet_0_net139),
    .X(clknet_1_1__leaf_net139));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net138 (.A(net138),
    .X(clknet_0_net138));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net138 (.A(clknet_0_net138),
    .X(clknet_1_0__leaf_net138));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net138 (.A(clknet_0_net138),
    .X(clknet_1_1__leaf_net138));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net873 (.A(net873),
    .X(clknet_0_net873));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net873 (.A(clknet_0_net873),
    .X(clknet_1_0__leaf_net873));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net873 (.A(clknet_0_net873),
    .X(clknet_1_1__leaf_net873));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net60 (.A(net60),
    .X(clknet_0_net60));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net60 (.A(clknet_0_net60),
    .X(clknet_1_0__leaf_net60));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net60 (.A(clknet_0_net60),
    .X(clknet_1_1__leaf_net60));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net872 (.A(net872),
    .X(clknet_0_net872));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net872 (.A(clknet_0_net872),
    .X(clknet_1_0__leaf_net872));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net872 (.A(clknet_0_net872),
    .X(clknet_1_1__leaf_net872));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net67 (.A(net67),
    .X(clknet_0_net67));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net67 (.A(clknet_0_net67),
    .X(clknet_1_0__leaf_net67));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net67 (.A(clknet_0_net67),
    .X(clknet_1_1__leaf_net67));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net70 (.A(net70),
    .X(clknet_0_net70));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net70 (.A(clknet_0_net70),
    .X(clknet_1_0__leaf_net70));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net70 (.A(clknet_0_net70),
    .X(clknet_1_1__leaf_net70));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net68 (.A(net68),
    .X(clknet_0_net68));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net68 (.A(clknet_0_net68),
    .X(clknet_1_0__leaf_net68));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net68 (.A(clknet_0_net68),
    .X(clknet_1_1__leaf_net68));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net75 (.A(net75),
    .X(clknet_0_net75));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net75 (.A(clknet_0_net75),
    .X(clknet_1_0__leaf_net75));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net75 (.A(clknet_0_net75),
    .X(clknet_1_1__leaf_net75));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net69 (.A(net69),
    .X(clknet_0_net69));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net69 (.A(clknet_0_net69),
    .X(clknet_1_0__leaf_net69));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net69 (.A(clknet_0_net69),
    .X(clknet_1_1__leaf_net69));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net48 (.A(net48),
    .X(clknet_0_net48));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net48 (.A(clknet_0_net48),
    .X(clknet_1_0__leaf_net48));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net48 (.A(clknet_0_net48),
    .X(clknet_1_1__leaf_net48));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net159 (.A(net159),
    .X(clknet_0_net159));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net159 (.A(clknet_0_net159),
    .X(clknet_1_0__leaf_net159));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net159 (.A(clknet_0_net159),
    .X(clknet_1_1__leaf_net159));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net167 (.A(net167),
    .X(clknet_0_net167));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net167 (.A(clknet_0_net167),
    .X(clknet_1_0__leaf_net167));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net167 (.A(clknet_0_net167),
    .X(clknet_1_1__leaf_net167));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net161 (.A(net161),
    .X(clknet_0_net161));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net161 (.A(clknet_0_net161),
    .X(clknet_1_0__leaf_net161));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net161 (.A(clknet_0_net161),
    .X(clknet_1_1__leaf_net161));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net160 (.A(net160),
    .X(clknet_0_net160));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net160 (.A(clknet_0_net160),
    .X(clknet_1_0__leaf_net160));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net160 (.A(clknet_0_net160),
    .X(clknet_1_1__leaf_net160));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net871 (.A(net871),
    .X(clknet_0_net871));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net871 (.A(clknet_0_net871),
    .X(clknet_1_0__leaf_net871));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net871 (.A(clknet_0_net871),
    .X(clknet_1_1__leaf_net871));
 sky130_fd_sc_hd__clkbuf_1 clone1 (.A(net1059),
    .X(net1081));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(net1004),
    .X(net1082));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(net399),
    .X(net1083));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(net411),
    .X(net1084));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(net870),
    .X(net1085));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(net663),
    .X(net1086));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(net896),
    .X(net1087));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(net680),
    .X(net1088));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(net524),
    .X(net1089));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(net877),
    .X(net1090));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(net982),
    .X(net1091));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(net72),
    .X(net1092));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(net275),
    .X(net1093));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(net780),
    .X(net1094));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(net944),
    .X(net1095));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(net914),
    .X(net1096));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(net906),
    .X(net1097));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(net788),
    .X(net1098));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(net569),
    .X(net1099));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(net190),
    .X(net1100));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(net826),
    .X(net1101));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(net264),
    .X(net1102));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(net286),
    .X(net1103));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(net233),
    .X(net1104));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(net351),
    .X(net1105));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(net76),
    .X(net1106));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(net952),
    .X(net1107));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(net187),
    .X(net1108));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(net869),
    .X(net1109));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(net29),
    .X(net1110));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(net761),
    .X(net1111));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(net905),
    .X(net1112));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(net375),
    .X(net1113));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(net310),
    .X(net1114));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(net933),
    .X(net1115));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(net268),
    .X(net1116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(net892),
    .X(net1117));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(net291),
    .X(net1118));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(net937),
    .X(net1119));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(net592),
    .X(net1120));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(net79),
    .X(net1121));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(net207),
    .X(net1122));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(net12),
    .X(net1123));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(net900),
    .X(net1124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(net306),
    .X(net1125));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(net319),
    .X(net1126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(net936),
    .X(net1127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(net740),
    .X(net1128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(net477),
    .X(net1129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(net522),
    .X(net1130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(net432),
    .X(net1131));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(net304),
    .X(net1132));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(net386),
    .X(net1133));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(net938),
    .X(net1134));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(net945),
    .X(net1135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(net552),
    .X(net1136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(net965),
    .X(net1137));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(net35),
    .X(net1138));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(net737),
    .X(net1139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(net959),
    .X(net1140));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(net879),
    .X(net1141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(net865),
    .X(net1142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(net383),
    .X(net1143));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(net926),
    .X(net1144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(net95),
    .X(net1145));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(net963),
    .X(net1146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(net887),
    .X(net1147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(net958),
    .X(net1148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(net868),
    .X(net1149));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(net677),
    .X(net1150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(net907),
    .X(net1151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(net146),
    .X(net1152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(net481),
    .X(net1153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(net957),
    .X(net1154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(net886),
    .X(net1155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(net114),
    .X(net1156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(net527),
    .X(net1157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(net908),
    .X(net1158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(net409),
    .X(net1159));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(net326),
    .X(net1160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(net754),
    .X(net1161));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(net732),
    .X(net1162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(net920),
    .X(net1163));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(net664),
    .X(net1164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(net980),
    .X(net1165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(net404),
    .X(net1166));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(net978),
    .X(net1167));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(net822),
    .X(net1168));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(net486),
    .X(net1169));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(net94),
    .X(net1170));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(net619),
    .X(net1171));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(net323),
    .X(net1172));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(net898),
    .X(net1173));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(net985),
    .X(net1174));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(net217),
    .X(net1175));
 sky130_fd_sc_hd__dlygate4sd3_1 hold96 (.A(net925),
    .X(net1176));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(net327),
    .X(net1177));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(net695),
    .X(net1178));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(net942),
    .X(net1179));
 sky130_fd_sc_hd__dlygate4sd3_1 hold100 (.A(net923),
    .X(net1180));
 sky130_fd_sc_hd__dlygate4sd3_1 hold101 (.A(net289),
    .X(net1181));
 sky130_fd_sc_hd__dlygate4sd3_1 hold102 (.A(net932),
    .X(net1182));
 sky130_fd_sc_hd__dlygate4sd3_1 hold103 (.A(net603),
    .X(net1183));
 sky130_fd_sc_hd__dlygate4sd3_1 hold104 (.A(net752),
    .X(net1184));
 sky130_fd_sc_hd__dlygate4sd3_1 hold105 (.A(net904),
    .X(net1185));
 sky130_fd_sc_hd__dlygate4sd3_1 hold106 (.A(net501),
    .X(net1186));
 sky130_fd_sc_hd__dlygate4sd3_1 hold107 (.A(net352),
    .X(net1187));
 sky130_fd_sc_hd__dlygate4sd3_1 hold108 (.A(net358),
    .X(net1188));
 sky130_fd_sc_hd__dlygate4sd3_1 hold109 (.A(net127),
    .X(net1189));
 sky130_fd_sc_hd__dlygate4sd3_1 hold110 (.A(net667),
    .X(net1190));
 sky130_fd_sc_hd__dlygate4sd3_1 hold111 (.A(net672),
    .X(net1191));
 sky130_fd_sc_hd__dlygate4sd3_1 hold112 (.A(net979),
    .X(net1192));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_A (.DIODE(clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(in0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(in1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(in10));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(in11));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(in12));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(in13));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(in14));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(in15));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(in16));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(in17));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(in18));
 sky130_fd_sc_hd__diode_2 ANTENNA_c252_A (.DIODE(in19));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(in2));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(in20));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(in21));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(in22));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(in23));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(in24));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(in3));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(in4));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(in5));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(in6));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_A (.DIODE(in7));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_A (.DIODE(in8));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_A (.DIODE(in9));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge789_A2 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge776_D (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge744_D (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_SET_B (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_SCE (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_X (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold28_A (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge776_RESET_B (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge740_RESET_B (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_B (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_A (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_A3 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA_c206_A3 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA_c203_S0 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_A2 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_SCD (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_X (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_B (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_B (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_A (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA_c229_Q (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge798_A0 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge759_A2 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge743_RESET_B (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_SCD (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_c230_X (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge788_S1 (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA_c532_A1 (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA_c411_RESET_B (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_A (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_X (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge771_RESET_B (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_S0 (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_A (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_SCD (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_A3 (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_A3 (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_SCD (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_X (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold86_A (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge788_S0 (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge784_A1 (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA_c407_SET_B (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA_c395_SCE (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA_c392_S1 (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA_c385_Q_N (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA_c650_A2 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA_c525_B (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_A (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA_c400_B (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA_c399_B (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA_c394_SCE (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA_c385_Q (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge774_SCE (.DIODE(net589));
 sky130_fd_sc_hd__diode_2 ANTENNA_c566_SCE (.DIODE(net589));
 sky130_fd_sc_hd__diode_2 ANTENNA_c563_DE (.DIODE(net589));
 sky130_fd_sc_hd__diode_2 ANTENNA_c561_SCE (.DIODE(net589));
 sky130_fd_sc_hd__diode_2 ANTENNA_c560_A2 (.DIODE(net589));
 sky130_fd_sc_hd__diode_2 ANTENNA_c557_A2 (.DIODE(net589));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_RESET_B (.DIODE(net589));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_D (.DIODE(net589));
 sky130_fd_sc_hd__diode_2 ANTENNA_c548_X (.DIODE(net589));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge782_SET_B (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c40_A2 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c37_A3 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c33_X (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c26_C (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c25_B (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_C (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout51_A (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c54_SET_B (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c34_X (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_s857_Q (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge798_S0 (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_C1 (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_B (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_s877_Q (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge798_S1 (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge784_S1 (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c571_B (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_D1 (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_B (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_S1 (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold74_A (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_s886_Q (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge754_SCE (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c647_S0 (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c642_D1 (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_SCE (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_B (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_B (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_A (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c534_C (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_s889_Q (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c675_B (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c670_A3 (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c667_S0 (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c656_B (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c549_SET_B (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c542_S1 (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_output29_A (.DIODE(net1058));
 sky130_fd_sc_hd__diode_2 ANTENNA_c373_S0 (.DIODE(net1058));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_A (.DIODE(net1058));
 sky130_fd_sc_hd__diode_2 ANTENNA_c251_A2 (.DIODE(net1058));
 sky130_fd_sc_hd__diode_2 ANTENNA_c250_A1 (.DIODE(net1058));
 sky130_fd_sc_hd__diode_2 ANTENNA_c242_C1 (.DIODE(net1058));
 sky130_fd_sc_hd__diode_2 ANTENNA_c240_X (.DIODE(net1058));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout39_X (.DIODE(net1068));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge740_SCD (.DIODE(net1068));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_S0 (.DIODE(net1068));
 sky130_fd_sc_hd__diode_2 ANTENNA_c437_S0 (.DIODE(net1068));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_SCD (.DIODE(net1068));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_S0 (.DIODE(net1068));
 sky130_fd_sc_hd__diode_2 ANTENNA_c434_B (.DIODE(net1068));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_D_N (.DIODE(net1068));
 sky130_fd_sc_hd__diode_2 ANTENNA_c428_B (.DIODE(net1068));
 sky130_fd_sc_hd__diode_2 ANTENNA_c691_A1 (.DIODE(net1068));
 sky130_fd_sc_hd__diode_2 ANTENNA_c556_B (.DIODE(net1068));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout40_X (.DIODE(net1069));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge740_SCE (.DIODE(net1069));
 sky130_fd_sc_hd__diode_2 ANTENNA_c561_D (.DIODE(net1069));
 sky130_fd_sc_hd__diode_2 ANTENNA_c538_A3 (.DIODE(net1069));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge795_A2 (.DIODE(net1069));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge788_A3 (.DIODE(net1069));
 sky130_fd_sc_hd__diode_2 ANTENNA_c411_SET_B (.DIODE(net1069));
 sky130_fd_sc_hd__diode_2 ANTENNA_c408_SET_B (.DIODE(net1069));
 sky130_fd_sc_hd__diode_2 ANTENNA_c407_SCD (.DIODE(net1069));
 sky130_fd_sc_hd__diode_2 ANTENNA_c403_SCE (.DIODE(net1069));
 sky130_fd_sc_hd__diode_2 ANTENNA_c532_S0 (.DIODE(net1069));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout41_X (.DIODE(net1070));
 sky130_fd_sc_hd__diode_2 ANTENNA_c81_A3 (.DIODE(net1070));
 sky130_fd_sc_hd__diode_2 ANTENNA_c80_D (.DIODE(net1070));
 sky130_fd_sc_hd__diode_2 ANTENNA_c79_S0 (.DIODE(net1070));
 sky130_fd_sc_hd__diode_2 ANTENNA_c78_S0 (.DIODE(net1070));
 sky130_fd_sc_hd__diode_2 ANTENNA_c77_S0 (.DIODE(net1070));
 sky130_fd_sc_hd__diode_2 ANTENNA_c76_D_N (.DIODE(net1070));
 sky130_fd_sc_hd__diode_2 ANTENNA_c70_SET_B (.DIODE(net1070));
 sky130_fd_sc_hd__diode_2 ANTENNA_c68_B (.DIODE(net1070));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge809_A3 (.DIODE(net1070));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge797_S1 (.DIODE(net1070));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout48_X (.DIODE(net1077));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_A2 (.DIODE(net1077));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge785_A0 (.DIODE(net1077));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_A1 (.DIODE(net1077));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_B (.DIODE(net1077));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout47_A (.DIODE(net1077));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout51_X (.DIODE(net1080));
 sky130_fd_sc_hd__diode_2 ANTENNA_c53_B (.DIODE(net1080));
 sky130_fd_sc_hd__diode_2 ANTENNA_c43_B (.DIODE(net1080));
 sky130_fd_sc_hd__diode_2 ANTENNA_c42_A (.DIODE(net1080));
 sky130_fd_sc_hd__diode_2 ANTENNA_c41_A2 (.DIODE(net1080));
 sky130_fd_sc_hd__diode_2 ANTENNA_c38_RESET_B (.DIODE(net1080));
 sky130_fd_sc_hd__diode_2 ANTENNA_c36_SET_B (.DIODE(net1080));
 sky130_fd_sc_hd__diode_2 ANTENNA_c35_A3 (.DIODE(net1080));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_A (.DIODE(net1080));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_A (.DIODE(net1080));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge762_RESET_B (.DIODE(net1080));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_3__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_2__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_1__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_0__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_X (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_45_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_44_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_43_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_42_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_41_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_40_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_4_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_3_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_2_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_1_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_0_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_0__f_clk_X (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_16_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_15_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_14_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_13_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_12_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_11_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_10_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_9_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_8_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_7_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_6_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_5_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_1__f_clk_X (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_39_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_38_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_37_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_36_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_35_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_34_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_33_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_32_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_31_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_30_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_2__f_clk_X (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_29_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_28_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_27_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_26_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_25_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_24_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_23_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_22_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_21_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_20_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_19_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_18_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_17_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_3__f_clk_X (.DIODE(clknet_2_3__leaf_clk));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_441 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_382 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_112 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_543 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_103 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_338 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_525 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_86 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_438 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_411 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_467 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_273 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_368 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_245 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_144 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_160 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_247 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_198 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_16 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_340 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_480 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_486 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_8 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_8 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_20 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_508 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_508 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_228 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_282 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_142 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_413 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_581 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_554 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_32 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_396 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_622 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_245 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_274 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_367 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_567 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_499 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_595 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_553 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_451 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_270 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_226 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_228 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_443 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_617 ();
endmodule
