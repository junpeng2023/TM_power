module netlist_1 (clk,
    in0,
    in1,
    in10,
    in11,
    in12,
    in13,
    in14,
    in15,
    in16,
    in17,
    in18,
    in19,
    in2,
    in20,
    in21,
    in22,
    in23,
    in24,
    in25,
    in26,
    in27,
    in28,
    in29,
    in3,
    in30,
    in31,
    in32,
    in33,
    in34,
    in35,
    in36,
    in37,
    in38,
    in39,
    in4,
    in40,
    in41,
    in42,
    in43,
    in44,
    in45,
    in46,
    in47,
    in48,
    in49,
    in5,
    in50,
    in51,
    in52,
    in53,
    in54,
    in55,
    in56,
    in57,
    in58,
    in59,
    in6,
    in60,
    in61,
    in62,
    in63,
    in64,
    in65,
    in66,
    in67,
    in68,
    in69,
    in7,
    in70,
    in71,
    in72,
    in73,
    in74,
    in75,
    in76,
    in77,
    in78,
    in79,
    in8,
    in80,
    in81,
    in82,
    in83,
    in84,
    in85,
    in86,
    in87,
    in88,
    in89,
    in9,
    in90,
    in91,
    in92,
    in93,
    in94,
    in95,
    in96,
    in97,
    in98,
    in99,
    out0,
    out1,
    out10,
    out11,
    out12,
    out13,
    out14,
    out15,
    out16,
    out17,
    out18,
    out19,
    out2,
    out20,
    out21,
    out22,
    out23,
    out24,
    out25,
    out26,
    out27,
    out28,
    out29,
    out3,
    out30,
    out31,
    out32,
    out33,
    out34,
    out35,
    out36,
    out37,
    out38,
    out39,
    out4,
    out40,
    out41,
    out42,
    out43,
    out44,
    out45,
    out46,
    out47,
    out48,
    out49,
    out5,
    out50,
    out51,
    out52,
    out53,
    out54,
    out55,
    out56,
    out57,
    out58,
    out59,
    out6,
    out60,
    out61,
    out62,
    out63,
    out64,
    out65,
    out66,
    out67,
    out68,
    out69,
    out7,
    out70,
    out71,
    out72,
    out73,
    out74,
    out75,
    out76,
    out77,
    out78,
    out79,
    out8,
    out80,
    out81,
    out82,
    out83,
    out84,
    out85,
    out86,
    out87,
    out88,
    out89,
    out9,
    out90,
    out91,
    out92,
    out93,
    out94,
    out95,
    out96,
    out97,
    out98,
    out99,
    rst);
 input clk;
 input in0;
 input in1;
 input in10;
 input in11;
 input in12;
 input in13;
 input in14;
 input in15;
 input in16;
 input in17;
 input in18;
 input in19;
 input in2;
 input in20;
 input in21;
 input in22;
 input in23;
 input in24;
 input in25;
 input in26;
 input in27;
 input in28;
 input in29;
 input in3;
 input in30;
 input in31;
 input in32;
 input in33;
 input in34;
 input in35;
 input in36;
 input in37;
 input in38;
 input in39;
 input in4;
 input in40;
 input in41;
 input in42;
 input in43;
 input in44;
 input in45;
 input in46;
 input in47;
 input in48;
 input in49;
 input in5;
 input in50;
 input in51;
 input in52;
 input in53;
 input in54;
 input in55;
 input in56;
 input in57;
 input in58;
 input in59;
 input in6;
 input in60;
 input in61;
 input in62;
 input in63;
 input in64;
 input in65;
 input in66;
 input in67;
 input in68;
 input in69;
 input in7;
 input in70;
 input in71;
 input in72;
 input in73;
 input in74;
 input in75;
 input in76;
 input in77;
 input in78;
 input in79;
 input in8;
 input in80;
 input in81;
 input in82;
 input in83;
 input in84;
 input in85;
 input in86;
 input in87;
 input in88;
 input in89;
 input in9;
 input in90;
 input in91;
 input in92;
 input in93;
 input in94;
 input in95;
 input in96;
 input in97;
 input in98;
 input in99;
 output out0;
 output out1;
 output out10;
 output out11;
 output out12;
 output out13;
 output out14;
 output out15;
 output out16;
 output out17;
 output out18;
 output out19;
 output out2;
 output out20;
 output out21;
 output out22;
 output out23;
 output out24;
 output out25;
 output out26;
 output out27;
 output out28;
 output out29;
 output out3;
 output out30;
 output out31;
 output out32;
 output out33;
 output out34;
 output out35;
 output out36;
 output out37;
 output out38;
 output out39;
 output out4;
 output out40;
 output out41;
 output out42;
 output out43;
 output out44;
 output out45;
 output out46;
 output out47;
 output out48;
 output out49;
 output out5;
 output out50;
 output out51;
 output out52;
 output out53;
 output out54;
 output out55;
 output out56;
 output out57;
 output out58;
 output out59;
 output out6;
 output out60;
 output out61;
 output out62;
 output out63;
 output out64;
 output out65;
 output out66;
 output out67;
 output out68;
 output out69;
 output out7;
 output out70;
 output out71;
 output out72;
 output out73;
 output out74;
 output out75;
 output out76;
 output out77;
 output out78;
 output out79;
 output out8;
 output out80;
 output out81;
 output out82;
 output out83;
 output out84;
 output out85;
 output out86;
 output out87;
 output out88;
 output out89;
 output out9;
 output out90;
 output out91;
 output out92;
 output out93;
 output out94;
 output out95;
 output out96;
 output out97;
 output out98;
 output out99;
 input rst;

 wire clknet_0_clk;
 wire clknet_0_net506;
 wire clknet_0_net561;
 wire clknet_0_net562;
 wire clknet_0_net563;
 wire clknet_1_0__leaf_net506;
 wire clknet_1_0__leaf_net561;
 wire clknet_1_0__leaf_net562;
 wire clknet_1_0__leaf_net563;
 wire clknet_1_1__leaf_net506;
 wire clknet_1_1__leaf_net561;
 wire clknet_1_1__leaf_net562;
 wire clknet_1_1__leaf_net563;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire net0;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net63;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net64;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net65;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net66;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net67;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net68;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net69;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net7;
 wire net70;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net71;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net72;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net73;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net74;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net75;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net76;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net77;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net78;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net79;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net8;
 wire net80;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net81;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net82;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net83;
 wire net830;
 wire net831;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;

 sky130_fd_sc_hd__diode_2 ANTENNA_c100_A3 (.DIODE(net1089));
 sky130_fd_sc_hd__diode_2 ANTENNA_c100_B1 (.DIODE(net1094));
 sky130_fd_sc_hd__diode_2 ANTENNA_c100_X (.DIODE(net688));
 sky130_fd_sc_hd__diode_2 ANTENNA_c102_A1 (.DIODE(net604));
 sky130_fd_sc_hd__diode_2 ANTENNA_c102_A2 (.DIODE(net659));
 sky130_fd_sc_hd__diode_2 ANTENNA_c102_B1_N (.DIODE(net1114));
 sky130_fd_sc_hd__diode_2 ANTENNA_c102_X (.DIODE(net735));
 sky130_fd_sc_hd__diode_2 ANTENNA_c103_A (.DIODE(net615));
 sky130_fd_sc_hd__diode_2 ANTENNA_c103_B (.DIODE(net658));
 sky130_fd_sc_hd__diode_2 ANTENNA_c104_A1 (.DIODE(net1083));
 sky130_fd_sc_hd__diode_2 ANTENNA_c104_A3 (.DIODE(net615));
 sky130_fd_sc_hd__diode_2 ANTENNA_c104_S0 (.DIODE(net659));
 sky130_fd_sc_hd__diode_2 ANTENNA_c104_S1 (.DIODE(net1089));
 sky130_fd_sc_hd__diode_2 ANTENNA_c105_A1 (.DIODE(net1094));
 sky130_fd_sc_hd__diode_2 ANTENNA_c105_A2 (.DIODE(net1103));
 sky130_fd_sc_hd__diode_2 ANTENNA_c105_B1_N (.DIODE(net1100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c106_A (.DIODE(net735));
 sky130_fd_sc_hd__diode_2 ANTENNA_c106_B (.DIODE(net601));
 sky130_fd_sc_hd__diode_2 ANTENNA_c107_B (.DIODE(net735));
 sky130_fd_sc_hd__diode_2 ANTENNA_c108_B (.DIODE(net607));
 sky130_fd_sc_hd__diode_2 ANTENNA_c109_S0 (.DIODE(net663));
 sky130_fd_sc_hd__diode_2 ANTENNA_c109_S1 (.DIODE(net1094));
 sky130_fd_sc_hd__diode_2 ANTENNA_c109_X (.DIODE(net722));
 sky130_fd_sc_hd__diode_2 ANTENNA_c110_A (.DIODE(net1108));
 sky130_fd_sc_hd__diode_2 ANTENNA_c110_B (.DIODE(net603));
 sky130_fd_sc_hd__diode_2 ANTENNA_c111_B (.DIODE(net623));
 sky130_fd_sc_hd__diode_2 ANTENNA_c112_A (.DIODE(net1114));
 sky130_fd_sc_hd__diode_2 ANTENNA_c113_A (.DIODE(net595));
 sky130_fd_sc_hd__diode_2 ANTENNA_c113_B (.DIODE(net623));
 sky130_fd_sc_hd__diode_2 ANTENNA_c114_A (.DIODE(net587));
 sky130_fd_sc_hd__diode_2 ANTENNA_c114_B (.DIODE(net722));
 sky130_fd_sc_hd__diode_2 ANTENNA_c115_B (.DIODE(net620));
 sky130_fd_sc_hd__diode_2 ANTENNA_c116_A (.DIODE(net1100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c116_Y (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_c119_B (.DIODE(net645));
 sky130_fd_sc_hd__diode_2 ANTENNA_c122_A (.DIODE(net620));
 sky130_fd_sc_hd__diode_2 ANTENNA_c125_B (.DIODE(net595));
 sky130_fd_sc_hd__diode_2 ANTENNA_c127_B (.DIODE(net1094));
 sky130_fd_sc_hd__diode_2 ANTENNA_c127_Y (.DIODE(net693));
 sky130_fd_sc_hd__diode_2 ANTENNA_c128_A2 (.DIODE(net693));
 sky130_fd_sc_hd__diode_2 ANTENNA_c129_A (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_c131_A2 (.DIODE(net603));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_A (.DIODE(net633));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_B (.DIODE(net1096));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_A (.DIODE(net1143));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_B (.DIODE(net1151));
 sky130_fd_sc_hd__diode_2 ANTENNA_c134_A (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_c134_B (.DIODE(net1100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_A (.DIODE(net1143));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_B (.DIODE(net1108));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_Y (.DIODE(net1093));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_B (.DIODE(net1097));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_Y (.DIODE(net1078));
 sky130_fd_sc_hd__diode_2 ANTENNA_c138_A2 (.DIODE(net1078));
 sky130_fd_sc_hd__diode_2 ANTENNA_c138_B1_N (.DIODE(net1101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c138_X (.DIODE(net1067));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_B (.DIODE(net570));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_Y (.DIODE(net1076));
 sky130_fd_sc_hd__diode_2 ANTENNA_c140_B (.DIODE(net1119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_A (.DIODE(net570));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_B (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_Y (.DIODE(net1156));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_A1 (.DIODE(net1093));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_A2 (.DIODE(net1100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_X (.DIODE(net1063));
 sky130_fd_sc_hd__diode_2 ANTENNA_c143_A (.DIODE(net1096));
 sky130_fd_sc_hd__diode_2 ANTENNA_c143_B (.DIODE(net759));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_A1 (.DIODE(net577));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_A2 (.DIODE(net1097));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_X (.DIODE(net1162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_B (.DIODE(net577));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_A0 (.DIODE(net1076));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_A1 (.DIODE(net1119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_A3 (.DIODE(net1099));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_S0 (.DIODE(net1093));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_X (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_A (.DIODE(net1063));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_A2 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_X (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_A1 (.DIODE(net1162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_A3 (.DIODE(net759));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_X (.DIODE(net1054));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_A1 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_A2 (.DIODE(net1054));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_X (.DIODE(net1053));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_A2 (.DIODE(net1099));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_X (.DIODE(net1057));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_A0 (.DIODE(net1053));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_A1 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_A2 (.DIODE(net1162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_A3 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_S0 (.DIODE(net1057));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_X (.DIODE(net1049));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_A (.DIODE(net603));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_B (.DIODE(net1114));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_Y (.DIODE(net1092));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_A (.DIODE(net593));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_B (.DIODE(net577));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_A (.DIODE(net577));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_B (.DIODE(net1117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_A1 (.DIODE(net582));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_A2 (.DIODE(net1100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_A3 (.DIODE(net597));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_B1 (.DIODE(net1084));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_X (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_c158_B (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_c158_Y (.DIODE(net724));
 sky130_fd_sc_hd__diode_2 ANTENNA_c159_B (.DIODE(net1084));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_A (.DIODE(net1097));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_B (.DIODE(net1084));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_Y (.DIODE(net1074));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_A (.DIODE(net1107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_B (.DIODE(net1114));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_Y (.DIODE(net1065));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_B (.DIODE(net519));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_Y (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_A (.DIODE(net584));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_B (.DIODE(net583));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_A0 (.DIODE(net724));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_A1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_S0 (.DIODE(net1084));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_S1 (.DIODE(net1108));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_A1 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_A2 (.DIODE(net604));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_B1_N (.DIODE(net1084));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_X (.DIODE(net1069));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_A3 (.DIODE(net1084));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_B1 (.DIODE(net1092));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_A (.DIODE(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_Y (.DIODE(net1088));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_A1 (.DIODE(net1092));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_A2 (.DIODE(net604));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_X (.DIODE(net1062));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_A1 (.DIODE(net1069));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_A2 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_A1 (.DIODE(net1092));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_B1_N (.DIODE(net1062));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_X (.DIODE(net1059));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_X (.DIODE(net1052));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_A1 (.DIODE(net1052));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_A2 (.DIODE(net1116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_A3 (.DIODE(net593));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_B1 (.DIODE(net1059));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_A2 (.DIODE(net1065));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_B1_N (.DIODE(net1052));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_A2 (.DIODE(net1052));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_A (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_B (.DIODE(net620));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_B (.DIODE(net633));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_A1 (.DIODE(net620));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_A2 (.DIODE(net627));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_B1_N (.DIODE(net1059));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_X (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_A (.DIODE(net1143));
 sky130_fd_sc_hd__diode_2 ANTENNA_c180_A2 (.DIODE(net1067));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_Y (.DIODE(net673));
 sky130_fd_sc_hd__diode_2 ANTENNA_c182_B (.DIODE(net673));
 sky130_fd_sc_hd__diode_2 ANTENNA_c182_Y (.DIODE(net1073));
 sky130_fd_sc_hd__diode_2 ANTENNA_c184_B (.DIODE(net1162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_A1 (.DIODE(net1093));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_B1_N (.DIODE(net583));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_X (.DIODE(net1087));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_B1_N (.DIODE(net1073));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_A2 (.DIODE(net1073));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_B1_N (.DIODE(net1087));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_X (.DIODE(net1056));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_A (.DIODE(net1073));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_B (.DIODE(net1117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_A1 (.DIODE(net1162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_A3 (.DIODE(net1056));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_B1 (.DIODE(net1107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c190_A2 (.DIODE(net615));
 sky130_fd_sc_hd__diode_2 ANTENNA_c190_B1_N (.DIODE(net1087));
 sky130_fd_sc_hd__diode_2 ANTENNA_c190_X (.DIODE(net1072));
 sky130_fd_sc_hd__diode_2 ANTENNA_c191_Y (.DIODE(net1163));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_A1 (.DIODE(net1087));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_A2 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_B1_N (.DIODE(net1084));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_X (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_A1 (.DIODE(net1163));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_A3 (.DIODE(net1117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_S1 (.DIODE(net1084));
 sky130_fd_sc_hd__diode_2 ANTENNA_c194_A2 (.DIODE(net1073));
 sky130_fd_sc_hd__diode_2 ANTENNA_c194_B1_N (.DIODE(net1056));
 sky130_fd_sc_hd__diode_2 ANTENNA_c194_X (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_A2 (.DIODE(net1072));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_A1 (.DIODE(net1056));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_B1 (.DIODE(net1105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_A2 (.DIODE(net1088));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_A3 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA_c198_B (.DIODE(net1121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_B (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_A2 (.DIODE(net1107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_X (.DIODE(net1048));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_A (.DIODE(net1048));
 sky130_fd_sc_hd__diode_2 ANTENNA_c203_A (.DIODE(net1163));
 sky130_fd_sc_hd__diode_2 ANTENNA_c205_B (.DIODE(net724));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_B (.DIODE(net1073));
 sky130_fd_sc_hd__diode_2 ANTENNA_c208_A2 (.DIODE(net636));
 sky130_fd_sc_hd__diode_2 ANTENNA_c208_B1_N (.DIODE(net1117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_B (.DIODE(net581));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_Y (.DIODE(net706));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_A3 (.DIODE(net1087));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_A2 (.DIODE(net1048));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_S0 (.DIODE(net650));
 sky130_fd_sc_hd__diode_2 ANTENNA_c215_B (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_B (.DIODE(net1048));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_X (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_c220_A3 (.DIODE(net659));
 sky130_fd_sc_hd__diode_2 ANTENNA_c220_X (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA_c221_A3 (.DIODE(net735));
 sky130_fd_sc_hd__diode_2 ANTENNA_c222_B (.DIODE(net595));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_A2 (.DIODE(net1083));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_B1_N (.DIODE(net1117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_B (.DIODE(net1083));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_A (.DIODE(net1055));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_B (.DIODE(net660));
 sky130_fd_sc_hd__diode_2 ANTENNA_c226_Y (.DIODE(net669));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_B (.DIODE(net1076));
 sky130_fd_sc_hd__diode_2 ANTENNA_c229_B1_N (.DIODE(net1048));
 sky130_fd_sc_hd__diode_2 ANTENNA_c229_X (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA_c232_B1_N (.DIODE(net1054));
 sky130_fd_sc_hd__diode_2 ANTENNA_c232_X (.DIODE(net696));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_A (.DIODE(net1121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_B (.DIODE(net669));
 sky130_fd_sc_hd__diode_2 ANTENNA_c234_Y (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA_c235_A (.DIODE(net659));
 sky130_fd_sc_hd__diode_2 ANTENNA_c235_B (.DIODE(net1123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c236_X (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_c237_Y (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_c239_A0 (.DIODE(net1057));
 sky130_fd_sc_hd__diode_2 ANTENNA_c239_S0 (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_c240_B1_N (.DIODE(net1087));
 sky130_fd_sc_hd__diode_2 ANTENNA_c241_B1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA_c264_A (.DIODE(net1097));
 sky130_fd_sc_hd__diode_2 ANTENNA_c264_B (.DIODE(net570));
 sky130_fd_sc_hd__diode_2 ANTENNA_c265_A (.DIODE(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA_c265_Y (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA_c266_A (.DIODE(net1099));
 sky130_fd_sc_hd__diode_2 ANTENNA_c266_B (.DIODE(net1116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c267_A1 (.DIODE(net1096));
 sky130_fd_sc_hd__diode_2 ANTENNA_c267_A2 (.DIODE(net1101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c267_X (.DIODE(net1071));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_A (.DIODE(net1099));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_B (.DIODE(net1067));
 sky130_fd_sc_hd__diode_2 ANTENNA_c272_A (.DIODE(net1095));
 sky130_fd_sc_hd__diode_2 ANTENNA_c272_B (.DIODE(net1097));
 sky130_fd_sc_hd__diode_2 ANTENNA_c272_Y (.DIODE(net1091));
 sky130_fd_sc_hd__diode_2 ANTENNA_c273_Y (.DIODE(net1159));
 sky130_fd_sc_hd__diode_2 ANTENNA_c274_Y (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c275_A (.DIODE(net1091));
 sky130_fd_sc_hd__diode_2 ANTENNA_c276_A (.DIODE(net1071));
 sky130_fd_sc_hd__diode_2 ANTENNA_c276_B (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_c276_Y (.DIODE(net1068));
 sky130_fd_sc_hd__diode_2 ANTENNA_c278_B (.DIODE(net1159));
 sky130_fd_sc_hd__diode_2 ANTENNA_c278_Y (.DIODE(net1046));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_A2 (.DIODE(net1159));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_X (.DIODE(net1044));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_A (.DIODE(net1098));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_Y (.DIODE(net1043));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_B (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA_c283_Y (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_B1_N (.DIODE(net1046));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_X (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_A1 (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_A2 (.DIODE(net1046));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_A3 (.DIODE(net1044));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_A4 (.DIODE(net1076));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_X (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c286_A (.DIODE(net1052));
 sky130_fd_sc_hd__diode_2 ANTENNA_c286_B (.DIODE(net519));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_A (.DIODE(net1084));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_Y (.DIODE(net689));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_A (.DIODE(net689));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_A (.DIODE(net601));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_Y (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_Y (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_B (.DIODE(net599));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_A2 (.DIODE(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_B1_N (.DIODE(net1114));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_A (.DIODE(net599));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_B (.DIODE(net1159));
 sky130_fd_sc_hd__diode_2 ANTENNA_c295_A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c295_Y (.DIODE(net1050));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_A1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_A2 (.DIODE(net1050));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_B1_N (.DIODE(net1034));
 sky130_fd_sc_hd__diode_2 ANTENNA_c297_A1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_Y (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_A2 (.DIODE(net586));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_X (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_A2 (.DIODE(net584));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_A3 (.DIODE(net1091));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_B1 (.DIODE(net1034));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_A (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_B (.DIODE(net1067));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_A2 (.DIODE(net593));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_B1_N (.DIODE(net582));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_A2 (.DIODE(net1050));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_B1_N (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_Y (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_A0 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_A1 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_S0 (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_S1 (.DIODE(net1034));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_A0 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_A3 (.DIODE(net1034));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_S0 (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_S1 (.DIODE(net1084));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_B (.DIODE(net613));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_Y (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_A2 (.DIODE(net1122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_B1_N (.DIODE(net1078));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_B (.DIODE(net1103));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_A (.DIODE(net627));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_B (.DIODE(net623));
 sky130_fd_sc_hd__diode_2 ANTENNA_c313_B (.DIODE(net1043));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_A (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_A2 (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_B1_N (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_Y (.DIODE(net1036));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_B (.DIODE(net1111));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_A1 (.DIODE(net599));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_B1_N (.DIODE(net1050));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_A1 (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_A2 (.DIODE(net623));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_B1_N (.DIODE(net1088));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_X (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c321_A2 (.DIODE(net607));
 sky130_fd_sc_hd__diode_2 ANTENNA_c321_B1_N (.DIODE(net673));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_A (.DIODE(net1116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_B (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_A1 (.DIODE(net1067));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_A2 (.DIODE(net1062));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_B1_N (.DIODE(net1036));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_A (.DIODE(net602));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_B (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_A1 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_A2 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_A2 (.DIODE(net1114));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_A3 (.DIODE(net599));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_S0 (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_S1 (.DIODE(net621));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_B1_N (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_A3 (.DIODE(net1088));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_B1 (.DIODE(net1089));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_X (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_A1 (.DIODE(net1073));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_A2 (.DIODE(net1163));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_B1_N (.DIODE(net1036));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_A1 (.DIODE(net583));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_A3 (.DIODE(net1144));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_A4 (.DIODE(net1089));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_B1 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_A2 (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_X (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_A2 (.DIODE(net1036));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_A3 (.DIODE(net1049));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_B1 (.DIODE(net1034));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_A2 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_c340_A2 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c340_B1_N (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_A (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_B (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_B1_N (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_X (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_A1 (.DIODE(net1043));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_B1_N (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c344_B1_N (.DIODE(net641));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_A3 (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_A4 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_B1 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_X (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_B1_N (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_X (.DIODE(net720));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_A (.DIODE(net1082));
 sky130_fd_sc_hd__diode_2 ANTENNA_c350_A (.DIODE(net1082));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_A1 (.DIODE(net1088));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_A3 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_S1 (.DIODE(net1034));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_A3 (.DIODE(net722));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_B1 (.DIODE(net696));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_A2 (.DIODE(net720));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_B1_N (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_A2 (.DIODE(net632));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_A2 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_B1_N (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_A (.DIODE(net621));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_B (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_B1_N (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_A1 (.DIODE(net1057));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_A2 (.DIODE(net650));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_A3 (.DIODE(net1119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_S0 (.DIODE(net1096));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_S1 (.DIODE(net1083));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_A1 (.DIODE(net654));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_A1 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_A2 (.DIODE(net621));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_A1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_A2 (.DIODE(net654));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_A1 (.DIODE(net575));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_S0 (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_S1 (.DIODE(net1089));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_X (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_A1 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_A2 (.DIODE(net1089));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_A3 (.DIODE(net650));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_S0 (.DIODE(net1048));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_X (.DIODE(net705));
 sky130_fd_sc_hd__diode_2 ANTENNA_c364_A3 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c364_A4 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c364_B1 (.DIODE(net706));
 sky130_fd_sc_hd__diode_2 ANTENNA_c365_B1_N (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA_c366_A (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_A2 (.DIODE(net1076));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_B1_N (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_c368_B1_N (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c369_X (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA_c371_A (.DIODE(net1082));
 sky130_fd_sc_hd__diode_2 ANTENNA_c373_A1 (.DIODE(net1117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c373_A3 (.DIODE(net1163));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_B (.DIODE(net1121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c397_A (.DIODE(net1099));
 sky130_fd_sc_hd__diode_2 ANTENNA_c397_B (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA_c398_B1_N (.DIODE(net1093));
 sky130_fd_sc_hd__diode_2 ANTENNA_c398_X (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_c399_A (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_c399_B (.DIODE(net1098));
 sky130_fd_sc_hd__diode_2 ANTENNA_c400_B (.DIODE(net1071));
 sky130_fd_sc_hd__diode_2 ANTENNA_c401_A (.DIODE(net1123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c401_B (.DIODE(net1063));
 sky130_fd_sc_hd__diode_2 ANTENNA_c401_Y (.DIODE(net1058));
 sky130_fd_sc_hd__diode_2 ANTENNA_c403_Y (.DIODE(net1127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c404_B (.DIODE(net1068));
 sky130_fd_sc_hd__diode_2 ANTENNA_c404_Y (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA_c405_A (.DIODE(net519));
 sky130_fd_sc_hd__diode_2 ANTENNA_c405_B (.DIODE(net1123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c405_Y (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA_c406_A1 (.DIODE(net1044));
 sky130_fd_sc_hd__diode_2 ANTENNA_c407_Y (.DIODE(net686));
 sky130_fd_sc_hd__diode_2 ANTENNA_c408_A (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_c409_A (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA_c409_Y (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_c410_A (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_c410_Y (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA_c411_B (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA_c412_B (.DIODE(net1095));
 sky130_fd_sc_hd__diode_2 ANTENNA_c412_Y (.DIODE(net692));
 sky130_fd_sc_hd__diode_2 ANTENNA_c413_A (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_c413_B (.DIODE(net1099));
 sky130_fd_sc_hd__diode_2 ANTENNA_c414_Y (.DIODE(net674));
 sky130_fd_sc_hd__diode_2 ANTENNA_c415_A (.DIODE(net1127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c416_B (.DIODE(net1043));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_A3 (.DIODE(net692));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_A4 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_B (.DIODE(net759));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_Y (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_A (.DIODE(net1093));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_B (.DIODE(net1127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_A (.DIODE(net1067));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_B (.DIODE(net1091));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_A1 (.DIODE(net1068));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_A3 (.DIODE(net1071));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_B1 (.DIODE(net1144));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_A2 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_A3 (.DIODE(net1063));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_B1 (.DIODE(net1074));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_B (.DIODE(net1092));
 sky130_fd_sc_hd__diode_2 ANTENNA_c424_A (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_A1 (.DIODE(net1107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_X (.DIODE(net679));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_A1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_A3 (.DIODE(net679));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_B1 (.DIODE(net1144));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_X (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA_c427_B1_N (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c427_X (.DIODE(net1148));
 sky130_fd_sc_hd__diode_2 ANTENNA_c428_Y (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_Y (.DIODE(net1028));
 sky130_fd_sc_hd__diode_2 ANTENNA_c430_B1_N (.DIODE(net1068));
 sky130_fd_sc_hd__diode_2 ANTENNA_c430_X (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c431_A1 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA_c431_A2 (.DIODE(net1127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c431_B1_N (.DIODE(net1028));
 sky130_fd_sc_hd__diode_2 ANTENNA_c431_X (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_A2 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_B1_N (.DIODE(net689));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_X (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_A0 (.DIODE(net1148));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_A1 (.DIODE(net1028));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_A3 (.DIODE(net1114));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_S0 (.DIODE(net1098));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_S1 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA_c434_A (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_Y (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_A (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c437_A (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_A (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_A (.DIODE(net1028));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_B (.DIODE(net679));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_A (.DIODE(net1112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_A2 (.DIODE(net1046));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_B1_N (.DIODE(net1056));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_A (.DIODE(net1078));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_A2 (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_B1_N (.DIODE(net1036));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_Y (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_A (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_B (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_Y (.DIODE(net666));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_A2 (.DIODE(net666));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_A3 (.DIODE(net1062));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_B1 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_Y (.DIODE(net675));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_B (.DIODE(net1043));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_A2 (.DIODE(net1028));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_A4 (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_A2 (.DIODE(net673));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_B1_N (.DIODE(net1052));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_B1_N (.DIODE(net1050));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_B1_N (.DIODE(net602));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_X (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_A1 (.DIODE(net1095));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_A2 (.DIODE(net1093));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_X (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_B1_N (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_X (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_A2 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_A3 (.DIODE(net1092));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_A4 (.DIODE(net1034));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_X (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_B1_N (.DIODE(net636));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_X (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_B (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_A1 (.DIODE(net586));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_A2 (.DIODE(net1092));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_B1_N (.DIODE(net1091));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_B1_N (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_A3 (.DIODE(net647));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_A4 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_B1 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_A (.DIODE(net680));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_A1 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_A2 (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_A3 (.DIODE(net692));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_A4 (.DIODE(net1112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_B1 (.DIODE(net1071));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_A1 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_A2 (.DIODE(net636));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_X (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_B1_N (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_A1 (.DIODE(net575));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_A2 (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_S1 (.DIODE(net1105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_A1 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_B1_N (.DIODE(net675));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_B (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_Y (.DIODE(net668));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_A1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_A2 (.DIODE(net586));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_X (.DIODE(net670));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_B1_N (.DIODE(net607));
 sky130_fd_sc_hd__diode_2 ANTENNA_c482_X (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_B1_N (.DIODE(net1053));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_A0 (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_A1 (.DIODE(net601));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_A2 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_S0 (.DIODE(net652));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_S1 (.DIODE(net1033));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_A1 (.DIODE(net583));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_A2 (.DIODE(net1037));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_B1_N (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_A (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_A1 (.DIODE(net663));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_A2 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_B1_N (.DIODE(net1083));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_X (.DIODE(net672));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_A (.DIODE(net607));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_A3 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_A4 (.DIODE(net672));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_B1 (.DIODE(net1083));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_X (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_A1 (.DIODE(net652));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_B1_N (.DIODE(net696));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_A (.DIODE(net541));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_A1 (.DIODE(net722));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_A2 (.DIODE(net663));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_S0 (.DIODE(net1055));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_A1 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_B1_N (.DIODE(net1148));
 sky130_fd_sc_hd__diode_2 ANTENNA_c494_B (.DIODE(net602));
 sky130_fd_sc_hd__diode_2 ANTENNA_c494_Y (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_A1 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_A2 (.DIODE(net1148));
 sky130_fd_sc_hd__diode_2 ANTENNA_c496_B1_N (.DIODE(net1114));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_A0 (.DIODE(net627));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_A2 (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_A3 (.DIODE(net652));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_S0 (.DIODE(net633));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_S1 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_A0 (.DIODE(net658));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_A3 (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_S0 (.DIODE(net627));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_B1_N (.DIODE(net1076));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_X (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_A (.DIODE(net541));
 sky130_fd_sc_hd__diode_2 ANTENNA_c502_B (.DIODE(net680));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_A (.DIODE(net1082));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_A2 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_S0 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_A0 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_A1 (.DIODE(net647));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_A2 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_S0 (.DIODE(net645));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_S1 (.DIODE(net688));
 sky130_fd_sc_hd__diode_2 ANTENNA_c528_B (.DIODE(net1044));
 sky130_fd_sc_hd__diode_2 ANTENNA_c528_Y (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_c530_A (.DIODE(net1057));
 sky130_fd_sc_hd__diode_2 ANTENNA_c531_A (.DIODE(net1101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c532_A (.DIODE(net573));
 sky130_fd_sc_hd__diode_2 ANTENNA_c533_A (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_c534_A (.DIODE(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA_c536_B (.DIODE(net1143));
 sky130_fd_sc_hd__diode_2 ANTENNA_c537_Y (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c538_B (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA_c539_Y (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c540_A (.DIODE(net1119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c541_A1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c541_B1 (.DIODE(net1101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c542_A (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c543_B (.DIODE(net674));
 sky130_fd_sc_hd__diode_2 ANTENNA_c544_A2 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c544_B1_N (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c544_X (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA_c545_B (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c546_Y (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA_c547_B (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_c547_Y (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_c548_A (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA_c548_Y (.DIODE(net677));
 sky130_fd_sc_hd__diode_2 ANTENNA_c549_A (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA_c549_B (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_c549_Y (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_A (.DIODE(net1098));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_A1 (.DIODE(net593));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_A2 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_A2 (.DIODE(net1074));
 sky130_fd_sc_hd__diode_2 ANTENNA_c554_A2 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c555_A (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_c556_B (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA_c557_A2 (.DIODE(net1069));
 sky130_fd_sc_hd__diode_2 ANTENNA_c558_A2 (.DIODE(net633));
 sky130_fd_sc_hd__diode_2 ANTENNA_c559_A (.DIODE(net597));
 sky130_fd_sc_hd__diode_2 ANTENNA_c560_A2 (.DIODE(net1044));
 sky130_fd_sc_hd__diode_2 ANTENNA_c561_B1_N (.DIODE(net1098));
 sky130_fd_sc_hd__diode_2 ANTENNA_c566_A1 (.DIODE(net519));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_Y (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_B1_N (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_A0 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_S0 (.DIODE(net1028));
 sky130_fd_sc_hd__diode_2 ANTENNA_c571_A2 (.DIODE(net597));
 sky130_fd_sc_hd__diode_2 ANTENNA_c571_X (.DIODE(net676));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_B1_N (.DIODE(net1143));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_B (.DIODE(net618));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_B1_N (.DIODE(net1049));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_X (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_B1 (.DIODE(net675));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_A (.DIODE(net1128));
 sky130_fd_sc_hd__diode_2 ANTENNA_c577_A2 (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_A2 (.DIODE(net674));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_B1_N (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_A2 (.DIODE(net1068));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_B1_N (.DIODE(net1103));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_A1 (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_A2 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_B1_N (.DIODE(net1054));
 sky130_fd_sc_hd__diode_2 ANTENNA_c582_B1_N (.DIODE(net1105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_A (.DIODE(net1128));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_X (.DIODE(net1153));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_A2 (.DIODE(net1105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_B1_N (.DIODE(net1076));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_A2 (.DIODE(net1055));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_A3 (.DIODE(net1121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_B1 (.DIODE(net1153));
 sky130_fd_sc_hd__diode_2 ANTENNA_c586_A2 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c586_B1_N (.DIODE(net1101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c587_A0 (.DIODE(net1074));
 sky130_fd_sc_hd__diode_2 ANTENNA_c587_A2 (.DIODE(net1153));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_A (.DIODE(net618));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_A0 (.DIODE(net1050));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_A1 (.DIODE(net1044));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_S1 (.DIODE(net677));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_X (.DIODE(net671));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_B (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_Y (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_A0 (.DIODE(net1116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_A2 (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_A3 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_S1 (.DIODE(net1046));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_A2 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_B1_N (.DIODE(net1153));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_A1 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_A2 (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_B1_N (.DIODE(net1153));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_A3 (.DIODE(net1072));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_B1 (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_B1_N (.DIODE(net643));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_A2 (.DIODE(net1028));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_B1_N (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_A2 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_B (.DIODE(net1049));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_Y (.DIODE(net1039));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_X (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_A1 (.DIODE(net643));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_A2 (.DIODE(net1117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_B1_N (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_A2 (.DIODE(net1039));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_A0 (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_A2 (.DIODE(net668));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_A3 (.DIODE(net1121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_S0 (.DIODE(net1039));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_S1 (.DIODE(net1095));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_A2 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_B1_N (.DIODE(net1039));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_A3 (.DIODE(net1039));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_B1 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c610_A2 (.DIODE(net1107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c611_A1 (.DIODE(net1054));
 sky130_fd_sc_hd__diode_2 ANTENNA_c611_A3 (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_A1 (.DIODE(net1062));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_A2 (.DIODE(net1039));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_A3 (.DIODE(net1056));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_S0 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c615_X (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_A1 (.DIODE(net1105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_A2 (.DIODE(net1078));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_A3 (.DIODE(net668));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_A4 (.DIODE(net1057));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_B1 (.DIODE(net1039));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_A0 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_A2 (.DIODE(net581));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_A3 (.DIODE(net1121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_S0 (.DIODE(net646));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_S1 (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_A2 (.DIODE(net1052));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_A3 (.DIODE(net1025));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_A4 (.DIODE(net670));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_B1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_A2 (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_A3 (.DIODE(net669));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_S0 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_S1 (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_A3 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_A4 (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_B1 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_A3 (.DIODE(net672));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_A4 (.DIODE(net670));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_B1 (.DIODE(net1059));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_A2 (.DIODE(net1065));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_A3 (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_B1 (.DIODE(net1132));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_A1 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_A2 (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_A3 (.DIODE(net1103));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_B1 (.DIODE(net1045));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_CLK_N (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_D (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_RESET_B (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_SCD (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_A2 (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_A3 (.DIODE(net1055));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_A0 (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_A2 (.DIODE(net646));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_S0 (.DIODE(net1025));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_A1 (.DIODE(net581));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_A2 (.DIODE(net1065));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_A3 (.DIODE(net1078));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_S1 (.DIODE(net1025));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_X (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_A1 (.DIODE(net584));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_B1_N (.DIODE(net674));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_A0 (.DIODE(net1055));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_A1 (.DIODE(net1039));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_A3 (.DIODE(net1105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_S0 (.DIODE(net1111));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_A2 (.DIODE(net1095));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_A3 (.DIODE(net1108));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_A4 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_B1 (.DIODE(net1033));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_A2 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_A4 (.DIODE(net1057));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_B1 (.DIODE(net1117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c633_A2 (.DIODE(net1127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c633_A4 (.DIODE(net672));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_CLK_N (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_D (.DIODE(net575));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_RESET_B (.DIODE(net1056));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_SCD (.DIODE(net1102));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_SET_B (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_A0 (.DIODE(net1108));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_A2 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_A3 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_X (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_CLK (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_RESET_B (.DIODE(net676));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_SCD (.DIODE(net1045));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_A2 (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_A3 (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_S0 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_S1 (.DIODE(net1151));
 sky130_fd_sc_hd__diode_2 ANTENNA_c660_A (.DIODE(net1122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c660_B (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c661_A (.DIODE(net570));
 sky130_fd_sc_hd__diode_2 ANTENNA_c662_A (.DIODE(net600));
 sky130_fd_sc_hd__diode_2 ANTENNA_c662_Y (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA_c663_B (.DIODE(net1063));
 sky130_fd_sc_hd__diode_2 ANTENNA_c664_A (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA_c665_A (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA_c666_B (.DIODE(net1058));
 sky130_fd_sc_hd__diode_2 ANTENNA_c667_A (.DIODE(net1156));
 sky130_fd_sc_hd__diode_2 ANTENNA_c667_B (.DIODE(net1058));
 sky130_fd_sc_hd__diode_2 ANTENNA_c668_A2 (.DIODE(net1049));
 sky130_fd_sc_hd__diode_2 ANTENNA_c669_A2 (.DIODE(net1119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c669_X (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_c670_B (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA_c671_B (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c674_A2 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA_c674_A3 (.DIODE(net1053));
 sky130_fd_sc_hd__diode_2 ANTENNA_c674_S1 (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA_c678_A2 (.DIODE(net1063));
 sky130_fd_sc_hd__diode_2 ANTENNA_c679_A2 (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA_c679_A3 (.DIODE(net1058));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_B (.DIODE(net1078));
 sky130_fd_sc_hd__diode_2 ANTENNA_c685_A1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c685_B1_N (.DIODE(net1074));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_A2 (.DIODE(net1122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_B1_N (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_A2 (.DIODE(net1053));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_A2 (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA_c691_B (.DIODE(net1059));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_A2 (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_B1_N (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA_c693_A (.DIODE(net1046));
 sky130_fd_sc_hd__diode_2 ANTENNA_c696_A2 (.DIODE(net1123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c698_A1 (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c698_A2 (.DIODE(net1063));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_A2 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_X (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA_c700_A1 (.DIODE(net1065));
 sky130_fd_sc_hd__diode_2 ANTENNA_c700_A2 (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA_c702_A1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c702_A2 (.DIODE(net751));
 sky130_fd_sc_hd__diode_2 ANTENNA_c703_A2 (.DIODE(net1151));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_B1_N (.DIODE(net1025));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_A2 (.DIODE(net1046));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_B1_N (.DIODE(net1069));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_A0 (.DIODE(net613));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_S1 (.DIODE(net666));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_B1_N (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_A2 (.DIODE(net1111));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_A3 (.DIODE(net1074));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_B1 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_A2 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_B1_N (.DIODE(net1112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_X (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_B1_N (.DIODE(net1111));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_B1_N (.DIODE(net1156));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_X (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_A2 (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_A3 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_S0 (.DIODE(net1072));
 sky130_fd_sc_hd__diode_2 ANTENNA_c720_A2 (.DIODE(net1059));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_A0 (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_A2 (.DIODE(net1072));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_A3 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_S0 (.DIODE(net1046));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_S1 (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_A3 (.DIODE(net1059));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_B1 (.DIODE(net1025));
 sky130_fd_sc_hd__diode_2 ANTENNA_c723_A2 (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA_c724_A2 (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c724_A3 (.DIODE(net1151));
 sky130_fd_sc_hd__diode_2 ANTENNA_c724_S1 (.DIODE(net1080));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_A0 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_A1 (.DIODE(net591));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_A3 (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_S1 (.DIODE(net1080));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A1 (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_B1_N (.DIODE(net1112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A2 (.DIODE(net591));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A3 (.DIODE(net1105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_B1 (.DIODE(net1122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_A1 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_B1 (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_CLK (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_SCD (.DIODE(net1069));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_A1 (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_B1 (.DIODE(net716));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_A1 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_A3 (.DIODE(net1108));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_S0 (.DIODE(net632));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_S1 (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_A1 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_A2 (.DIODE(net1091));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_A3 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_B1 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_A3 (.DIODE(net1025));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_B1 (.DIODE(net1074));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_A1 (.DIODE(net1069));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_A2 (.DIODE(net578));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_A2 (.DIODE(net1069));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_B1 (.DIODE(net1080));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_A3 (.DIODE(net751));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_A3 (.DIODE(net1144));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_S1 (.DIODE(net1059));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_A2 (.DIODE(net781));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_A3 (.DIODE(net1119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_S1 (.DIODE(net1080));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_A1 (.DIODE(net781));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_A2 (.DIODE(net1108));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_A3 (.DIODE(net1069));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_A0 (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_A2 (.DIODE(net578));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_S0 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c742_B1 (.DIODE(net1033));
 sky130_fd_sc_hd__diode_2 ANTENNA_c743_A1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c743_A2 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_c743_A3 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA_c743_A4 (.DIODE(net1096));
 sky130_fd_sc_hd__diode_2 ANTENNA_c744_A1 (.DIODE(net1107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c744_A3 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_c745_B1 (.DIODE(net1080));
 sky130_fd_sc_hd__diode_2 ANTENNA_c747_CLK (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c747_D (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_c747_Q (.DIODE(net490));
 sky130_fd_sc_hd__diode_2 ANTENNA_c747_SCD (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c747_SCE (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_A1 (.DIODE(net1111));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_A3 (.DIODE(net1156));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_S0 (.DIODE(net1072));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_S1 (.DIODE(net716));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_A1 (.DIODE(net1076));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_S0 (.DIODE(net490));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_S1 (.DIODE(net1103));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_A0 (.DIODE(net1068));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_A1 (.DIODE(net1033));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_A3 (.DIODE(net1123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_S1 (.DIODE(net716));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_A0 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_A1 (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_A2 (.DIODE(net1112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_A3 (.DIODE(net1074));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_S0 (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_A3 (.DIODE(net587));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_S0 (.DIODE(net1151));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_A0 (.DIODE(net632));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_A2 (.DIODE(net1105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_S1 (.DIODE(net1080));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A0 (.DIODE(net1102));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A1 (.DIODE(net1063));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_S0 (.DIODE(net1119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_S1 (.DIODE(net1074));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A0 (.DIODE(net1059));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A1 (.DIODE(net1103));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A2 (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_A0 (.DIODE(net1044));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_A1 (.DIODE(net641));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_A2 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_S0 (.DIODE(net1078));
 sky130_fd_sc_hd__diode_2 ANTENNA_c757_A0 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_c757_A2 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA_c757_S0 (.DIODE(net751));
 sky130_fd_sc_hd__diode_2 ANTENNA_c757_S1 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_A0 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_A3 (.DIODE(net1060));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_S0 (.DIODE(net1103));
 sky130_fd_sc_hd__diode_2 ANTENNA_c759_A1 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_c759_S0 (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_c760_A0 (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA_c760_A1 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA_c760_A2 (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA_c760_S0 (.DIODE(net1033));
 sky130_fd_sc_hd__diode_2 ANTENNA_c760_S1 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA_c761_A0 (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_c761_S0 (.DIODE(net1102));
 sky130_fd_sc_hd__diode_2 ANTENNA_c762_A0 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_c762_A1 (.DIODE(net1054));
 sky130_fd_sc_hd__diode_2 ANTENNA_c762_A3 (.DIODE(net641));
 sky130_fd_sc_hd__diode_2 ANTENNA_c762_S0 (.DIODE(net1080));
 sky130_fd_sc_hd__diode_2 ANTENNA_c763_A0 (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_c763_A3 (.DIODE(net490));
 sky130_fd_sc_hd__diode_2 ANTENNA_c763_S0 (.DIODE(net1065));
 sky130_fd_sc_hd__diode_2 ANTENNA_c764_A0 (.DIODE(net1053));
 sky130_fd_sc_hd__diode_2 ANTENNA_c764_A1 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA_c764_A3 (.DIODE(net590));
 sky130_fd_sc_hd__diode_2 ANTENNA_c765_A1 (.DIODE(net1103));
 sky130_fd_sc_hd__diode_2 ANTENNA_c765_A2 (.DIODE(net1072));
 sky130_fd_sc_hd__diode_2 ANTENNA_c765_S0 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA_c765_S1 (.DIODE(net1096));
 sky130_fd_sc_hd__diode_2 ANTENNA_c766_A1 (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA_c766_A2 (.DIODE(net590));
 sky130_fd_sc_hd__diode_2 ANTENNA_c766_A3 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_c766_S0 (.DIODE(net751));
 sky130_fd_sc_hd__diode_2 ANTENNA_c767_A3 (.DIODE(net1025));
 sky130_fd_sc_hd__diode_2 ANTENNA_c767_S1 (.DIODE(net1080));
 sky130_fd_sc_hd__diode_2 ANTENNA_c768_A1 (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA_c768_A3 (.DIODE(net587));
 sky130_fd_sc_hd__diode_2 ANTENNA_c769_A1 (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_A (.DIODE(clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_X (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_0__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_1__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_1__f_clk_X (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_2__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_2__f_clk_X (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_3__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_3__f_clk_X (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone22_A (.DIODE(net1128));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone22_X (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone5_X (.DIODE(net1033));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout175_A (.DIODE(net1025));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout175_X (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout176_X (.DIODE(net1025));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout178_A (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout178_X (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout179_A (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout179_X (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout180_X (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout181_A (.DIODE(net1144));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout181_X (.DIODE(net1034));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout182_X (.DIODE(net1038));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout203_A (.DIODE(net1089));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout203_X (.DIODE(net1085));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout204_X (.DIODE(net1089));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold58_A (.DIODE(net1081));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_X (.DIODE(net575));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_X (.DIODE(net1123));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_X (.DIODE(net577));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_X (.DIODE(net578));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_X (.DIODE(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_X (.DIODE(net1121));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_X (.DIODE(net581));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_X (.DIODE(net582));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_X (.DIODE(net583));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(net850));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_X (.DIODE(net584));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_X (.DIODE(net519));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_X (.DIODE(net1117));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_X (.DIODE(net586));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_A (.DIODE(net853));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_X (.DIODE(net587));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_A (.DIODE(net854));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_A (.DIODE(net855));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_X (.DIODE(net1116));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_A (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_X (.DIODE(net590));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_A (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_X (.DIODE(net591));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_A (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_X (.DIODE(net1114));
 sky130_fd_sc_hd__diode_2 ANTENNA_input28_A (.DIODE(net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_input28_X (.DIODE(net593));
 sky130_fd_sc_hd__diode_2 ANTENNA_input29_A (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_X (.DIODE(net1119));
 sky130_fd_sc_hd__diode_2 ANTENNA_input30_A (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_input30_X (.DIODE(net595));
 sky130_fd_sc_hd__diode_2 ANTENNA_input31_A (.DIODE(net862));
 sky130_fd_sc_hd__diode_2 ANTENNA_input31_X (.DIODE(net596));
 sky130_fd_sc_hd__diode_2 ANTENNA_input32_A (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_input32_X (.DIODE(net597));
 sky130_fd_sc_hd__diode_2 ANTENNA_input33_A (.DIODE(net864));
 sky130_fd_sc_hd__diode_2 ANTENNA_input33_X (.DIODE(net598));
 sky130_fd_sc_hd__diode_2 ANTENNA_input34_A (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_input34_X (.DIODE(net599));
 sky130_fd_sc_hd__diode_2 ANTENNA_input35_A (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_input35_X (.DIODE(net600));
 sky130_fd_sc_hd__diode_2 ANTENNA_input36_A (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_input36_X (.DIODE(net601));
 sky130_fd_sc_hd__diode_2 ANTENNA_input37_A (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_input37_X (.DIODE(net602));
 sky130_fd_sc_hd__diode_2 ANTENNA_input38_A (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_input38_X (.DIODE(net603));
 sky130_fd_sc_hd__diode_2 ANTENNA_input39_A (.DIODE(net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_input39_X (.DIODE(net604));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_X (.DIODE(net1113));
 sky130_fd_sc_hd__diode_2 ANTENNA_input40_A (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA_input41_A (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_input42_A (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_input42_X (.DIODE(net607));
 sky130_fd_sc_hd__diode_2 ANTENNA_input43_A (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_input44_A (.DIODE(net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_input44_X (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA_input45_A (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA_input46_A (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_input46_X (.DIODE(net1107));
 sky130_fd_sc_hd__diode_2 ANTENNA_input47_A (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_input47_X (.DIODE(net1105));
 sky130_fd_sc_hd__diode_2 ANTENNA_input48_A (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_input48_X (.DIODE(net613));
 sky130_fd_sc_hd__diode_2 ANTENNA_input49_A (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_X (.DIODE(net1108));
 sky130_fd_sc_hd__diode_2 ANTENNA_input50_A (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_input50_X (.DIODE(net615));
 sky130_fd_sc_hd__diode_2 ANTENNA_input51_A (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_input51_X (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA_input52_A (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_input52_X (.DIODE(net1104));
 sky130_fd_sc_hd__diode_2 ANTENNA_input53_A (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_input53_X (.DIODE(net618));
 sky130_fd_sc_hd__diode_2 ANTENNA_input54_A (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_input55_A (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_input55_X (.DIODE(net620));
 sky130_fd_sc_hd__diode_2 ANTENNA_input56_A (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_input56_X (.DIODE(net621));
 sky130_fd_sc_hd__diode_2 ANTENNA_input57_A (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_input57_X (.DIODE(net1102));
 sky130_fd_sc_hd__diode_2 ANTENNA_input58_A (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_input58_X (.DIODE(net623));
 sky130_fd_sc_hd__diode_2 ANTENNA_input59_A (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_X (.DIODE(net570));
 sky130_fd_sc_hd__diode_2 ANTENNA_input60_A (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_input61_A (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_input61_X (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA_input62_A (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_input62_X (.DIODE(net627));
 sky130_fd_sc_hd__diode_2 ANTENNA_input63_A (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_input64_A (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_input65_A (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_input66_A (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_input67_A (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_input67_X (.DIODE(net632));
 sky130_fd_sc_hd__diode_2 ANTENNA_input68_A (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_input68_X (.DIODE(net633));
 sky130_fd_sc_hd__diode_2 ANTENNA_input69_A (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_X (.DIODE(net1100));
 sky130_fd_sc_hd__diode_2 ANTENNA_input70_A (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_input71_A (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_input71_X (.DIODE(net636));
 sky130_fd_sc_hd__diode_2 ANTENNA_input72_A (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_input73_A (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_input74_A (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_input75_A (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_input76_A (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_input76_X (.DIODE(net641));
 sky130_fd_sc_hd__diode_2 ANTENNA_input77_A (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_input78_A (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_input78_X (.DIODE(net643));
 sky130_fd_sc_hd__diode_2 ANTENNA_input79_A (.DIODE(net910));
 sky130_fd_sc_hd__diode_2 ANTENNA_input79_X (.DIODE(net1098));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_X (.DIODE(net1099));
 sky130_fd_sc_hd__diode_2 ANTENNA_input80_A (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_input80_X (.DIODE(net645));
 sky130_fd_sc_hd__diode_2 ANTENNA_input81_A (.DIODE(net912));
 sky130_fd_sc_hd__diode_2 ANTENNA_input81_X (.DIODE(net646));
 sky130_fd_sc_hd__diode_2 ANTENNA_input82_A (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA_input82_X (.DIODE(net647));
 sky130_fd_sc_hd__diode_2 ANTENNA_input83_A (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA_input84_A (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_input85_A (.DIODE(net916));
 sky130_fd_sc_hd__diode_2 ANTENNA_input85_X (.DIODE(net650));
 sky130_fd_sc_hd__diode_2 ANTENNA_input86_A (.DIODE(net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_input87_A (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_input87_X (.DIODE(net652));
 sky130_fd_sc_hd__diode_2 ANTENNA_input88_A (.DIODE(net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_input89_A (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_input89_X (.DIODE(net654));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_X (.DIODE(net573));
 sky130_fd_sc_hd__diode_2 ANTENNA_input90_A (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_input90_X (.DIODE(net1095));
 sky130_fd_sc_hd__diode_2 ANTENNA_input91_A (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_input92_A (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_input93_A (.DIODE(net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_input93_X (.DIODE(net658));
 sky130_fd_sc_hd__diode_2 ANTENNA_input94_A (.DIODE(net925));
 sky130_fd_sc_hd__diode_2 ANTENNA_input94_X (.DIODE(net659));
 sky130_fd_sc_hd__diode_2 ANTENNA_input95_A (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_input95_X (.DIODE(net660));
 sky130_fd_sc_hd__diode_2 ANTENNA_input96_A (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_input97_A (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_input98_A (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_input98_X (.DIODE(net663));
 sky130_fd_sc_hd__diode_2 ANTENNA_input99_A (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_X (.DIODE(net1096));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap186_X (.DIODE(net751));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap187_A (.DIODE(net1058));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap190_X (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap192_X (.DIODE(net1055));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap194_A (.DIODE(net1156));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap194_X (.DIODE(net759));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap197_X (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap198_A (.DIODE(net1091));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap200_X (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap202_X (.DIODE(net1083));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge782_A4 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge784_A0 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge784_S1 (.DIODE(net1128));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge786_A1 (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge786_A3 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge786_S1 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge787_A1 (.DIODE(net595));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge787_B1 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge788_A4 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge788_X (.DIODE(net1128));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge789_A1 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge789_A2 (.DIODE(net613));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge789_S1 (.DIODE(net1128));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge790_A1 (.DIODE(net686));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge790_A2 (.DIODE(net641));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge790_S1 (.DIODE(net632));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge791_A3 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge791_S1 (.DIODE(net1116));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge792_A0 (.DIODE(net1036));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge792_A2 (.DIODE(net676));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge792_A3 (.DIODE(net591));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge792_S0 (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge792_S1 (.DIODE(net1117));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge793_CLK_N (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge793_D (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge793_RESET_B (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge793_SCD (.DIODE(net587));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge794_A1 (.DIODE(net660));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge794_A2 (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge794_S0 (.DIODE(net575));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge794_S1 (.DIODE(net663));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge795_A0 (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge795_A1 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge795_A2 (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge795_A3 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge795_S1 (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge796_A0 (.DIODE(net1062));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge796_A1 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge797_CLK (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge800_Y (.DIODE(net534));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge801_CLK_N (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge805_CLK (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge806_CLK (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge806_Q (.DIODE(net1128));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge807_CLK (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge807_Q (.DIODE(net1082));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge808_CLK (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge808_Q_N (.DIODE(net541));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge809_CLK (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge810_CLK (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge811_CLK (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge812_CLK (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge813_GATE_N (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge814_GATE_N (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge815_GATE (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge815_Q (.DIODE(net680));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge815_RESET_B (.DIODE(net534));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge817_GATE_N (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_output101_A (.DIODE(net666));
 sky130_fd_sc_hd__diode_2 ANTENNA_output102_A (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_output103_A (.DIODE(net668));
 sky130_fd_sc_hd__diode_2 ANTENNA_output104_A (.DIODE(net669));
 sky130_fd_sc_hd__diode_2 ANTENNA_output105_A (.DIODE(net670));
 sky130_fd_sc_hd__diode_2 ANTENNA_output106_A (.DIODE(net671));
 sky130_fd_sc_hd__diode_2 ANTENNA_output107_A (.DIODE(net672));
 sky130_fd_sc_hd__diode_2 ANTENNA_output108_A (.DIODE(net673));
 sky130_fd_sc_hd__diode_2 ANTENNA_output109_A (.DIODE(net674));
 sky130_fd_sc_hd__diode_2 ANTENNA_output110_A (.DIODE(net675));
 sky130_fd_sc_hd__diode_2 ANTENNA_output111_A (.DIODE(net676));
 sky130_fd_sc_hd__diode_2 ANTENNA_output112_A (.DIODE(net677));
 sky130_fd_sc_hd__diode_2 ANTENNA_output114_A (.DIODE(net679));
 sky130_fd_sc_hd__diode_2 ANTENNA_output115_A (.DIODE(net680));
 sky130_fd_sc_hd__diode_2 ANTENNA_output116_A (.DIODE(net1058));
 sky130_fd_sc_hd__diode_2 ANTENNA_output117_A (.DIODE(net1049));
 sky130_fd_sc_hd__diode_2 ANTENNA_output120_A (.DIODE(net1054));
 sky130_fd_sc_hd__diode_2 ANTENNA_output121_A (.DIODE(net686));
 sky130_fd_sc_hd__diode_2 ANTENNA_output123_A (.DIODE(net688));
 sky130_fd_sc_hd__diode_2 ANTENNA_output124_A (.DIODE(net689));
 sky130_fd_sc_hd__diode_2 ANTENNA_output127_A (.DIODE(net692));
 sky130_fd_sc_hd__diode_2 ANTENNA_output128_A (.DIODE(net693));
 sky130_fd_sc_hd__diode_2 ANTENNA_output131_A (.DIODE(net696));
 sky130_fd_sc_hd__diode_2 ANTENNA_output132_A (.DIODE(net1071));
 sky130_fd_sc_hd__diode_2 ANTENNA_output133_A (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_output137_A (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA_output140_A (.DIODE(net705));
 sky130_fd_sc_hd__diode_2 ANTENNA_output141_A (.DIODE(net706));
 sky130_fd_sc_hd__diode_2 ANTENNA_output142_A (.DIODE(net1025));
 sky130_fd_sc_hd__diode_2 ANTENNA_output146_A (.DIODE(net1048));
 sky130_fd_sc_hd__diode_2 ANTENNA_output148_A (.DIODE(net1088));
 sky130_fd_sc_hd__diode_2 ANTENNA_output149_A (.DIODE(net1082));
 sky130_fd_sc_hd__diode_2 ANTENNA_output151_A (.DIODE(net716));
 sky130_fd_sc_hd__diode_2 ANTENNA_output155_A (.DIODE(net720));
 sky130_fd_sc_hd__diode_2 ANTENNA_output157_A (.DIODE(net722));
 sky130_fd_sc_hd__diode_2 ANTENNA_output158_A (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_output159_A (.DIODE(net724));
 sky130_fd_sc_hd__diode_2 ANTENNA_output160_A (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA_output161_A (.DIODE(net1087));
 sky130_fd_sc_hd__diode_2 ANTENNA_output167_A (.DIODE(net1066));
 sky130_fd_sc_hd__diode_2 ANTENNA_output169_A (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_output170_A (.DIODE(net735));
 sky130_fd_sc_hd__diode_2 ANTENNA_output173_A (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer12_X (.DIODE(net781));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer33_A (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer34_A (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer53_X (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer56_A (.DIODE(net1034));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer6_X (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer7_A (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer8_A (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer8_X (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_s818_CLK (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s819_CLK (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s820_Q (.DIODE(net1080));
 sky130_fd_sc_hd__diode_2 ANTENNA_s821_Q (.DIODE(net716));
 sky130_fd_sc_hd__diode_2 ANTENNA_s822_CLK (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s823_CLK (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s824_CLK (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s825_CLK (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire191_X (.DIODE(net756));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Left_203 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Left_202 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Left_201 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Left_200 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Left_199 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Left_198 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Left_197 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Left_196 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Left_195 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Left_194 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Left_193 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Left_192 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Left_191 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Left_190 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Left_189 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Left_188 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Left_187 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Left_186 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Left_185 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Left_184 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Left_183 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_182 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_181 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_180 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_179 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_178 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_177 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_176 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_175 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_174 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_173 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_172 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_171 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_170 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_169 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_168 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_167 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_166 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_165 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_164 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_163 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_162 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_161 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Right_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Right_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Right_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Right_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Right_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Right_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Right_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Right_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Right_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Right_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Right_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Right_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Right_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Right_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Right_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Right_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Right_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Right_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Right_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Right_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Right_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_204 ();
 sky130_fd_sc_hd__a31o_1 c100 (.A1(net662),
    .A2(net608),
    .A3(net1090),
    .B1(net1094),
    .X(net688));
 sky130_fd_sc_hd__xnor2_2 c101 (.A(net629),
    .B(net648),
    .Y(net699));
 sky130_fd_sc_hd__a21bo_4 c102 (.A1(net604),
    .A2(net659),
    .B1_N(net1115),
    .X(net735));
 sky130_fd_sc_hd__xnor2_1 c103 (.A(net615),
    .B(net658),
    .Y(net0));
 sky130_fd_sc_hd__mux4_2 c104 (.A0(net657),
    .A1(net1083),
    .A2(net605),
    .A3(net615),
    .S0(net659),
    .S1(net1090),
    .X(net1));
 sky130_fd_sc_hd__a21bo_1 c105 (.A1(net1094),
    .A2(net1103),
    .B1_N(net1100),
    .X(net2));
 sky130_fd_sc_hd__xnor2_1 c106 (.A(net735),
    .B(net601),
    .Y(net3));
 sky130_fd_sc_hd__xnor2_2 c107 (.A(net664),
    .B(net735),
    .Y(net703));
 sky130_fd_sc_hd__xnor2_1 c108 (.A(net1),
    .B(net607),
    .Y(net728));
 sky130_fd_sc_hd__mux4_2 c109 (.A0(net631),
    .A1(net653),
    .A2(net2),
    .A3(net728),
    .S0(net663),
    .S1(net1094),
    .X(net722));
 sky130_fd_sc_hd__xnor2_1 c110 (.A(net1109),
    .B(net603),
    .Y(net704));
 sky130_fd_sc_hd__xnor2_1 c111 (.A(net657),
    .B(net623),
    .Y(net4));
 sky130_fd_sc_hd__xnor2_1 c112 (.A(net1114),
    .B(net699),
    .Y(net721));
 sky130_fd_sc_hd__xnor2_4 c113 (.A(net595),
    .B(net623),
    .Y(net5));
 sky130_fd_sc_hd__xnor2_1 c114 (.A(net587),
    .B(net722),
    .Y(net701));
 sky130_fd_sc_hd__xnor2_1 c115 (.A(net4),
    .B(net620),
    .Y(net6));
 sky130_fd_sc_hd__xnor2_2 c116 (.A(net571),
    .B(net703),
    .Y(net7));
 sky130_fd_sc_hd__xnor2_1 c117 (.A(net648),
    .B(net605),
    .Y(net736));
 sky130_fd_sc_hd__xnor2_4 c118 (.A(net662),
    .B(net5),
    .Y(net731));
 sky130_fd_sc_hd__xnor2_4 c119 (.A(net731),
    .B(net645),
    .Y(net8));
 sky130_fd_sc_hd__xnor2_1 c120 (.A(net8),
    .B(net648),
    .Y(net695));
 sky130_fd_sc_hd__xnor2_2 c121 (.A(net1),
    .B(net8),
    .Y(net9));
 sky130_fd_sc_hd__xnor2_2 c122 (.A(net620),
    .B(net8),
    .Y(net10));
 sky130_fd_sc_hd__xnor2_1 c123 (.A(net9),
    .B(net605),
    .Y(net710));
 sky130_fd_sc_hd__xnor2_1 c124 (.A(net9),
    .B(net10),
    .Y(net717));
 sky130_fd_sc_hd__xnor2_1 c125 (.A(net10),
    .B(net595),
    .Y(net11));
 sky130_fd_sc_hd__xnor2_1 c126 (.A(net6),
    .B(net8),
    .Y(net715));
 sky130_fd_sc_hd__xnor2_1 c127 (.A(net5),
    .B(net1094),
    .Y(net693));
 sky130_fd_sc_hd__a21bo_1 c128 (.A1(net2),
    .A2(net693),
    .B1_N(net717),
    .X(net737));
 sky130_fd_sc_hd__xnor2_1 c129 (.A(net7),
    .B(net737),
    .Y(net730));
 sky130_fd_sc_hd__xnor2_1 c130 (.A(net11),
    .B(net10),
    .Y(net12));
 sky130_fd_sc_hd__a21bo_1 c131 (.A1(net12),
    .A2(net603),
    .B1_N(net737),
    .X(net712));
 sky130_fd_sc_hd__xnor2_4 c132 (.A(net633),
    .B(net1096),
    .Y(net13));
 sky130_fd_sc_hd__xnor2_4 c133 (.A(net1110),
    .B(net1113),
    .Y(net738));
 sky130_fd_sc_hd__xnor2_4 c134 (.A(net765),
    .B(net1100),
    .Y(net14));
 sky130_fd_sc_hd__xnor2_4 c135 (.A(net1110),
    .B(net1108),
    .Y(net15));
 sky130_fd_sc_hd__xnor2_4 c136 (.A(net770),
    .B(net14),
    .Y(net16));
 sky130_fd_sc_hd__xnor2_2 c137 (.A(net771),
    .B(net1097),
    .Y(net17));
 sky130_fd_sc_hd__a21bo_1 c138 (.A1(net16),
    .A2(net1078),
    .B1_N(net1102),
    .X(net18));
 sky130_fd_sc_hd__xnor2_2 c139 (.A(net766),
    .B(net570),
    .Y(net19));
 sky130_fd_sc_hd__xnor2_4 c140 (.A(net1119),
    .B(net772),
    .Y(net729));
 sky130_fd_sc_hd__xnor2_4 c141 (.A(net570),
    .B(net762),
    .Y(net732));
 sky130_fd_sc_hd__a31o_1 c142 (.A1(net15),
    .A2(net1100),
    .A3(net766),
    .B1(net729),
    .X(net20));
 sky130_fd_sc_hd__xnor2_4 c143 (.A(net1096),
    .B(net759),
    .Y(net21));
 sky130_fd_sc_hd__a21bo_4 c144 (.A1(net577),
    .A2(net1097),
    .B1_N(net21),
    .X(net22));
 sky130_fd_sc_hd__xnor2_4 c145 (.A(net16),
    .B(net577),
    .Y(net23));
 sky130_fd_sc_hd__mux4_2 c146 (.A0(net1076),
    .A1(net1119),
    .A2(net729),
    .A3(net1099),
    .S0(net1093),
    .S1(net14),
    .X(net24));
 sky130_fd_sc_hd__xnor2_4 c147 (.A(net1064),
    .B(net729),
    .Y(net25));
 sky130_fd_sc_hd__xnor2_2 c148 (.A(net729),
    .B(net23),
    .Y(net26));
 sky130_fd_sc_hd__a21bo_2 c149 (.A1(net25),
    .A2(net24),
    .B1_N(net23),
    .X(net27));
 sky130_fd_sc_hd__a31o_2 c150 (.A1(net22),
    .A2(net25),
    .A3(net759),
    .B1(net23),
    .X(net685));
 sky130_fd_sc_hd__a21bo_2 c151 (.A1(net24),
    .A2(net1054),
    .B1_N(net23),
    .X(net28));
 sky130_fd_sc_hd__a21bo_2 c152 (.A1(net25),
    .A2(net1099),
    .B1_N(net729),
    .X(net29));
 sky130_fd_sc_hd__mux4_2 c153 (.A0(net1053),
    .A1(net24),
    .A2(net22),
    .A3(net27),
    .S0(net1057),
    .S1(net754),
    .X(net682));
 sky130_fd_sc_hd__xnor2_4 c154 (.A(net603),
    .B(net1115),
    .Y(net30));
 sky130_fd_sc_hd__xnor2_4 c155 (.A(net593),
    .B(net577),
    .Y(net733));
 sky130_fd_sc_hd__xnor2_4 c156 (.A(net577),
    .B(net1118),
    .Y(net31));
 sky130_fd_sc_hd__a31o_4 c157 (.A1(net582),
    .A2(net1100),
    .A3(net597),
    .B1(net1086),
    .X(net32));
 sky130_fd_sc_hd__xnor2_4 c158 (.A(net594),
    .B(net32),
    .Y(net724));
 sky130_fd_sc_hd__xnor2_2 c159 (.A(net13),
    .B(net1085),
    .Y(net33));
 sky130_fd_sc_hd__xnor2_2 c160 (.A(net1097),
    .B(net1086),
    .Y(net34));
 sky130_fd_sc_hd__xnor2_4 c161 (.A(net1107),
    .B(net1115),
    .Y(net35));
 sky130_fd_sc_hd__xnor2_4 c162 (.A(net35),
    .B(net761),
    .Y(net36));
 sky130_fd_sc_hd__xnor2_4 c163 (.A(net733),
    .B(net519),
    .Y(net37));
 sky130_fd_sc_hd__xnor2_1 c164 (.A(net584),
    .B(net583),
    .Y(net38));
 sky130_fd_sc_hd__mux4_2 c165 (.A0(net724),
    .A1(net37),
    .A2(net31),
    .A3(net754),
    .S0(net1085),
    .S1(net1108),
    .X(net39));
 sky130_fd_sc_hd__a21bo_1 c166 (.A1(net32),
    .A2(net604),
    .B1_N(net1086),
    .X(net40));
 sky130_fd_sc_hd__a31o_2 c167 (.A1(net38),
    .A2(net761),
    .A3(net1086),
    .B1(net1092),
    .X(net41));
 sky130_fd_sc_hd__xnor2_2 c168 (.A(net579),
    .B(net733),
    .Y(net713));
 sky130_fd_sc_hd__a21bo_1 c169 (.A1(net1092),
    .A2(net604),
    .B1_N(net41),
    .X(net42));
 sky130_fd_sc_hd__a21bo_4 c170 (.A1(net1069),
    .A2(net37),
    .B1_N(net39),
    .X(net43));
 sky130_fd_sc_hd__a21bo_1 c171 (.A1(net1092),
    .A2(net41),
    .B1_N(net1062),
    .X(net44));
 sky130_fd_sc_hd__a21bo_4 c172 (.A1(net31),
    .A2(net594),
    .B1_N(net43),
    .X(net45));
 sky130_fd_sc_hd__a31o_4 c173 (.A1(net1052),
    .A2(net1116),
    .A3(net593),
    .B1(net1061),
    .X(net46));
 sky130_fd_sc_hd__a21bo_4 c174 (.A1(net39),
    .A2(net1065),
    .B1_N(net1052),
    .X(net734));
 sky130_fd_sc_hd__a21bo_1 c175 (.A1(net734),
    .A2(net1052),
    .B1_N(net46),
    .X(net47));
 sky130_fd_sc_hd__xnor2_1 c176 (.A(net24),
    .B(net620),
    .Y(net48));
 sky130_fd_sc_hd__xnor2_4 c177 (.A(net633),
    .B(net734),
    .Y(net49));
 sky130_fd_sc_hd__a21bo_2 c178 (.A1(net620),
    .A2(net627),
    .B1_N(net1059),
    .X(net50));
 sky130_fd_sc_hd__xnor2_4 c179 (.A(net1110),
    .B(net628),
    .Y(net51));
 sky130_fd_sc_hd__a21bo_1 c180 (.A1(net625),
    .A2(net1067),
    .B1_N(net39),
    .X(net52));
 sky130_fd_sc_hd__xnor2_4 c181 (.A(net51),
    .B(net624),
    .Y(net673));
 sky130_fd_sc_hd__xnor2_2 c182 (.A(net614),
    .B(net673),
    .Y(net53));
 sky130_fd_sc_hd__xnor2_2 c183 (.A(net52),
    .B(net614),
    .Y(net54));
 sky130_fd_sc_hd__xnor2_2 c184 (.A(net49),
    .B(net22),
    .Y(net55));
 sky130_fd_sc_hd__a21bo_2 c185 (.A1(net1093),
    .A2(net625),
    .B1_N(net583),
    .X(net726));
 sky130_fd_sc_hd__a21bo_4 c186 (.A1(net54),
    .A2(net49),
    .B1_N(net53),
    .X(net56));
 sky130_fd_sc_hd__a21bo_2 c187 (.A1(net754),
    .A2(net1073),
    .B1_N(net1087),
    .X(net57));
 sky130_fd_sc_hd__xnor2_4 c188 (.A(net1073),
    .B(net1118),
    .Y(net58));
 sky130_fd_sc_hd__a31o_4 c189 (.A1(net55),
    .A2(net22),
    .A3(net1056),
    .B1(net1107),
    .X(net59));
 sky130_fd_sc_hd__a21bo_2 c190 (.A1(net619),
    .A2(net615),
    .B1_N(net1087),
    .X(net60));
 sky130_fd_sc_hd__xnor2_4 c191 (.A(net789),
    .B(net56),
    .Y(net61));
 sky130_fd_sc_hd__a21bo_1 c192 (.A1(net726),
    .A2(net50),
    .B1_N(net1086),
    .X(net62));
 sky130_fd_sc_hd__mux4_2 c193 (.A0(net38),
    .A1(net1037),
    .A2(net606),
    .A3(net1118),
    .S0(net59),
    .S1(net1086),
    .X(net63));
 sky130_fd_sc_hd__a21bo_1 c194 (.A1(net624),
    .A2(net53),
    .B1_N(net1056),
    .X(net64));
 sky130_fd_sc_hd__a21bo_2 c195 (.A1(net59),
    .A2(net1072),
    .B1_N(net38),
    .X(net65));
 sky130_fd_sc_hd__a31o_4 c196 (.A1(net63),
    .A2(net57),
    .A3(net65),
    .B1(net1106),
    .X(net66));
 sky130_fd_sc_hd__a31o_1 c197 (.A1(net66),
    .A2(net1088),
    .A3(net64),
    .B1(net59),
    .X(net67));
 sky130_fd_sc_hd__xnor2_4 c198 (.A(net639),
    .B(net1121),
    .Y(net709));
 sky130_fd_sc_hd__xnor2_1 c199 (.A(net630),
    .B(net50),
    .Y(net708));
 sky130_fd_sc_hd__xnor2_4 c200 (.A(net635),
    .B(net709),
    .Y(net68));
 sky130_fd_sc_hd__a21bo_1 c201 (.A1(net789),
    .A2(net1107),
    .B1_N(net709),
    .X(net711));
 sky130_fd_sc_hd__xnor2_4 c202 (.A(net1048),
    .B(net65),
    .Y(net69));
 sky130_fd_sc_hd__xnor2_1 c203 (.A(net1037),
    .B(net58),
    .Y(net70));
 sky130_fd_sc_hd__xnor2_2 c204 (.A(net638),
    .B(net637),
    .Y(net71));
 sky130_fd_sc_hd__xnor2_2 c205 (.A(net35),
    .B(net724),
    .Y(net72));
 sky130_fd_sc_hd__xnor2_2 c206 (.A(net69),
    .B(net709),
    .Y(net73));
 sky130_fd_sc_hd__xnor2_1 c207 (.A(net47),
    .B(net1073),
    .Y(net74));
 sky130_fd_sc_hd__a21bo_1 c208 (.A1(net70),
    .A2(net636),
    .B1_N(net1118),
    .X(net75));
 sky130_fd_sc_hd__xnor2_2 c209 (.A(net69),
    .B(net581),
    .Y(net76));
 sky130_fd_sc_hd__xnor2_1 c210 (.A(net73),
    .B(net75),
    .Y(net77));
 sky130_fd_sc_hd__xnor2_2 c211 (.A(net785),
    .B(net635),
    .Y(net706));
 sky130_fd_sc_hd__xnor2_1 c212 (.A(net77),
    .B(net649),
    .Y(net78));
 sky130_fd_sc_hd__mux4_2 c213 (.A0(net74),
    .A1(net78),
    .A2(net70),
    .A3(net726),
    .S0(net786),
    .S1(net73),
    .X(net79));
 sky130_fd_sc_hd__mux4_2 c214 (.A0(net628),
    .A1(net708),
    .A2(net711),
    .A3(net71),
    .S0(net650),
    .S1(net76),
    .X(net698));
 sky130_fd_sc_hd__xnor2_2 c215 (.A(net71),
    .B(net1011),
    .Y(net80));
 sky130_fd_sc_hd__xnor2_4 c216 (.A(net72),
    .B(net651),
    .Y(net81));
 sky130_fd_sc_hd__xnor2_4 c217 (.A(net81),
    .B(net1048),
    .Y(net82));
 sky130_fd_sc_hd__a21bo_1 c218 (.A1(net79),
    .A2(net82),
    .B1_N(net81),
    .X(net83));
 sky130_fd_sc_hd__a21bo_1 c219 (.A1(net82),
    .A2(net83),
    .B1_N(net81),
    .X(net84));
 sky130_fd_sc_hd__a31o_1 c220 (.A1(net39),
    .A2(net74),
    .A3(net659),
    .B1(net656),
    .X(net725));
 sky130_fd_sc_hd__a31o_2 c221 (.A1(net653),
    .A2(net68),
    .A3(net735),
    .B1(net800),
    .X(net85));
 sky130_fd_sc_hd__xnor2_4 c222 (.A(net68),
    .B(net595),
    .Y(net86));
 sky130_fd_sc_hd__a21bo_1 c223 (.A1(net634),
    .A2(net1083),
    .B1_N(net1118),
    .X(net87));
 sky130_fd_sc_hd__xnor2_4 c224 (.A(net758),
    .B(net1083),
    .Y(net88));
 sky130_fd_sc_hd__xnor2_1 c225 (.A(net1055),
    .B(net1094),
    .Y(net89));
 sky130_fd_sc_hd__xnor2_4 c226 (.A(net82),
    .B(net758),
    .Y(net669));
 sky130_fd_sc_hd__xnor2_1 c227 (.A(net87),
    .B(net1077),
    .Y(net90));
 sky130_fd_sc_hd__xnor2_4 c228 (.A(net608),
    .B(net86),
    .Y(net91));
 sky130_fd_sc_hd__a21bo_1 c229 (.A1(net90),
    .A2(net85),
    .B1_N(net711),
    .X(net702));
 sky130_fd_sc_hd__xnor2_2 c230 (.A(net758),
    .B(net88),
    .Y(net700));
 sky130_fd_sc_hd__xnor2_2 c231 (.A(net85),
    .B(net700),
    .Y(net92));
 sky130_fd_sc_hd__a21bo_2 c232 (.A1(net606),
    .A2(net47),
    .B1_N(net685),
    .X(net696));
 sky130_fd_sc_hd__xnor2_1 c233 (.A(net1121),
    .B(net669),
    .Y(net93));
 sky130_fd_sc_hd__xnor2_4 c234 (.A(net51),
    .B(net606),
    .Y(net94));
 sky130_fd_sc_hd__xnor2_1 c235 (.A(net659),
    .B(net576),
    .Y(net95));
 sky130_fd_sc_hd__a21bo_1 c236 (.A1(net801),
    .A2(net95),
    .B1_N(net608),
    .X(net723));
 sky130_fd_sc_hd__xnor2_2 c237 (.A(net91),
    .B(net88),
    .Y(net96));
 sky130_fd_sc_hd__xnor2_1 c238 (.A(net91),
    .B(net92),
    .Y(net727));
 sky130_fd_sc_hd__mux4_1 c239 (.A0(net29),
    .A1(net92),
    .A2(net727),
    .A3(net80),
    .S0(net1020),
    .S1(net89),
    .X(net97));
 sky130_fd_sc_hd__a21bo_1 c240 (.A1(net97),
    .A2(net80),
    .B1_N(net726),
    .X(net718));
 sky130_fd_sc_hd__a31o_1 c241 (.A1(net92),
    .A2(net86),
    .A3(net718),
    .B1(net94),
    .X(net739));
 sky130_fd_sc_hd__xnor2_4 c264 (.A(net573),
    .B(net570),
    .Y(net98));
 sky130_fd_sc_hd__xnor2_4 c265 (.A(net579),
    .B(net98),
    .Y(net99));
 sky130_fd_sc_hd__xnor2_4 c266 (.A(net572),
    .B(net1116),
    .Y(net719));
 sky130_fd_sc_hd__a21bo_1 c267 (.A1(net1096),
    .A2(net1102),
    .B1_N(net764),
    .X(net697));
 sky130_fd_sc_hd__xnor2_4 c268 (.A(net1099),
    .B(net1067),
    .Y(net100));
 sky130_fd_sc_hd__xnor2_2 c269 (.A(net764),
    .B(net784),
    .Y(net101));
 sky130_fd_sc_hd__xnor2_4 c270 (.A(net766),
    .B(net754),
    .Y(net102));
 sky130_fd_sc_hd__xnor2_2 c271 (.A(net719),
    .B(net764),
    .Y(net103));
 sky130_fd_sc_hd__xnor2_4 c272 (.A(net1095),
    .B(net1097),
    .Y(net104));
 sky130_fd_sc_hd__xnor2_4 c273 (.A(net750),
    .B(net764),
    .Y(net105));
 sky130_fd_sc_hd__xnor2_4 c274 (.A(net719),
    .B(net103),
    .Y(net106));
 sky130_fd_sc_hd__xnor2_2 c275 (.A(net1091),
    .B(net750),
    .Y(net107));
 sky130_fd_sc_hd__xnor2_2 c276 (.A(net1071),
    .B(net765),
    .Y(net108));
 sky130_fd_sc_hd__xnor2_4 c277 (.A(net100),
    .B(net1051),
    .Y(net109));
 sky130_fd_sc_hd__xnor2_2 c278 (.A(net763),
    .B(net105),
    .Y(net110));
 sky130_fd_sc_hd__xnor2_4 c279 (.A(net763),
    .B(net1051),
    .Y(net111));
 sky130_fd_sc_hd__a21bo_1 c280 (.A1(net101),
    .A2(net105),
    .B1_N(net111),
    .X(net112));
 sky130_fd_sc_hd__xnor2_4 c281 (.A(net1098),
    .B(net111),
    .Y(net113));
 sky130_fd_sc_hd__xnor2_4 c282 (.A(net760),
    .B(net99),
    .Y(net114));
 sky130_fd_sc_hd__xnor2_4 c283 (.A(net760),
    .B(net109),
    .Y(net115));
 sky130_fd_sc_hd__a21bo_1 c284 (.A1(net109),
    .A2(net763),
    .B1_N(net1047),
    .X(net116));
 sky130_fd_sc_hd__a41o_4 c285 (.A1(net1042),
    .A2(net1047),
    .A3(net1045),
    .A4(net1076),
    .B1(net1051),
    .X(net117));
 sky130_fd_sc_hd__xnor2_4 c286 (.A(net519),
    .B(net45),
    .Y(net118));
 sky130_fd_sc_hd__xnor2_4 c287 (.A(net1085),
    .B(net31),
    .Y(net689));
 sky130_fd_sc_hd__xnor2_2 c288 (.A(net689),
    .B(net118),
    .Y(net119));
 sky130_fd_sc_hd__xnor2_4 c289 (.A(net761),
    .B(net41),
    .Y(net120));
 sky130_fd_sc_hd__xnor2_4 c290 (.A(net601),
    .B(net102),
    .Y(net121));
 sky130_fd_sc_hd__xnor2_4 c291 (.A(net31),
    .B(net754),
    .Y(net122));
 sky130_fd_sc_hd__xnor2_2 c292 (.A(net825),
    .B(net599),
    .Y(net123));
 sky130_fd_sc_hd__a21bo_2 c293 (.A1(net118),
    .A2(net579),
    .B1_N(net1115),
    .X(net124));
 sky130_fd_sc_hd__xnor2_1 c294 (.A(net599),
    .B(net105),
    .Y(net125));
 sky130_fd_sc_hd__xnor2_2 c295 (.A(net121),
    .B(net33),
    .Y(net126));
 sky130_fd_sc_hd__a21bo_4 c296 (.A1(net122),
    .A2(net1050),
    .B1_N(net1035),
    .X(net127));
 sky130_fd_sc_hd__a21bo_1 c297 (.A1(net37),
    .A2(net33),
    .B1_N(net738),
    .X(net128));
 sky130_fd_sc_hd__xnor2_2 c298 (.A(net102),
    .B(net46),
    .Y(net129));
 sky130_fd_sc_hd__a21bo_2 c299 (.A1(net41),
    .A2(net586),
    .B1_N(net120),
    .X(net130));
 sky130_fd_sc_hd__a31o_1 c300 (.A1(net128),
    .A2(net584),
    .A3(net104),
    .B1(net1035),
    .X(net131));
 sky130_fd_sc_hd__xnor2_4 c301 (.A(net755),
    .B(net1067),
    .Y(net132));
 sky130_fd_sc_hd__a21bo_2 c302 (.A1(net753),
    .A2(net593),
    .B1_N(net582),
    .X(net133));
 sky130_fd_sc_hd__xnor2_2 c303 (.A(net127),
    .B(net120),
    .Y(net134));
 sky130_fd_sc_hd__a21bo_2 c304 (.A1(net124),
    .A2(net1050),
    .B1_N(net1041),
    .X(net135));
 sky130_fd_sc_hd__xnor2_4 c305 (.A(net135),
    .B(net133),
    .Y(net136));
 sky130_fd_sc_hd__mux4_2 c306 (.A0(net130),
    .A1(net136),
    .A2(net134),
    .A3(net132),
    .S0(net1041),
    .S1(net1035),
    .X(net137));
 sky130_fd_sc_hd__mux4_1 c307 (.A0(net27),
    .A1(net125),
    .A2(net753),
    .A3(net1035),
    .S0(net755),
    .S1(net1086),
    .X(net138));
 sky130_fd_sc_hd__xnor2_2 c308 (.A(net66),
    .B(net613),
    .Y(net139));
 sky130_fd_sc_hd__a21bo_1 c309 (.A1(net52),
    .A2(net1122),
    .B1_N(net1079),
    .X(net140));
 sky130_fd_sc_hd__xnor2_1 c310 (.A(net120),
    .B(net1103),
    .Y(net141));
 sky130_fd_sc_hd__xnor2_2 c311 (.A(net140),
    .B(net67),
    .Y(net142));
 sky130_fd_sc_hd__xnor2_2 c312 (.A(net627),
    .B(net623),
    .Y(net143));
 sky130_fd_sc_hd__xnor2_1 c313 (.A(net143),
    .B(net1043),
    .Y(net144));
 sky130_fd_sc_hd__xnor2_1 c314 (.A(net609),
    .B(net142),
    .Y(net145));
 sky130_fd_sc_hd__a21bo_1 c315 (.A1(net138),
    .A2(net609),
    .B1_N(net1030),
    .X(net146));
 sky130_fd_sc_hd__xnor2_1 c316 (.A(net824),
    .B(net143),
    .Y(net147));
 sky130_fd_sc_hd__xnor2_2 c317 (.A(net67),
    .B(net56),
    .Y(net148));
 sky130_fd_sc_hd__xnor2_1 c318 (.A(net55),
    .B(net1111),
    .Y(net149));
 sky130_fd_sc_hd__a21bo_1 c319 (.A1(net599),
    .A2(net148),
    .B1_N(net1050),
    .X(net150));
 sky130_fd_sc_hd__a21bo_1 c320 (.A1(net1029),
    .A2(net623),
    .B1_N(net1088),
    .X(net151));
 sky130_fd_sc_hd__a21bo_1 c321 (.A1(net142),
    .A2(net607),
    .B1_N(net673),
    .X(net152));
 sky130_fd_sc_hd__xnor2_1 c322 (.A(net1116),
    .B(net1019),
    .Y(net153));
 sky130_fd_sc_hd__xnor2_1 c323 (.A(net109),
    .B(net1124),
    .Y(net154));
 sky130_fd_sc_hd__a21bo_2 c324 (.A1(net1067),
    .A2(net1062),
    .B1_N(net1036),
    .X(net155));
 sky130_fd_sc_hd__xnor2_1 c325 (.A(net602),
    .B(net1041),
    .Y(net156));
 sky130_fd_sc_hd__xnor2_1 c326 (.A(net155),
    .B(net140),
    .Y(net707));
 sky130_fd_sc_hd__a21bo_1 c327 (.A1(net1019),
    .A2(net1016),
    .B1_N(net152),
    .X(net157));
 sky130_fd_sc_hd__mux4_1 c328 (.A0(net156),
    .A1(net149),
    .A2(net1115),
    .A3(net599),
    .S0(net1030),
    .S1(net621),
    .X(net158));
 sky130_fd_sc_hd__a21bo_1 c329 (.A1(net141),
    .A2(net158),
    .B1_N(net1019),
    .X(net159));
 sky130_fd_sc_hd__xnor2_2 c330 (.A(net698),
    .B(net54),
    .Y(net160));
 sky130_fd_sc_hd__xnor2_1 c331 (.A(net79),
    .B(net156),
    .Y(net161));
 sky130_fd_sc_hd__a41o_2 c332 (.A1(net83),
    .A2(net59),
    .A3(net1088),
    .A4(net1129),
    .B1(net1090),
    .X(net162));
 sky130_fd_sc_hd__a21bo_1 c333 (.A1(net53),
    .A2(net1037),
    .B1_N(net1036),
    .X(net163));
 sky130_fd_sc_hd__a41o_2 c334 (.A1(net583),
    .A2(net83),
    .A3(net1038),
    .A4(net1090),
    .B1(net1016),
    .X(net687));
 sky130_fd_sc_hd__a41o_1 c335 (.A1(net48),
    .A2(net1030),
    .A3(net123),
    .A4(net144),
    .B1(net825),
    .X(net164));
 sky130_fd_sc_hd__xnor2_2 c336 (.A(net610),
    .B(net73),
    .Y(net165));
 sky130_fd_sc_hd__a21bo_1 c337 (.A1(net156),
    .A2(net790),
    .B1_N(net161),
    .X(net166));
 sky130_fd_sc_hd__a41o_1 c338 (.A1(net107),
    .A2(net1036),
    .A3(net1049),
    .A4(net58),
    .B1(net1035),
    .X(net667));
 sky130_fd_sc_hd__a21bo_1 c339 (.A1(net149),
    .A2(net27),
    .B1_N(net687),
    .X(net167));
 sky130_fd_sc_hd__a21bo_1 c340 (.A1(net157),
    .A2(net1019),
    .B1_N(net1016),
    .X(net168));
 sky130_fd_sc_hd__xnor2_4 c341 (.A(net27),
    .B(net1024),
    .Y(net169));
 sky130_fd_sc_hd__a21bo_1 c342 (.A1(net637),
    .A2(net783),
    .B1_N(net1023),
    .X(net170));
 sky130_fd_sc_hd__a21bo_1 c343 (.A1(net1043),
    .A2(net165),
    .B1_N(net1023),
    .X(net171));
 sky130_fd_sc_hd__a21bo_1 c344 (.A1(net160),
    .A2(net169),
    .B1_N(net641),
    .X(net172));
 sky130_fd_sc_hd__a41o_2 c345 (.A1(net144),
    .A2(net146),
    .A3(net626),
    .A4(net1023),
    .B1(net1015),
    .X(net173));
 sky130_fd_sc_hd__a21bo_1 c346 (.A1(net75),
    .A2(net165),
    .B1_N(net171),
    .X(net174));
 sky130_fd_sc_hd__a21bo_1 c347 (.A1(net174),
    .A2(net823),
    .B1_N(net687),
    .X(net175));
 sky130_fd_sc_hd__a21bo_1 c348 (.A1(net161),
    .A2(net48),
    .B1_N(net1023),
    .X(net720));
 sky130_fd_sc_hd__buf_1 c349 (.A(net1082),
    .X(net176));
 sky130_fd_sc_hd__clkbuf_2 c350 (.A(net1082),
    .X(net177));
 sky130_fd_sc_hd__mux4_2 c351 (.A0(net171),
    .A1(net713),
    .A2(net177),
    .A3(net1024),
    .S0(net172),
    .S1(net1152),
    .X(net178));
 sky130_fd_sc_hd__a41o_1 c352 (.A1(net93),
    .A2(net640),
    .A3(net722),
    .A4(net642),
    .B1(net696),
    .X(net179));
 sky130_fd_sc_hd__a21bo_1 c353 (.A1(net134),
    .A2(net720),
    .B1_N(net1023),
    .X(net180));
 sky130_fd_sc_hd__a21bo_1 c354 (.A1(net168),
    .A2(net632),
    .B1_N(net776),
    .X(net181));
 sky130_fd_sc_hd__a21bo_1 c355 (.A1(net179),
    .A2(net1018),
    .B1_N(net1011),
    .X(net182));
 sky130_fd_sc_hd__xnor2_1 c356 (.A(net621),
    .B(net626),
    .Y(net183));
 sky130_fd_sc_hd__a21bo_1 c357 (.A1(net56),
    .A2(net789),
    .B1_N(net173),
    .X(net684));
 sky130_fd_sc_hd__mux4_1 c358 (.A0(net0),
    .A1(net29),
    .A2(net650),
    .A3(net1120),
    .S0(net574),
    .S1(net767),
    .X(net184));
 sky130_fd_sc_hd__a21bo_1 c359 (.A1(net654),
    .A2(net826),
    .B1_N(net184),
    .X(net185));
 sky130_fd_sc_hd__a21bo_1 c360 (.A1(net32),
    .A2(net621),
    .B1_N(net642),
    .X(net186));
 sky130_fd_sc_hd__a21bo_1 c361 (.A1(net117),
    .A2(net654),
    .B1_N(net183),
    .X(net187));
 sky130_fd_sc_hd__mux4_2 c362 (.A0(net88),
    .A1(net575),
    .A2(net85),
    .A3(net825),
    .S0(net702),
    .S1(net1089),
    .X(net188));
 sky130_fd_sc_hd__mux4_1 c363 (.A0(net146),
    .A1(net32),
    .A2(net1089),
    .A3(net650),
    .S0(net711),
    .S1(net80),
    .X(net705));
 sky130_fd_sc_hd__a41o_2 c364 (.A1(net168),
    .A2(net184),
    .A3(net1023),
    .A4(net1019),
    .B1(net706),
    .X(net189));
 sky130_fd_sc_hd__a21bo_1 c365 (.A1(net89),
    .A2(net183),
    .B1_N(net94),
    .X(net691));
 sky130_fd_sc_hd__xnor2_1 c366 (.A(net94),
    .B(net185),
    .Y(net190));
 sky130_fd_sc_hd__a21bo_1 c367 (.A1(net166),
    .A2(net1077),
    .B1_N(net1013),
    .X(net191));
 sky130_fd_sc_hd__a21bo_1 c368 (.A1(net190),
    .A2(net189),
    .B1_N(net1018),
    .X(net192));
 sky130_fd_sc_hd__a21bo_1 c369 (.A1(net80),
    .A2(net85),
    .B1_N(net189),
    .X(net193));
 sky130_fd_sc_hd__xnor2_1 c370 (.A(net165),
    .B(net91),
    .Y(net194));
 sky130_fd_sc_hd__buf_1 c371 (.A(net1082),
    .X(net195));
 sky130_fd_sc_hd__a21bo_1 c372 (.A1(net187),
    .A2(net189),
    .B1_N(net718),
    .X(net196));
 sky130_fd_sc_hd__a41o_1 c373 (.A1(net1118),
    .A2(net196),
    .A3(net61),
    .A4(net195),
    .B1(net189),
    .X(net197));
 sky130_fd_sc_hd__xnor2_4 c396 (.A(net114),
    .B(net580),
    .Y(net198));
 sky130_fd_sc_hd__xnor2_4 c397 (.A(net572),
    .B(net756),
    .Y(net199));
 sky130_fd_sc_hd__a21bo_4 c398 (.A1(net199),
    .A2(net764),
    .B1_N(net15),
    .X(net200));
 sky130_fd_sc_hd__xnor2_4 c399 (.A(net1098),
    .B(net1042),
    .Y(net201));
 sky130_fd_sc_hd__xnor2_4 c400 (.A(net111),
    .B(net1071),
    .Y(net202));
 sky130_fd_sc_hd__xnor2_1 c401 (.A(net1123),
    .B(net1063),
    .Y(net681));
 sky130_fd_sc_hd__xnor2_4 c402 (.A(net98),
    .B(net749),
    .Y(net203));
 sky130_fd_sc_hd__xnor2_4 c403 (.A(net201),
    .B(net198),
    .Y(net204));
 sky130_fd_sc_hd__xnor2_4 c404 (.A(net114),
    .B(net1068),
    .Y(net205));
 sky130_fd_sc_hd__xnor2_4 c405 (.A(net519),
    .B(net1123),
    .Y(net206));
 sky130_fd_sc_hd__a41o_2 c406 (.A1(net1045),
    .A2(net114),
    .A3(net749),
    .A4(net199),
    .B1(net752),
    .X(net207));
 sky130_fd_sc_hd__xnor2_4 c407 (.A(net202),
    .B(net199),
    .Y(net686));
 sky130_fd_sc_hd__xnor2_4 c408 (.A(net200),
    .B(net748),
    .Y(net208));
 sky130_fd_sc_hd__xnor2_4 c409 (.A(net206),
    .B(net752),
    .Y(net209));
 sky130_fd_sc_hd__xnor2_4 c410 (.A(net200),
    .B(net748),
    .Y(net210));
 sky130_fd_sc_hd__xnor2_4 c411 (.A(net203),
    .B(net205),
    .Y(net211));
 sky130_fd_sc_hd__xnor2_4 c412 (.A(net25),
    .B(net1095),
    .Y(net692));
 sky130_fd_sc_hd__xnor2_4 c413 (.A(net209),
    .B(net572),
    .Y(net212));
 sky130_fd_sc_hd__xnor2_4 c414 (.A(net212),
    .B(net749),
    .Y(net674));
 sky130_fd_sc_hd__xnor2_4 c415 (.A(net1127),
    .B(net212),
    .Y(net213));
 sky130_fd_sc_hd__xnor2_4 c416 (.A(net211),
    .B(net113),
    .Y(net214));
 sky130_fd_sc_hd__a41o_2 c417 (.A1(net1133),
    .A2(net101),
    .A3(net692),
    .A4(net200),
    .B1(net748),
    .X(net215));
 sky130_fd_sc_hd__xnor2_4 c418 (.A(net753),
    .B(net759),
    .Y(net216));
 sky130_fd_sc_hd__xnor2_2 c419 (.A(net1093),
    .B(net204),
    .Y(net217));
 sky130_fd_sc_hd__xnor2_2 c420 (.A(net18),
    .B(net1091),
    .Y(net218));
 sky130_fd_sc_hd__a31o_1 c421 (.A1(net217),
    .A2(net1068),
    .A3(net1071),
    .B1(net1038),
    .X(net219));
 sky130_fd_sc_hd__a41o_4 c422 (.A1(net111),
    .A2(net210),
    .A3(net1064),
    .A4(net212),
    .B1(net1074),
    .X(net220));
 sky130_fd_sc_hd__xnor2_4 c423 (.A(net30),
    .B(net127),
    .Y(net221));
 sky130_fd_sc_hd__xnor2_2 c424 (.A(net216),
    .B(net131),
    .Y(net222));
 sky130_fd_sc_hd__a21bo_2 c425 (.A1(net611),
    .A2(net207),
    .B1_N(net796),
    .X(net679));
 sky130_fd_sc_hd__a31o_2 c426 (.A1(net99),
    .A2(net46),
    .A3(net679),
    .B1(net1038),
    .X(net223));
 sky130_fd_sc_hd__a21bo_4 c427 (.A1(net218),
    .A2(net742),
    .B1_N(net121),
    .X(net224));
 sky130_fd_sc_hd__xnor2_4 c428 (.A(net46),
    .B(net220),
    .Y(net225));
 sky130_fd_sc_hd__xnor2_2 c429 (.A(net219),
    .B(net220),
    .Y(net226));
 sky130_fd_sc_hd__a21bo_1 c430 (.A1(net124),
    .A2(net222),
    .B1_N(net1068),
    .X(net227));
 sky130_fd_sc_hd__a21bo_1 c431 (.A1(net223),
    .A2(net1145),
    .B1_N(net226),
    .X(net228));
 sky130_fd_sc_hd__a21bo_2 c432 (.A1(net128),
    .A2(net228),
    .B1_N(net689),
    .X(net229));
 sky130_fd_sc_hd__mux4_2 c433 (.A0(net224),
    .A1(net1028),
    .A2(net742),
    .A3(net1115),
    .S0(net1098),
    .S1(net206),
    .X(net230));
 sky130_fd_sc_hd__xnor2_4 c434 (.A(net225),
    .B(net124),
    .Y(net231));
 sky130_fd_sc_hd__xnor2_4 c435 (.A(net796),
    .B(net231),
    .Y(net232));
 sky130_fd_sc_hd__xnor2_4 c436 (.A(net232),
    .B(net132),
    .Y(net233));
 sky130_fd_sc_hd__xnor2_2 c437 (.A(net230),
    .B(net1027),
    .Y(net234));
 sky130_fd_sc_hd__xnor2_1 c438 (.A(net229),
    .B(net792),
    .Y(net235));
 sky130_fd_sc_hd__xnor2_4 c439 (.A(net1028),
    .B(net679),
    .Y(net236));
 sky130_fd_sc_hd__xnor2_1 c440 (.A(net1112),
    .B(net233),
    .Y(net237));
 sky130_fd_sc_hd__a21bo_1 c441 (.A1(net1047),
    .A2(net234),
    .B1_N(net155),
    .X(net238));
 sky130_fd_sc_hd__a21bo_1 c442 (.A1(net235),
    .A2(net125),
    .B1_N(net57),
    .X(net239));
 sky130_fd_sc_hd__xnor2_4 c443 (.A(net220),
    .B(net58),
    .Y(net240));
 sky130_fd_sc_hd__xnor2_1 c444 (.A(net1079),
    .B(net155),
    .Y(net241));
 sky130_fd_sc_hd__a21bo_1 c445 (.A1(net159),
    .A2(net1042),
    .B1_N(net1036),
    .X(net242));
 sky130_fd_sc_hd__a21bo_1 c446 (.A1(net133),
    .A2(net100),
    .B1_N(net16),
    .X(net243));
 sky130_fd_sc_hd__xnor2_2 c447 (.A(net148),
    .B(net222),
    .Y(net244));
 sky130_fd_sc_hd__xnor2_4 c448 (.A(net616),
    .B(net106),
    .Y(net666));
 sky130_fd_sc_hd__a31o_1 c449 (.A1(net238),
    .A2(net666),
    .A3(net1062),
    .B1(net1016),
    .X(net245));
 sky130_fd_sc_hd__xnor2_4 c450 (.A(net240),
    .B(net1125),
    .Y(net675));
 sky130_fd_sc_hd__xnor2_2 c451 (.A(net218),
    .B(net1043),
    .Y(net246));
 sky130_fd_sc_hd__a41o_1 c452 (.A1(net152),
    .A2(net226),
    .A3(net155),
    .A4(net1160),
    .B1(net238),
    .X(net247));
 sky130_fd_sc_hd__a21bo_1 c453 (.A1(net245),
    .A2(net673),
    .B1_N(net45),
    .X(net248));
 sky130_fd_sc_hd__a21bo_1 c454 (.A1(net247),
    .A2(net233),
    .B1_N(net220),
    .X(net249));
 sky130_fd_sc_hd__a21bo_1 c455 (.A1(net153),
    .A2(net247),
    .B1_N(net1050),
    .X(net250));
 sky130_fd_sc_hd__xnor2_1 c456 (.A(net813),
    .B(net59),
    .Y(net251));
 sky130_fd_sc_hd__a21bo_1 c457 (.A1(net131),
    .A2(net251),
    .B1_N(net602),
    .X(net252));
 sky130_fd_sc_hd__xnor2_1 c458 (.A(net243),
    .B(net245),
    .Y(net253));
 sky130_fd_sc_hd__a21bo_1 c459 (.A1(net1095),
    .A2(net15),
    .B1_N(net246),
    .X(net254));
 sky130_fd_sc_hd__a21bo_1 c460 (.A1(net249),
    .A2(net250),
    .B1_N(net254),
    .X(net255));
 sky130_fd_sc_hd__a41o_2 c461 (.A1(net253),
    .A2(net1008),
    .A3(net30),
    .A4(net1035),
    .B1(net795),
    .X(net256));
 sky130_fd_sc_hd__a21bo_1 c462 (.A1(net78),
    .A2(net610),
    .B1_N(net636),
    .X(net257));
 sky130_fd_sc_hd__xnor2_1 c463 (.A(net251),
    .B(net1160),
    .Y(net258));
 sky130_fd_sc_hd__a21bo_1 c464 (.A1(net586),
    .A2(net30),
    .B1_N(net104),
    .X(net259));
 sky130_fd_sc_hd__a21bo_1 c465 (.A1(net16),
    .A2(net240),
    .B1_N(net162),
    .X(net260));
 sky130_fd_sc_hd__clkbuf_1 c466 (.A(net552),
    .X(net261));
 sky130_fd_sc_hd__a41o_1 c467 (.A1(net176),
    .A2(net100),
    .A3(net647),
    .A4(net232),
    .B1(net1015),
    .X(net262));
 sky130_fd_sc_hd__buf_1 c468 (.A(net680),
    .X(net263));
 sky130_fd_sc_hd__a41o_1 c469 (.A1(net64),
    .A2(net129),
    .A3(net692),
    .A4(net1112),
    .B1(net697),
    .X(net264));
 sky130_fd_sc_hd__a21bo_1 c470 (.A1(net209),
    .A2(net168),
    .B1_N(net794),
    .X(net265));
 sky130_fd_sc_hd__a21bo_2 c471 (.A1(net265),
    .A2(net636),
    .B1_N(net742),
    .X(net266));
 sky130_fd_sc_hd__a21bo_1 c472 (.A1(net259),
    .A2(net263),
    .B1_N(net1030),
    .X(net267));
 sky130_fd_sc_hd__mux4_1 c473 (.A0(net248),
    .A1(net575),
    .A2(net1160),
    .A3(net233),
    .S0(net239),
    .S1(net1106),
    .X(net268));
 sky130_fd_sc_hd__dlymetal6s2s_1 c474 (.A(net552),
    .X(net269));
 sky130_fd_sc_hd__a21bo_1 c475 (.A1(net205),
    .A2(net262),
    .B1_N(net264),
    .X(net270));
 sky130_fd_sc_hd__a21bo_1 c476 (.A1(net58),
    .A2(net262),
    .B1_N(net675),
    .X(net271));
 sky130_fd_sc_hd__clkbuf_1 c477 (.A(net552),
    .X(net272));
 sky130_fd_sc_hd__a21bo_1 c478 (.A1(net267),
    .A2(net272),
    .B1_N(net259),
    .X(net273));
 sky130_fd_sc_hd__xnor2_4 c479 (.A(net177),
    .B(net229),
    .Y(net668));
 sky130_fd_sc_hd__a21bo_2 c480 (.A1(net162),
    .A2(net586),
    .B1_N(net269),
    .X(net670));
 sky130_fd_sc_hd__a21bo_1 c481 (.A1(net100),
    .A2(net273),
    .B1_N(net607),
    .X(net274));
 sky130_fd_sc_hd__a21bo_1 c482 (.A1(net274),
    .A2(net270),
    .B1_N(net269),
    .X(net275));
 sky130_fd_sc_hd__a21bo_1 c483 (.A1(net246),
    .A2(net261),
    .B1_N(net1053),
    .X(net276));
 sky130_fd_sc_hd__mux4_2 c484 (.A0(net626),
    .A1(net601),
    .A2(net1015),
    .A3(net178),
    .S0(net652),
    .S1(net1033),
    .X(net694));
 sky130_fd_sc_hd__a21bo_1 c485 (.A1(net583),
    .A2(net1037),
    .B1_N(net1016),
    .X(net277));
 sky130_fd_sc_hd__xnor2_1 c486 (.A(net244),
    .B(net189),
    .Y(net278));
 sky130_fd_sc_hd__a21bo_2 c487 (.A1(net663),
    .A2(net200),
    .B1_N(net767),
    .X(net672));
 sky130_fd_sc_hd__xnor2_1 c488 (.A(net607),
    .B(net3),
    .Y(net279));
 sky130_fd_sc_hd__a41o_1 c489 (.A1(net181),
    .A2(net277),
    .A3(net96),
    .A4(net672),
    .B1(net767),
    .X(net280));
 sky130_fd_sc_hd__a21bo_1 c490 (.A1(net652),
    .A2(net95),
    .B1_N(net696),
    .X(net281));
 sky130_fd_sc_hd__clkbuf_1 c491 (.A(net541),
    .X(net282));
 sky130_fd_sc_hd__mux4_1 c492 (.A0(net178),
    .A1(net722),
    .A2(net663),
    .A3(net123),
    .S0(net1055),
    .S1(net189),
    .X(net283));
 sky130_fd_sc_hd__a21bo_1 c493 (.A1(net96),
    .A2(net661),
    .B1_N(net1148),
    .X(net678));
 sky130_fd_sc_hd__xnor2_2 c494 (.A(net182),
    .B(net602),
    .Y(net284));
 sky130_fd_sc_hd__a21bo_1 c495 (.A1(net228),
    .A2(net1147),
    .B1_N(net189),
    .X(net285));
 sky130_fd_sc_hd__a21bo_1 c496 (.A1(net123),
    .A2(net276),
    .B1_N(net1115),
    .X(net286));
 sky130_fd_sc_hd__mux4_1 c497 (.A0(net627),
    .A1(net191),
    .A2(net1011),
    .A3(net652),
    .S0(net633),
    .S1(net1015),
    .X(net287));
 sky130_fd_sc_hd__mux4_1 c498 (.A0(net658),
    .A1(net286),
    .A2(net189),
    .A3(net1011),
    .S0(net627),
    .S1(net694),
    .X(net288));
 sky130_fd_sc_hd__xnor2_1 c499 (.A(net95),
    .B(net92),
    .Y(net289));
 sky130_fd_sc_hd__a21bo_1 c500 (.A1(net186),
    .A2(net194),
    .B1_N(net1077),
    .X(net290));
 sky130_fd_sc_hd__clkbuf_1 c501 (.A(net541),
    .X(net291));
 sky130_fd_sc_hd__xnor2_1 c502 (.A(net3),
    .B(net680),
    .Y(net292));
 sky130_fd_sc_hd__clkbuf_1 c503 (.A(net1082),
    .X(net293));
 sky130_fd_sc_hd__mux4_1 c504 (.A0(net292),
    .A1(net293),
    .A2(net173),
    .A3(net163),
    .S0(net1024),
    .S1(net285),
    .X(net294));
 sky130_fd_sc_hd__mux4_1 c505 (.A0(net254),
    .A1(net647),
    .A2(net244),
    .A3(net283),
    .S0(net645),
    .S1(net688),
    .X(net295));
 sky130_fd_sc_hd__xnor2_4 c528 (.A(net213),
    .B(net1045),
    .Y(net296));
 sky130_fd_sc_hd__xnor2_4 c529 (.A(net203),
    .B(net211),
    .Y(net297));
 sky130_fd_sc_hd__xnor2_4 c530 (.A(net1057),
    .B(net297),
    .Y(net298));
 sky130_fd_sc_hd__xnor2_4 c531 (.A(net1101),
    .B(net215),
    .Y(net299));
 sky130_fd_sc_hd__xnor2_4 c532 (.A(net1097),
    .B(net21),
    .Y(net300));
 sky130_fd_sc_hd__xnor2_4 c533 (.A(net296),
    .B(net300),
    .Y(net301));
 sky130_fd_sc_hd__xnor2_1 c534 (.A(net579),
    .B(net298),
    .Y(net302));
 sky130_fd_sc_hd__xnor2_1 c535 (.A(net298),
    .B(net300),
    .Y(net303));
 sky130_fd_sc_hd__xnor2_4 c536 (.A(net798),
    .B(net600),
    .Y(net304));
 sky130_fd_sc_hd__xnor2_4 c537 (.A(net301),
    .B(net208),
    .Y(net305));
 sky130_fd_sc_hd__xnor2_2 c538 (.A(net199),
    .B(net756),
    .Y(net306));
 sky130_fd_sc_hd__xnor2_1 c539 (.A(net302),
    .B(net213),
    .Y(net307));
 sky130_fd_sc_hd__xnor2_2 c540 (.A(net1120),
    .B(net306),
    .Y(net308));
 sky130_fd_sc_hd__a41o_2 c541 (.A1(net117),
    .A2(net298),
    .A3(net308),
    .A4(net302),
    .B1(net1102),
    .X(net309));
 sky130_fd_sc_hd__xnor2_4 c542 (.A(net1012),
    .B(net299),
    .Y(net310));
 sky130_fd_sc_hd__xnor2_2 c543 (.A(net308),
    .B(net674),
    .Y(net311));
 sky130_fd_sc_hd__a21bo_2 c544 (.A1(net308),
    .A2(net1017),
    .B1_N(net1012),
    .X(net312));
 sky130_fd_sc_hd__xnor2_4 c545 (.A(net297),
    .B(net305),
    .Y(net313));
 sky130_fd_sc_hd__xnor2_4 c546 (.A(net304),
    .B(net313),
    .Y(net314));
 sky130_fd_sc_hd__xnor2_4 c547 (.A(net299),
    .B(net1032),
    .Y(net315));
 sky130_fd_sc_hd__xnor2_2 c548 (.A(net312),
    .B(net311),
    .Y(net677));
 sky130_fd_sc_hd__xnor2_4 c549 (.A(net314),
    .B(net315),
    .Y(net316));
 sky130_fd_sc_hd__xnor2_4 c550 (.A(net644),
    .B(net236),
    .Y(net317));
 sky130_fd_sc_hd__a21bo_1 c551 (.A1(net593),
    .A2(net130),
    .B1_N(net198),
    .X(net318));
 sky130_fd_sc_hd__xnor2_1 c552 (.A(net231),
    .B(net207),
    .Y(net319));
 sky130_fd_sc_hd__a21bo_1 c553 (.A1(net208),
    .A2(net1075),
    .B1_N(net317),
    .X(net320));
 sky130_fd_sc_hd__a41o_1 c554 (.A1(net212),
    .A2(net122),
    .A3(net236),
    .A4(net778),
    .B1(net317),
    .X(net321));
 sky130_fd_sc_hd__xnor2_1 c555 (.A(net130),
    .B(net321),
    .Y(net322));
 sky130_fd_sc_hd__xnor2_1 c556 (.A(net309),
    .B(net762),
    .Y(net323));
 sky130_fd_sc_hd__a21bo_1 c557 (.A1(net101),
    .A2(net1070),
    .B1_N(net208),
    .X(net324));
 sky130_fd_sc_hd__a21bo_1 c558 (.A1(net317),
    .A2(net633),
    .B1_N(net748),
    .X(net325));
 sky130_fd_sc_hd__xnor2_1 c559 (.A(net597),
    .B(net318),
    .Y(net326));
 sky130_fd_sc_hd__a21bo_1 c560 (.A1(net326),
    .A2(net1045),
    .B1_N(net799),
    .X(net327));
 sky130_fd_sc_hd__a21bo_1 c561 (.A1(net323),
    .A2(net322),
    .B1_N(net1098),
    .X(net328));
 sky130_fd_sc_hd__xnor2_1 c562 (.A(net236),
    .B(net300),
    .Y(net329));
 sky130_fd_sc_hd__xnor2_1 c563 (.A(net327),
    .B(net298),
    .Y(net330));
 sky130_fd_sc_hd__xnor2_1 c564 (.A(net321),
    .B(net330),
    .Y(net331));
 sky130_fd_sc_hd__a21bo_1 c565 (.A1(net326),
    .A2(net328),
    .B1_N(net779),
    .X(net332));
 sky130_fd_sc_hd__a21bo_1 c566 (.A1(net519),
    .A2(net327),
    .B1_N(net323),
    .X(net333));
 sky130_fd_sc_hd__xnor2_2 c567 (.A(net333),
    .B(net332),
    .Y(net334));
 sky130_fd_sc_hd__a21bo_2 c568 (.A1(net319),
    .A2(net13),
    .B1_N(net796),
    .X(net335));
 sky130_fd_sc_hd__a21bo_1 c569 (.A1(net328),
    .A2(net217),
    .B1_N(net1027),
    .X(net336));
 sky130_fd_sc_hd__mux4_1 c570 (.A0(net334),
    .A1(net332),
    .A2(net317),
    .A3(net329),
    .S0(net1028),
    .S1(net335),
    .X(net337));
 sky130_fd_sc_hd__a21bo_2 c571 (.A1(net336),
    .A2(net597),
    .B1_N(net335),
    .X(net676));
 sky130_fd_sc_hd__a21bo_1 c572 (.A1(net150),
    .A2(net336),
    .B1_N(net1110),
    .X(net338));
 sky130_fd_sc_hd__xnor2_1 c573 (.A(net310),
    .B(net618),
    .Y(net339));
 sky130_fd_sc_hd__a21bo_2 c574 (.A1(net215),
    .A2(net335),
    .B1_N(net1049),
    .X(net340));
 sky130_fd_sc_hd__a31o_1 c575 (.A1(net298),
    .A2(net135),
    .A3(net150),
    .B1(net675),
    .X(net341));
 sky130_fd_sc_hd__clkbuf_1 c576 (.A(net1141),
    .X(net342));
 sky130_fd_sc_hd__a21bo_1 c577 (.A1(net198),
    .A2(net340),
    .B1_N(net155),
    .X(net343));
 sky130_fd_sc_hd__a21bo_1 c578 (.A1(net323),
    .A2(net674),
    .B1_N(net1009),
    .X(net344));
 sky130_fd_sc_hd__clkbuf_1 c579 (.A(net543),
    .X(net345));
 sky130_fd_sc_hd__a21bo_1 c580 (.A1(net318),
    .A2(net108),
    .B1_N(net1104),
    .X(net346));
 sky130_fd_sc_hd__a21bo_1 c581 (.A1(net1041),
    .A2(net117),
    .B1_N(net1054),
    .X(net347));
 sky130_fd_sc_hd__a21bo_1 c582 (.A1(net346),
    .A2(net154),
    .B1_N(net1106),
    .X(net348));
 sky130_fd_sc_hd__buf_6 c583 (.A(net1007),
    .X(net349));
 sky130_fd_sc_hd__a21bo_1 c584 (.A1(net343),
    .A2(net1106),
    .B1_N(net1077),
    .X(net350));
 sky130_fd_sc_hd__a31o_4 c585 (.A1(net748),
    .A2(net1055),
    .A3(net580),
    .B1(net1006),
    .X(net351));
 sky130_fd_sc_hd__a21bo_1 c586 (.A1(net330),
    .A2(net1008),
    .B1_N(net1101),
    .X(net352));
 sky130_fd_sc_hd__mux4_2 c587 (.A0(net1075),
    .A1(net219),
    .A2(net1006),
    .A3(net301),
    .S0(net351),
    .S1(net320),
    .X(net353));
 sky130_fd_sc_hd__xnor2_1 c588 (.A(net618),
    .B(net319),
    .Y(net354));
 sky130_fd_sc_hd__mux4_2 c589 (.A0(net126),
    .A1(net1045),
    .A2(net346),
    .A3(net353),
    .S0(net325),
    .S1(net677),
    .X(net671));
 sky130_fd_sc_hd__xnor2_1 c590 (.A(net320),
    .B(net609),
    .Y(net355));
 sky130_fd_sc_hd__mux4_1 c591 (.A0(net1116),
    .A1(net155),
    .A2(net340),
    .A3(net121),
    .S0(net347),
    .S1(net1047),
    .X(net356));
 sky130_fd_sc_hd__a21bo_1 c592 (.A1(net348),
    .A2(net62),
    .B1_N(net1006),
    .X(net357));
 sky130_fd_sc_hd__a21bo_1 c593 (.A1(net62),
    .A2(net1010),
    .B1_N(net1006),
    .X(net358));
 sky130_fd_sc_hd__a31o_1 c594 (.A1(net264),
    .A2(net259),
    .A3(net1072),
    .B1(net791),
    .X(net359));
 sky130_fd_sc_hd__a21bo_1 c595 (.A1(net311),
    .A2(net304),
    .B1_N(net643),
    .X(net690));
 sky130_fd_sc_hd__clkbuf_1 c596 (.A(net547),
    .X(net360));
 sky130_fd_sc_hd__a21bo_1 c597 (.A1(net158),
    .A2(net226),
    .B1_N(net257),
    .X(net361));
 sky130_fd_sc_hd__a21bo_1 c598 (.A1(net241),
    .A2(net232),
    .B1_N(net169),
    .X(net362));
 sky130_fd_sc_hd__xnor2_1 c599 (.A(net313),
    .B(net797),
    .Y(net363));
 sky130_fd_sc_hd__xnor2_2 c600 (.A(net306),
    .B(net1131),
    .Y(net364));
 sky130_fd_sc_hd__a21bo_1 c601 (.A1(net235),
    .A2(net137),
    .B1_N(net268),
    .X(net365));
 sky130_fd_sc_hd__clkbuf_1 c602 (.A(net547),
    .X(net366));
 sky130_fd_sc_hd__a21bo_1 c603 (.A1(net643),
    .A2(net1118),
    .B1_N(net1009),
    .X(net367));
 sky130_fd_sc_hd__a21bo_1 c604 (.A1(net242),
    .A2(net1039),
    .B1_N(net137),
    .X(net368));
 sky130_fd_sc_hd__mux4_1 c605 (.A0(net365),
    .A1(net361),
    .A2(net668),
    .A3(net580),
    .S0(net1040),
    .S1(net1095),
    .X(net369));
 sky130_fd_sc_hd__clkbuf_1 c606 (.A(net547),
    .X(net370));
 sky130_fd_sc_hd__a21bo_1 c607 (.A1(net233),
    .A2(net1134),
    .B1_N(net169),
    .X(net371));
 sky130_fd_sc_hd__a21bo_1 c608 (.A1(net354),
    .A2(net257),
    .B1_N(net1040),
    .X(net372));
 sky130_fd_sc_hd__a31o_1 c609 (.A1(net352),
    .A2(net371),
    .A3(net1040),
    .B1(net744),
    .X(net373));
 sky130_fd_sc_hd__a21bo_1 c610 (.A1(net372),
    .A2(net611),
    .B1_N(net530),
    .X(net374));
 sky130_fd_sc_hd__mux4_1 c611 (.A0(net169),
    .A1(net685),
    .A2(net233),
    .A3(net365),
    .S0(net787),
    .S1(net221),
    .X(net375));
 sky130_fd_sc_hd__mux4_1 c612 (.A0(net366),
    .A1(net42),
    .A2(net1039),
    .A3(net57),
    .S0(net1021),
    .S1(net556),
    .X(net376));
 sky130_fd_sc_hd__clkbuf_1 c613 (.A(net547),
    .X(net377));
 sky130_fd_sc_hd__clkbuf_1 c614 (.A(net567),
    .X(net378));
 sky130_fd_sc_hd__a21bo_1 c615 (.A1(net239),
    .A2(net376),
    .B1_N(net557),
    .X(net379));
 sky130_fd_sc_hd__a41o_1 c616 (.A1(net1106),
    .A2(net1079),
    .A3(net668),
    .A4(net1057),
    .B1(net1040),
    .X(net380));
 sky130_fd_sc_hd__mux4_1 c617 (.A0(net223),
    .A1(net374),
    .A2(net581),
    .A3(net1121),
    .S0(net646),
    .S1(net1020),
    .X(net381));
 sky130_fd_sc_hd__clkbuf_1 c618 (.A(net564),
    .X(net683));
 sky130_fd_sc_hd__a41o_1 c619 (.A1(net285),
    .A2(net45),
    .A3(net1026),
    .A4(net670),
    .B1(net117),
    .X(net382));
 sky130_fd_sc_hd__mux4_1 c620 (.A0(net163),
    .A1(net269),
    .A2(net275),
    .A3(net669),
    .S0(net266),
    .S1(net1013),
    .X(net383));
 sky130_fd_sc_hd__a41o_1 c621 (.A1(net339),
    .A2(net381),
    .A3(net256),
    .A4(net1020),
    .B1(net223),
    .X(net384));
 sky130_fd_sc_hd__a41o_1 c622 (.A1(net331),
    .A2(net368),
    .A3(net672),
    .A4(net670),
    .B1(net1060),
    .X(net385));
 sky130_fd_sc_hd__a41o_1 c623 (.A1(net137),
    .A2(net1065),
    .A3(net1013),
    .A4(net269),
    .B1(net1049),
    .X(net386));
 sky130_fd_sc_hd__a31o_1 c624 (.A1(net170),
    .A2(net1042),
    .A3(net1104),
    .B1(net1044),
    .X(net387));
 sky130_fd_sc_hd__sdfbbn_1 c625 (.CLK_N(clknet_2_2__leaf_clk),
    .D(net173),
    .RESET_B(net1031),
    .SCD(net188),
    .SCE(net381),
    .SET_B(net557),
    .Q(net388));
 sky130_fd_sc_hd__a31o_1 c626 (.A1(net388),
    .A2(net116),
    .A3(net757),
    .B1(net546),
    .X(net389));
 sky130_fd_sc_hd__mux4_1 c627 (.A0(net340),
    .A1(net362),
    .A2(net646),
    .A3(net269),
    .S0(net1026),
    .S1(net542),
    .X(net390));
 sky130_fd_sc_hd__mux4_2 c628 (.A0(net356),
    .A1(net581),
    .A2(net1065),
    .A3(net1079),
    .S0(net368),
    .S1(net1026),
    .X(net391));
 sky130_fd_sc_hd__a21bo_1 c629 (.A1(net584),
    .A2(net291),
    .B1_N(net674),
    .X(net392));
 sky130_fd_sc_hd__mux4_1 c630 (.A0(net1055),
    .A1(net1040),
    .A2(net289),
    .A3(net1105),
    .S0(net1111),
    .S1(net556),
    .X(net393));
 sky130_fd_sc_hd__a41o_1 c631 (.A1(net353),
    .A2(net655),
    .A3(net1109),
    .A4(net170),
    .B1(net1033),
    .X(net394));
 sky130_fd_sc_hd__a41o_1 c632 (.A1(net393),
    .A2(net115),
    .A3(net390),
    .A4(net29),
    .B1(net1118),
    .X(net395));
 sky130_fd_sc_hd__a41o_1 c633 (.A1(net782),
    .A2(net1146),
    .A3(net389),
    .A4(net672),
    .B1(net392),
    .X(net396));
 sky130_fd_sc_hd__sdfbbn_1 c634 (.CLK_N(clknet_2_2__leaf_clk),
    .D(net575),
    .RESET_B(net1056),
    .SCD(net1101),
    .SCE(net285),
    .SET_B(net391),
    .Q(net398),
    .Q_N(net397));
 sky130_fd_sc_hd__mux4_2 c635 (.A0(net1109),
    .A1(net395),
    .A2(net284),
    .A3(net115),
    .S0(net397),
    .S1(net394),
    .X(net399));
 sky130_fd_sc_hd__sdfrbp_1 c636 (.CLK(clknet_2_2__leaf_clk),
    .D(net278),
    .RESET_B(net676),
    .SCD(net1044),
    .SCE(net829),
    .Q(net400));
 sky130_fd_sc_hd__mux4_1 c637 (.A0(net831),
    .A1(net816),
    .A2(net340),
    .A3(net399),
    .S0(net391),
    .S1(net1113),
    .X(net401));
 sky130_fd_sc_hd__xnor2_1 c660 (.A(net1122),
    .B(net106),
    .Y(net402));
 sky130_fd_sc_hd__xnor2_1 c661 (.A(net570),
    .B(net214),
    .Y(net403));
 sky130_fd_sc_hd__xnor2_2 c662 (.A(net1110),
    .B(net310),
    .Y(net404));
 sky130_fd_sc_hd__xnor2_1 c663 (.A(net214),
    .B(net1063),
    .Y(net405));
 sky130_fd_sc_hd__xnor2_1 c664 (.A(net756),
    .B(net214),
    .Y(net406));
 sky130_fd_sc_hd__xnor2_2 c665 (.A(net316),
    .B(net309),
    .Y(net407));
 sky130_fd_sc_hd__xnor2_1 c666 (.A(net303),
    .B(net1058),
    .Y(net408));
 sky130_fd_sc_hd__xnor2_2 c667 (.A(net1066),
    .B(net1058),
    .Y(net409));
 sky130_fd_sc_hd__a21bo_1 c668 (.A1(net211),
    .A2(net1132),
    .B1_N(net409),
    .X(net410));
 sky130_fd_sc_hd__a21bo_1 c669 (.A1(net408),
    .A2(net1120),
    .B1_N(net409),
    .X(net411));
 sky130_fd_sc_hd__xnor2_1 c670 (.A(net402),
    .B(net316),
    .Y(net412));
 sky130_fd_sc_hd__xnor2_1 c671 (.A(net407),
    .B(net115),
    .Y(net413));
 sky130_fd_sc_hd__a21bo_1 c672 (.A1(net409),
    .A2(net309),
    .B1_N(net407),
    .X(net414));
 sky130_fd_sc_hd__a21bo_1 c673 (.A1(net414),
    .A2(net413),
    .B1_N(net408),
    .X(net415));
 sky130_fd_sc_hd__mux4_1 c674 (.A0(net302),
    .A1(net303),
    .A2(net312),
    .A3(net1053),
    .S0(net410),
    .S1(net316),
    .X(net416));
 sky130_fd_sc_hd__xnor2_1 c675 (.A(net410),
    .B(net214),
    .Y(net417));
 sky130_fd_sc_hd__xnor2_1 c676 (.A(net403),
    .B(net414),
    .Y(net418));
 sky130_fd_sc_hd__clkbuf_1 c677 (.A(net544),
    .X(net419));
 sky130_fd_sc_hd__a31o_1 c678 (.A1(net414),
    .A2(net1064),
    .A3(net300),
    .B1(net207),
    .X(net420));
 sky130_fd_sc_hd__a31o_1 c679 (.A1(net405),
    .A2(net404),
    .A3(net1058),
    .B1(net414),
    .X(net421));
 sky130_fd_sc_hd__xnor2_1 c680 (.A(net417),
    .B(net416),
    .Y(net422));
 sky130_fd_sc_hd__clkbuf_1 c681 (.A(net544),
    .X(net423));
 sky130_fd_sc_hd__clkbuf_1 c682 (.A(net544),
    .X(net424));
 sky130_fd_sc_hd__buf_1 c683 (.A(net543),
    .X(net425));
 sky130_fd_sc_hd__xnor2_1 c684 (.A(net329),
    .B(net1078),
    .Y(net426));
 sky130_fd_sc_hd__a21bo_1 c685 (.A1(net106),
    .A2(net325),
    .B1_N(net1075),
    .X(net427));
 sky130_fd_sc_hd__xnor2_1 c686 (.A(net424),
    .B(net423),
    .Y(net428));
 sky130_fd_sc_hd__clkbuf_1 c687 (.A(net543),
    .X(net429));
 sky130_fd_sc_hd__a21bo_1 c688 (.A1(net324),
    .A2(net1122),
    .B1_N(net1027),
    .X(net430));
 sky130_fd_sc_hd__a21bo_1 c689 (.A1(net426),
    .A2(net1053),
    .B1_N(net427),
    .X(net431));
 sky130_fd_sc_hd__a21bo_1 c690 (.A1(net427),
    .A2(net314),
    .B1_N(net779),
    .X(net432));
 sky130_fd_sc_hd__xnor2_1 c691 (.A(net335),
    .B(net1061),
    .Y(net433));
 sky130_fd_sc_hd__a21bo_1 c692 (.A1(net428),
    .A2(net1027),
    .B1_N(net314),
    .X(net434));
 sky130_fd_sc_hd__xnor2_1 c693 (.A(net1046),
    .B(net429),
    .Y(net435));
 sky130_fd_sc_hd__xnor2_1 c694 (.A(net300),
    .B(net433),
    .Y(net436));
 sky130_fd_sc_hd__a21bo_1 c695 (.A1(net322),
    .A2(net409),
    .B1_N(net433),
    .X(net437));
 sky130_fd_sc_hd__a21bo_1 c696 (.A1(net416),
    .A2(net1123),
    .B1_N(net437),
    .X(net438));
 sky130_fd_sc_hd__a31o_1 c697 (.A1(net419),
    .A2(net317),
    .A3(net432),
    .B1(net409),
    .X(net439));
 sky130_fd_sc_hd__a21bo_1 c698 (.A1(net227),
    .A2(net1064),
    .B1_N(net425),
    .X(net440));
 sky130_fd_sc_hd__a31o_1 c699 (.A1(net435),
    .A2(net1017),
    .A3(net427),
    .B1(net439),
    .X(net441));
 sky130_fd_sc_hd__a21bo_1 c700 (.A1(net1065),
    .A2(net755),
    .B1_N(net437),
    .X(net442));
 sky130_fd_sc_hd__a21bo_1 c701 (.A1(net437),
    .A2(net317),
    .B1_N(net438),
    .X(net443));
 sky130_fd_sc_hd__a21bo_1 c702 (.A1(net105),
    .A2(net751),
    .B1_N(net438),
    .X(net444));
 sky130_fd_sc_hd__a31o_1 c703 (.A1(net436),
    .A2(net1113),
    .A3(net438),
    .B1(net442),
    .X(net445));
 sky130_fd_sc_hd__a21bo_1 c704 (.A1(net432),
    .A2(net427),
    .B1_N(net1026),
    .X(net446));
 sky130_fd_sc_hd__clkbuf_1 c705 (.A(net549),
    .X(net447));
 sky130_fd_sc_hd__clkbuf_1 c706 (.A(net548),
    .X(net448));
 sky130_fd_sc_hd__a21bo_1 c707 (.A1(net446),
    .A2(net1047),
    .B1_N(net1070),
    .X(net449));
 sky130_fd_sc_hd__mux4_1 c708 (.A0(net613),
    .A1(net417),
    .A2(net432),
    .A3(net438),
    .S0(net310),
    .S1(net666),
    .X(net450));
 sky130_fd_sc_hd__a21bo_1 c709 (.A1(net431),
    .A2(net403),
    .B1_N(net1012),
    .X(net451));
 sky130_fd_sc_hd__a21bo_1 c710 (.A1(net406),
    .A2(net1111),
    .B1_N(net335),
    .X(net452));
 sky130_fd_sc_hd__clkbuf_1 c711 (.A(net525),
    .X(net453));
 sky130_fd_sc_hd__a31o_1 c712 (.A1(net325),
    .A2(net301),
    .A3(net1075),
    .B1(net1016),
    .X(net454));
 sky130_fd_sc_hd__a21bo_1 c713 (.A1(net332),
    .A2(net121),
    .B1_N(net1112),
    .X(net455));
 sky130_fd_sc_hd__a21bo_1 c714 (.A1(net422),
    .A2(net425),
    .B1_N(net1111),
    .X(net456));
 sky130_fd_sc_hd__a21bo_1 c715 (.A1(net413),
    .A2(net135),
    .B1_N(net335),
    .X(net457));
 sky130_fd_sc_hd__a21bo_1 c716 (.A1(net207),
    .A2(net451),
    .B1_N(net1066),
    .X(net458));
 sky130_fd_sc_hd__clkbuf_1 c717 (.A(net524),
    .X(net459));
 sky130_fd_sc_hd__buf_1 c718 (.A(net565),
    .X(net460));
 sky130_fd_sc_hd__mux4_1 c719 (.A0(net460),
    .A1(net430),
    .A2(net791),
    .A3(net334),
    .S0(net60),
    .S1(net452),
    .X(net461));
 sky130_fd_sc_hd__a21bo_1 c720 (.A1(net358),
    .A2(net1061),
    .B1_N(net460),
    .X(net462));
 sky130_fd_sc_hd__mux4_1 c721 (.A0(net404),
    .A1(net448),
    .A2(net60),
    .A3(net256),
    .S0(net1046),
    .S1(net455),
    .X(net463));
 sky130_fd_sc_hd__a31o_1 c722 (.A1(net459),
    .A2(net440),
    .A3(net1061),
    .B1(net1026),
    .X(net464));
 sky130_fd_sc_hd__a31o_1 c723 (.A1(net449),
    .A2(net458),
    .A3(net464),
    .B1(net827),
    .X(net465));
 sky130_fd_sc_hd__mux4_1 c724 (.A0(net412),
    .A1(net464),
    .A2(net307),
    .A3(net1113),
    .S0(net445),
    .S1(net1081),
    .X(net466));
 sky130_fd_sc_hd__mux4_1 c725 (.A0(net315),
    .A1(net591),
    .A2(net460),
    .A3(net458),
    .S0(net532),
    .S1(net1081),
    .X(net467));
 sky130_fd_sc_hd__a21bo_1 c726 (.A1(net756),
    .A2(net439),
    .B1_N(net1112),
    .X(net468));
 sky130_fd_sc_hd__a31o_1 c727 (.A1(net263),
    .A2(net591),
    .A3(net1106),
    .B1(net1122),
    .X(net469));
 sky130_fd_sc_hd__a41o_1 c728 (.A1(net1017),
    .A2(net268),
    .A3(net341),
    .A4(net802),
    .B1(net1010),
    .X(net470));
 sky130_fd_sc_hd__sdfrbp_1 c729 (.CLK(clknet_2_1__leaf_clk),
    .D(net415),
    .RESET_B(net367),
    .SCD(net1070),
    .SCE(net434),
    .Q(net472),
    .Q_N(net471));
 sky130_fd_sc_hd__a31o_1 c730 (.A1(net762),
    .A2(net438),
    .A3(net367),
    .B1(net716),
    .X(net473));
 sky130_fd_sc_hd__mux4_1 c731 (.A0(net271),
    .A1(net1009),
    .A2(net471),
    .A3(net1109),
    .S0(net632),
    .S1(net1010),
    .X(net474));
 sky130_fd_sc_hd__a31o_1 c732 (.A1(net50),
    .A2(net104),
    .A3(net1017),
    .B1(net744),
    .X(net475));
 sky130_fd_sc_hd__a31o_1 c733 (.A1(net345),
    .A2(net442),
    .A3(net1026),
    .B1(net1075),
    .X(net476));
 sky130_fd_sc_hd__a21bo_1 c734 (.A1(net1070),
    .A2(net1122),
    .B1_N(net803),
    .X(net477));
 sky130_fd_sc_hd__a31o_1 c735 (.A1(net350),
    .A2(net1070),
    .A3(net535),
    .B1(net559),
    .X(net478));
 sky130_fd_sc_hd__a31o_1 c736 (.A1(net478),
    .A2(net773),
    .A3(net751),
    .B1(net549),
    .X(net479));
 sky130_fd_sc_hd__mux4_1 c737 (.A0(net472),
    .A1(net445),
    .A2(net442),
    .A3(net747),
    .S0(net462),
    .S1(net1061),
    .X(net480));
 sky130_fd_sc_hd__mux4_1 c738 (.A0(net420),
    .A1(net434),
    .A2(net781),
    .A3(net1120),
    .S0(net803),
    .S1(net1081),
    .X(net481));
 sky130_fd_sc_hd__clkbuf_1 c739 (.A(net566),
    .X(net482));
 sky130_fd_sc_hd__a31o_1 c740 (.A1(net781),
    .A2(net1109),
    .A3(net1069),
    .B1(net830),
    .X(net483));
 sky130_fd_sc_hd__mux4_1 c741 (.A0(net379),
    .A1(net468),
    .A2(net1122),
    .A3(net462),
    .S0(net349),
    .S1(net476),
    .X(net484));
 sky130_fd_sc_hd__a31o_1 c742 (.A1(net370),
    .A2(net453),
    .A3(net482),
    .B1(net1033),
    .X(net485));
 sky130_fd_sc_hd__a41o_1 c743 (.A1(net115),
    .A2(net84),
    .A3(net225),
    .A4(net574),
    .B1(net462),
    .X(net665));
 sky130_fd_sc_hd__a41o_1 c744 (.A1(net611),
    .A2(net479),
    .A3(net84),
    .A4(net442),
    .B1(net476),
    .X(net486));
 sky130_fd_sc_hd__a31o_1 c745 (.A1(net485),
    .A2(net788),
    .A3(net554),
    .B1(net1081),
    .X(net487));
 sky130_fd_sc_hd__a31o_1 c746 (.A1(net456),
    .A2(net450),
    .A3(net487),
    .B1(net529),
    .X(net488));
 sky130_fd_sc_hd__sdfbbp_1 c747 (.CLK(clknet_2_3__leaf_clk),
    .D(net1032),
    .RESET_B(net483),
    .SCD(net1021),
    .SCE(net266),
    .SET_B(net555),
    .Q(net490),
    .Q_N(net489));
 sky130_fd_sc_hd__mux4_1 c748 (.A0(net341),
    .A1(net1111),
    .A2(net386),
    .A3(net732),
    .S0(net1072),
    .S1(net716),
    .X(net491));
 sky130_fd_sc_hd__mux4_1 c749 (.A0(net447),
    .A1(net1077),
    .A2(net363),
    .A3(net402),
    .S0(net490),
    .S1(net1104),
    .X(net492));
 sky130_fd_sc_hd__mux4_2 c750 (.A0(net1068),
    .A1(net1033),
    .A2(net394),
    .A3(net1123),
    .S0(net533),
    .S1(net716),
    .X(net493));
 sky130_fd_sc_hd__mux4_2 c751 (.A0(net266),
    .A1(net1012),
    .A2(net1112),
    .A3(net1075),
    .S0(net441),
    .S1(net553),
    .X(net494));
 sky130_fd_sc_hd__mux4_1 c752 (.A0(net470),
    .A1(net359),
    .A2(net387),
    .A3(net587),
    .S0(net568),
    .S1(net828),
    .X(net495));
 sky130_fd_sc_hd__mux4_1 c753 (.A0(net632),
    .A1(net474),
    .A2(net1106),
    .A3(net489),
    .S0(net542),
    .S1(net1154),
    .X(net496));
 sky130_fd_sc_hd__mux4_1 c754 (.A0(net1101),
    .A1(net1064),
    .A2(net477),
    .A3(net492),
    .S0(net1120),
    .S1(net1075),
    .X(net497));
 sky130_fd_sc_hd__mux4_1 c755 (.A0(net1060),
    .A1(net1104),
    .A2(net723),
    .A3(net560),
    .S0(clknet_1_1__leaf_net561),
    .S1(clknet_1_1__leaf_net562),
    .X(net498));
 sky130_fd_sc_hd__mux4_1 c756 (.A0(net1044),
    .A1(net641),
    .A2(net122),
    .A3(net498),
    .S0(net1079),
    .S1(clknet_1_0__leaf_net561),
    .X(net499));
 sky130_fd_sc_hd__mux4_1 c757 (.A0(net284),
    .A1(net347),
    .A2(net225),
    .A3(net380),
    .S0(net751),
    .S1(net1021),
    .X(net500));
 sky130_fd_sc_hd__mux4_1 c758 (.A0(net210),
    .A1(net1126),
    .A2(net392),
    .A3(net1060),
    .S0(net1104),
    .S1(net558),
    .X(net501));
 sky130_fd_sc_hd__mux4_1 c759 (.A0(net491),
    .A1(net136),
    .A2(net469),
    .A3(net500),
    .S0(net1010),
    .S1(clknet_1_0__leaf_net562),
    .X(net502));
 sky130_fd_sc_hd__mux4_1 c760 (.A0(net441),
    .A1(net256),
    .A2(net399),
    .A3(net398),
    .S0(net774),
    .S1(net210),
    .X(net503));
 sky130_fd_sc_hd__mux4_1 c761 (.A0(net1013),
    .A1(net457),
    .A2(net499),
    .A3(net502),
    .S0(net1101),
    .S1(net535),
    .X(net504));
 sky130_fd_sc_hd__mux4_1 c762 (.A0(net411),
    .A1(net685),
    .A2(net378),
    .A3(net641),
    .S0(net1080),
    .S1(clknet_1_1__leaf_net563),
    .X(net505));
 sky130_fd_sc_hd__mux4_1 c763 (.A0(net791),
    .A1(net462),
    .A2(net475),
    .A3(net490),
    .S0(net36),
    .S1(clknet_1_0__leaf_net563),
    .X(net506));
 sky130_fd_sc_hd__mux4_2 c764 (.A0(net28),
    .A1(net391),
    .A2(net493),
    .A3(net590),
    .S0(net398),
    .S1(net545),
    .X(net507));
 sky130_fd_sc_hd__mux4_1 c765 (.A0(clknet_1_0__leaf_net506),
    .A1(net1104),
    .A2(net60),
    .A3(net396),
    .S0(net210),
    .S1(net574),
    .X(net508));
 sky130_fd_sc_hd__mux4_1 c766 (.A0(net279),
    .A1(net1010),
    .A2(net590),
    .A3(net136),
    .S0(net751),
    .S1(net555),
    .X(net509));
 sky130_fd_sc_hd__mux4_1 c767 (.A0(net454),
    .A1(net501),
    .A2(net509),
    .A3(net1026),
    .S0(net546),
    .S1(net559),
    .X(net510));
 sky130_fd_sc_hd__mux4_1 c768 (.A0(net505),
    .A1(net275),
    .A2(net377),
    .A3(net587),
    .S0(clknet_1_1__leaf_net506),
    .X(net511));
 sky130_fd_sc_hd__mux4_2 c769 (.A0(net342),
    .A1(net280),
    .A2(net510),
    .A3(net507),
    .S0(net545),
    .S1(net551),
    .X(net512));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net506 (.A(net506),
    .X(clknet_0_net506));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net561 (.A(net561),
    .X(clknet_0_net561));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net562 (.A(net562),
    .X(clknet_0_net562));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net563 (.A(net563),
    .X(clknet_0_net563));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net506 (.A(clknet_0_net506),
    .X(clknet_1_0__leaf_net506));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net561 (.A(clknet_0_net561),
    .X(clknet_1_0__leaf_net561));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net562 (.A(clknet_0_net562),
    .X(clknet_1_0__leaf_net562));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net563 (.A(clknet_0_net563),
    .X(clknet_1_0__leaf_net563));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net506 (.A(clknet_0_net506),
    .X(clknet_1_1__leaf_net506));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net561 (.A(clknet_0_net561),
    .X(clknet_1_1__leaf_net561));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net562 (.A(clknet_0_net562),
    .X(clknet_1_1__leaf_net562));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net563 (.A(clknet_0_net563),
    .X(clknet_1_1__leaf_net563));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_2 clone22 (.A(net1141),
    .X(net791));
 sky130_fd_sc_hd__buf_1 clone5 (.A(net780),
    .X(net774));
 sky130_fd_sc_hd__clkbuf_1 fanout175 (.A(net1026),
    .X(net740));
 sky130_fd_sc_hd__clkbuf_1 fanout176 (.A(net707),
    .X(net741));
 sky130_fd_sc_hd__clkbuf_1 fanout178 (.A(net1031),
    .X(net743));
 sky130_fd_sc_hd__clkbuf_2 fanout179 (.A(net1031),
    .X(net744));
 sky130_fd_sc_hd__buf_1 fanout180 (.A(net667),
    .X(net745));
 sky130_fd_sc_hd__buf_6 fanout181 (.A(net1038),
    .X(net746));
 sky130_fd_sc_hd__buf_6 fanout182 (.A(net119),
    .X(net747));
 sky130_fd_sc_hd__clkbuf_1 fanout203 (.A(net1090),
    .X(net768));
 sky130_fd_sc_hd__clkbuf_1 fanout204 (.A(net588),
    .X(net769));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(net1081),
    .X(net827));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(net560),
    .X(net828));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(net539),
    .X(net829));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(net530),
    .X(net830));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(net400),
    .X(net831));
 sky130_fd_sc_hd__clkbuf_8 input1 (.A(net832),
    .X(net519));
 sky130_fd_sc_hd__buf_2 input10 (.A(net841),
    .X(net575));
 sky130_fd_sc_hd__buf_6 input11 (.A(net842),
    .X(net576));
 sky130_fd_sc_hd__buf_4 input12 (.A(net843),
    .X(net577));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(net844),
    .X(net578));
 sky130_fd_sc_hd__clkbuf_8 input14 (.A(net845),
    .X(net579));
 sky130_fd_sc_hd__buf_6 input15 (.A(net846),
    .X(net580));
 sky130_fd_sc_hd__clkbuf_2 input16 (.A(net847),
    .X(net581));
 sky130_fd_sc_hd__dlymetal6s2s_1 input17 (.A(net848),
    .X(net582));
 sky130_fd_sc_hd__clkbuf_2 input18 (.A(net849),
    .X(net583));
 sky130_fd_sc_hd__buf_2 input19 (.A(net850),
    .X(net584));
 sky130_fd_sc_hd__buf_1 input2 (.A(net833),
    .X(net550));
 sky130_fd_sc_hd__buf_6 input20 (.A(net851),
    .X(net585));
 sky130_fd_sc_hd__clkbuf_2 input21 (.A(net852),
    .X(net586));
 sky130_fd_sc_hd__buf_2 input22 (.A(net853),
    .X(net587));
 sky130_fd_sc_hd__clkbuf_1 input23 (.A(net854),
    .X(net588));
 sky130_fd_sc_hd__clkbuf_2 input24 (.A(net855),
    .X(net589));
 sky130_fd_sc_hd__buf_1 input25 (.A(net856),
    .X(net590));
 sky130_fd_sc_hd__clkbuf_2 input26 (.A(net857),
    .X(net591));
 sky130_fd_sc_hd__clkbuf_1 input27 (.A(net858),
    .X(net592));
 sky130_fd_sc_hd__clkbuf_4 input28 (.A(net859),
    .X(net593));
 sky130_fd_sc_hd__clkbuf_2 input29 (.A(net860),
    .X(net594));
 sky130_fd_sc_hd__buf_6 input3 (.A(net834),
    .X(net568));
 sky130_fd_sc_hd__buf_4 input30 (.A(net861),
    .X(net595));
 sky130_fd_sc_hd__clkbuf_1 input31 (.A(net862),
    .X(net596));
 sky130_fd_sc_hd__buf_2 input32 (.A(net863),
    .X(net597));
 sky130_fd_sc_hd__buf_1 input33 (.A(net864),
    .X(net598));
 sky130_fd_sc_hd__clkbuf_4 input34 (.A(net865),
    .X(net599));
 sky130_fd_sc_hd__buf_8 input35 (.A(net866),
    .X(net600));
 sky130_fd_sc_hd__clkbuf_4 input36 (.A(net867),
    .X(net601));
 sky130_fd_sc_hd__buf_2 input37 (.A(net868),
    .X(net602));
 sky130_fd_sc_hd__clkbuf_4 input38 (.A(net869),
    .X(net603));
 sky130_fd_sc_hd__clkbuf_2 input39 (.A(net870),
    .X(net604));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(net835),
    .X(net569));
 sky130_fd_sc_hd__dlymetal6s2s_1 input40 (.A(net871),
    .X(net605));
 sky130_fd_sc_hd__clkbuf_2 input41 (.A(net872),
    .X(net606));
 sky130_fd_sc_hd__clkbuf_4 input42 (.A(net873),
    .X(net607));
 sky130_fd_sc_hd__buf_2 input43 (.A(net874),
    .X(net608));
 sky130_fd_sc_hd__buf_2 input44 (.A(net875),
    .X(net609));
 sky130_fd_sc_hd__dlymetal6s2s_1 input45 (.A(net876),
    .X(net610));
 sky130_fd_sc_hd__buf_4 input46 (.A(net877),
    .X(net611));
 sky130_fd_sc_hd__clkbuf_1 input47 (.A(net878),
    .X(net612));
 sky130_fd_sc_hd__buf_2 input48 (.A(net879),
    .X(net613));
 sky130_fd_sc_hd__clkbuf_2 input49 (.A(net880),
    .X(net614));
 sky130_fd_sc_hd__buf_4 input5 (.A(net836),
    .X(net570));
 sky130_fd_sc_hd__clkbuf_2 input50 (.A(net881),
    .X(net615));
 sky130_fd_sc_hd__buf_2 input51 (.A(net882),
    .X(net616));
 sky130_fd_sc_hd__clkbuf_1 input52 (.A(net883),
    .X(net617));
 sky130_fd_sc_hd__clkbuf_2 input53 (.A(net884),
    .X(net618));
 sky130_fd_sc_hd__clkbuf_1 input54 (.A(net885),
    .X(net619));
 sky130_fd_sc_hd__buf_2 input55 (.A(net886),
    .X(net620));
 sky130_fd_sc_hd__buf_2 input56 (.A(net887),
    .X(net621));
 sky130_fd_sc_hd__buf_1 input57 (.A(net888),
    .X(net622));
 sky130_fd_sc_hd__buf_4 input58 (.A(net889),
    .X(net623));
 sky130_fd_sc_hd__clkbuf_2 input59 (.A(net890),
    .X(net624));
 sky130_fd_sc_hd__buf_2 input6 (.A(net837),
    .X(net571));
 sky130_fd_sc_hd__buf_1 input60 (.A(net891),
    .X(net625));
 sky130_fd_sc_hd__clkbuf_2 input61 (.A(net892),
    .X(net626));
 sky130_fd_sc_hd__buf_2 input62 (.A(net893),
    .X(net627));
 sky130_fd_sc_hd__clkbuf_2 input63 (.A(net894),
    .X(net628));
 sky130_fd_sc_hd__buf_1 input64 (.A(net895),
    .X(net629));
 sky130_fd_sc_hd__buf_1 input65 (.A(net896),
    .X(net630));
 sky130_fd_sc_hd__clkbuf_1 input66 (.A(net897),
    .X(net631));
 sky130_fd_sc_hd__clkbuf_4 input67 (.A(net898),
    .X(net632));
 sky130_fd_sc_hd__clkbuf_8 input68 (.A(net899),
    .X(net633));
 sky130_fd_sc_hd__clkbuf_1 input69 (.A(net900),
    .X(net634));
 sky130_fd_sc_hd__buf_6 input7 (.A(net838),
    .X(net572));
 sky130_fd_sc_hd__buf_2 input70 (.A(net901),
    .X(net635));
 sky130_fd_sc_hd__clkbuf_2 input71 (.A(net902),
    .X(net636));
 sky130_fd_sc_hd__dlymetal6s2s_1 input72 (.A(net903),
    .X(net637));
 sky130_fd_sc_hd__buf_1 input73 (.A(net904),
    .X(net638));
 sky130_fd_sc_hd__clkbuf_2 input74 (.A(net905),
    .X(net639));
 sky130_fd_sc_hd__clkbuf_1 input75 (.A(net906),
    .X(net640));
 sky130_fd_sc_hd__buf_2 input76 (.A(net907),
    .X(net641));
 sky130_fd_sc_hd__buf_1 input77 (.A(net908),
    .X(net642));
 sky130_fd_sc_hd__dlymetal6s2s_1 input78 (.A(net909),
    .X(net643));
 sky130_fd_sc_hd__buf_4 input79 (.A(net910),
    .X(net644));
 sky130_fd_sc_hd__buf_6 input8 (.A(net839),
    .X(net573));
 sky130_fd_sc_hd__clkbuf_4 input80 (.A(net911),
    .X(net645));
 sky130_fd_sc_hd__clkbuf_2 input81 (.A(net912),
    .X(net646));
 sky130_fd_sc_hd__dlymetal6s2s_1 input82 (.A(net913),
    .X(net647));
 sky130_fd_sc_hd__clkbuf_2 input83 (.A(net914),
    .X(net648));
 sky130_fd_sc_hd__buf_1 input84 (.A(net915),
    .X(net649));
 sky130_fd_sc_hd__clkbuf_2 input85 (.A(net916),
    .X(net650));
 sky130_fd_sc_hd__clkbuf_2 input86 (.A(net917),
    .X(net651));
 sky130_fd_sc_hd__clkbuf_2 input87 (.A(net918),
    .X(net652));
 sky130_fd_sc_hd__clkbuf_1 input88 (.A(net919),
    .X(net653));
 sky130_fd_sc_hd__buf_1 input89 (.A(net920),
    .X(net654));
 sky130_fd_sc_hd__buf_6 input9 (.A(net840),
    .X(net574));
 sky130_fd_sc_hd__clkbuf_2 input90 (.A(net921),
    .X(net655));
 sky130_fd_sc_hd__clkbuf_1 input91 (.A(net922),
    .X(net656));
 sky130_fd_sc_hd__buf_1 input92 (.A(net923),
    .X(net657));
 sky130_fd_sc_hd__buf_1 input93 (.A(net924),
    .X(net658));
 sky130_fd_sc_hd__clkbuf_4 input94 (.A(net925),
    .X(net659));
 sky130_fd_sc_hd__buf_1 input95 (.A(net926),
    .X(net660));
 sky130_fd_sc_hd__clkbuf_1 input96 (.A(net927),
    .X(net661));
 sky130_fd_sc_hd__clkbuf_2 input97 (.A(net928),
    .X(net662));
 sky130_fd_sc_hd__buf_2 input98 (.A(net929),
    .X(net663));
 sky130_fd_sc_hd__buf_1 input99 (.A(net930),
    .X(net664));
 sky130_fd_sc_hd__buf_6 max_cap177 (.A(net221),
    .X(net742));
 sky130_fd_sc_hd__buf_6 max_cap183 (.A(net749),
    .X(net748));
 sky130_fd_sc_hd__buf_4 max_cap184 (.A(net202),
    .X(net749));
 sky130_fd_sc_hd__buf_6 max_cap185 (.A(net102),
    .X(net750));
 sky130_fd_sc_hd__buf_4 max_cap186 (.A(net752),
    .X(net751));
 sky130_fd_sc_hd__buf_4 max_cap187 (.A(net681),
    .X(net752));
 sky130_fd_sc_hd__buf_4 max_cap188 (.A(net132),
    .X(net753));
 sky130_fd_sc_hd__buf_4 max_cap190 (.A(net120),
    .X(net755));
 sky130_fd_sc_hd__clkbuf_2 max_cap192 (.A(net21),
    .X(net757));
 sky130_fd_sc_hd__buf_4 max_cap193 (.A(net86),
    .X(net758));
 sky130_fd_sc_hd__buf_4 max_cap194 (.A(net1066),
    .X(net759));
 sky130_fd_sc_hd__buf_4 max_cap195 (.A(net103),
    .X(net760));
 sky130_fd_sc_hd__buf_4 max_cap196 (.A(net33),
    .X(net761));
 sky130_fd_sc_hd__buf_8 max_cap197 (.A(net14),
    .X(net762));
 sky130_fd_sc_hd__buf_4 max_cap198 (.A(net1091),
    .X(net763));
 sky130_fd_sc_hd__buf_6 max_cap199 (.A(net98),
    .X(net764));
 sky130_fd_sc_hd__buf_6 max_cap200 (.A(net738),
    .X(net765));
 sky130_fd_sc_hd__buf_4 max_cap201 (.A(net13),
    .X(net766));
 sky130_fd_sc_hd__clkbuf_2 max_cap202 (.A(net699),
    .X(net767));
 sky130_fd_sc_hd__a41o_1 merge782 (.A1(net418),
    .A2(net303),
    .A3(net421),
    .A4(net411),
    .B1(net422),
    .X(net513));
 sky130_fd_sc_hd__a31o_1 merge783 (.A1(net167),
    .A2(net793),
    .A3(net145),
    .B1(net175),
    .X(net514));
 sky130_fd_sc_hd__mux4_1 merge784 (.A0(net99),
    .A1(net418),
    .A2(net217),
    .A3(net406),
    .S0(net420),
    .S1(net1007),
    .X(net515));
 sky130_fd_sc_hd__mux4_1 merge785 (.A0(net281),
    .A1(net192),
    .A2(net189),
    .A3(net288),
    .S0(net195),
    .S1(net276),
    .X(net516));
 sky130_fd_sc_hd__mux4_1 merge786 (.A0(net357),
    .A1(net616),
    .A2(net352),
    .A3(net164),
    .S0(net814),
    .S1(net744),
    .X(net517));
 sky130_fd_sc_hd__a31o_1 merge787 (.A1(net595),
    .A2(net175),
    .A3(net176),
    .B1(net1024),
    .X(net518));
 sky130_fd_sc_hd__a41o_4 merge788 (.A1(net344),
    .A2(net338),
    .A3(net328),
    .A4(net216),
    .X(net540));
 sky130_fd_sc_hd__mux4_1 merge789 (.A0(net407),
    .A1(net334),
    .A2(net613),
    .A3(net443),
    .S0(net442),
    .S1(net1128),
    .X(net520));
 sky130_fd_sc_hd__mux4_1 merge790 (.A0(net258),
    .A1(net686),
    .A2(net641),
    .A3(net222),
    .S0(net260),
    .S1(net632),
    .X(net521));
 sky130_fd_sc_hd__mux4_1 merge791 (.A0(net425),
    .A1(net407),
    .A2(net415),
    .A3(net206),
    .S0(net815),
    .S1(net589),
    .X(net522));
 sky130_fd_sc_hd__mux4_1 merge792 (.A0(net147),
    .A1(net360),
    .A2(net676),
    .A3(net591),
    .S0(net365),
    .S1(net1118),
    .X(net523));
 sky130_fd_sc_hd__sdfbbn_1 merge793 (.CLK_N(clknet_2_1__leaf_clk),
    .D(net252),
    .RESET_B(net106),
    .SCD(net587),
    .SCE(net452),
    .SET_B(net444),
    .Q(net525),
    .Q_N(net524));
 sky130_fd_sc_hd__mux4_1 merge794 (.A0(net191),
    .A1(net1094),
    .A2(net1031),
    .A3(net180),
    .S0(net575),
    .S1(net663),
    .X(net526));
 sky130_fd_sc_hd__mux4_1 merge795 (.A0(net455),
    .A1(net312),
    .A2(net791),
    .A3(net193),
    .S0(net282),
    .S1(net290),
    .X(net527));
 sky130_fd_sc_hd__mux4_1 merge796 (.A0(net1062),
    .A1(net216),
    .A2(net814),
    .A3(net237),
    .S0(net476),
    .S1(net457),
    .X(net528));
 sky130_fd_sc_hd__dfrbp_1 merge797 (.CLK(clknet_2_1__leaf_clk),
    .D(net373),
    .RESET_B(net369),
    .Q(net530),
    .Q_N(net529));
 sky130_fd_sc_hd__xnor2_1 merge798 (.A(net197),
    .B(net526),
    .Y(net531));
 sky130_fd_sc_hd__dfrbp_1 merge799 (.CLK(clknet_2_0__leaf_clk),
    .D(net461),
    .RESET_B(net465),
    .Q(net533),
    .Q_N(net532));
 sky130_fd_sc_hd__xnor2_2 merge800 (.A(net514),
    .B(net521),
    .Y(net534));
 sky130_fd_sc_hd__dfrtn_1 merge801 (.CLK_N(clknet_2_1__leaf_clk),
    .D(net473),
    .RESET_B(net480),
    .Q(net535));
 sky130_fd_sc_hd__xnor2_2 merge802 (.A(net512),
    .B(net494),
    .Y(net536));
 sky130_fd_sc_hd__xnor2_1 merge803 (.A(net515),
    .B(net522),
    .Y(net537));
 sky130_fd_sc_hd__xnor2_1 merge804 (.A(net287),
    .B(net295),
    .Y(net538));
 sky130_fd_sc_hd__dfrtp_1 merge805 (.CLK(clknet_2_2__leaf_clk),
    .D(net382),
    .RESET_B(net383),
    .Q(net539));
 sky130_fd_sc_hd__dfrtp_4 merge806 (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net337),
    .Q(net540));
 sky130_fd_sc_hd__dfrtp_1 merge807 (.CLK(clknet_2_2__leaf_clk),
    .D(net518),
    .RESET_B(net531),
    .Q(net714));
 sky130_fd_sc_hd__dfsbp_2 merge808 (.CLK(clknet_2_2__leaf_clk),
    .D(net294),
    .SET_B(net516),
    .Q(net542),
    .Q_N(net541));
 sky130_fd_sc_hd__dfsbp_1 merge809 (.CLK(clknet_2_1__leaf_clk),
    .D(net513),
    .SET_B(net537),
    .Q(net544),
    .Q_N(net543));
 sky130_fd_sc_hd__dfstp_1 merge810 (.CLK(clknet_2_3__leaf_clk),
    .D(net536),
    .SET_B(net495),
    .Q(net545));
 sky130_fd_sc_hd__dfstp_1 merge811 (.CLK(clknet_2_3__leaf_clk),
    .D(net384),
    .SET_B(net385),
    .Q(net546));
 sky130_fd_sc_hd__dfstp_1 merge812 (.CLK(clknet_2_3__leaf_clk),
    .D(net517),
    .SET_B(net523),
    .Q(net547));
 sky130_fd_sc_hd__dlrbn_1 merge813 (.D(net466),
    .GATE_N(clknet_2_1__leaf_clk),
    .RESET_B(net520),
    .Q(net549),
    .Q_N(net548));
 sky130_fd_sc_hd__dlrbn_1 merge814 (.GATE_N(clknet_2_3__leaf_clk),
    .RESET_B(net508),
    .Q(net551),
    .Q_N(net511));
 sky130_fd_sc_hd__dlrbp_2 merge815 (.D(net538),
    .GATE(clknet_2_2__leaf_clk),
    .RESET_B(net534),
    .Q(net680),
    .Q_N(net552));
 sky130_fd_sc_hd__dlrbp_1 merge816 (.D(net481),
    .GATE(clknet_2_0__leaf_clk),
    .RESET_B(net486),
    .Q(net554),
    .Q_N(net553));
 sky130_fd_sc_hd__dlrtn_1 merge817 (.D(net488),
    .GATE_N(clknet_2_3__leaf_clk),
    .RESET_B(net504),
    .Q(net555));
 sky130_fd_sc_hd__clkbuf_1 output100 (.A(net665),
    .X(net931));
 sky130_fd_sc_hd__clkbuf_1 output101 (.A(net666),
    .X(net932));
 sky130_fd_sc_hd__clkbuf_1 output102 (.A(net745),
    .X(net933));
 sky130_fd_sc_hd__clkbuf_1 output103 (.A(net668),
    .X(net934));
 sky130_fd_sc_hd__clkbuf_1 output104 (.A(net669),
    .X(net935));
 sky130_fd_sc_hd__clkbuf_1 output105 (.A(net670),
    .X(net936));
 sky130_fd_sc_hd__clkbuf_1 output106 (.A(net671),
    .X(net937));
 sky130_fd_sc_hd__clkbuf_1 output107 (.A(net672),
    .X(net938));
 sky130_fd_sc_hd__clkbuf_1 output108 (.A(net673),
    .X(net939));
 sky130_fd_sc_hd__clkbuf_1 output109 (.A(net674),
    .X(net940));
 sky130_fd_sc_hd__clkbuf_1 output110 (.A(net675),
    .X(net941));
 sky130_fd_sc_hd__clkbuf_1 output111 (.A(net676),
    .X(net942));
 sky130_fd_sc_hd__clkbuf_1 output112 (.A(net677),
    .X(net943));
 sky130_fd_sc_hd__clkbuf_1 output113 (.A(net678),
    .X(net944));
 sky130_fd_sc_hd__clkbuf_1 output114 (.A(net679),
    .X(net945));
 sky130_fd_sc_hd__clkbuf_1 output115 (.A(net680),
    .X(net946));
 sky130_fd_sc_hd__clkbuf_1 output116 (.A(net1058),
    .X(net947));
 sky130_fd_sc_hd__clkbuf_1 output117 (.A(net1049),
    .X(net948));
 sky130_fd_sc_hd__clkbuf_1 output118 (.A(net683),
    .X(net949));
 sky130_fd_sc_hd__clkbuf_1 output119 (.A(net684),
    .X(net950));
 sky130_fd_sc_hd__clkbuf_1 output120 (.A(net1054),
    .X(net951));
 sky130_fd_sc_hd__clkbuf_1 output121 (.A(net686),
    .X(net952));
 sky130_fd_sc_hd__clkbuf_1 output122 (.A(net687),
    .X(net953));
 sky130_fd_sc_hd__clkbuf_1 output123 (.A(net688),
    .X(net954));
 sky130_fd_sc_hd__clkbuf_1 output124 (.A(net689),
    .X(net955));
 sky130_fd_sc_hd__clkbuf_1 output125 (.A(net690),
    .X(net956));
 sky130_fd_sc_hd__clkbuf_1 output126 (.A(net691),
    .X(net957));
 sky130_fd_sc_hd__clkbuf_1 output127 (.A(net692),
    .X(net958));
 sky130_fd_sc_hd__clkbuf_1 output128 (.A(net693),
    .X(net959));
 sky130_fd_sc_hd__clkbuf_1 output129 (.A(net694),
    .X(net960));
 sky130_fd_sc_hd__clkbuf_1 output130 (.A(net695),
    .X(net961));
 sky130_fd_sc_hd__clkbuf_1 output131 (.A(net696),
    .X(net962));
 sky130_fd_sc_hd__clkbuf_1 output132 (.A(net1071),
    .X(net963));
 sky130_fd_sc_hd__clkbuf_1 output133 (.A(net777),
    .X(net964));
 sky130_fd_sc_hd__clkbuf_1 output134 (.A(net699),
    .X(net965));
 sky130_fd_sc_hd__clkbuf_1 output135 (.A(net700),
    .X(net966));
 sky130_fd_sc_hd__clkbuf_1 output136 (.A(net701),
    .X(net967));
 sky130_fd_sc_hd__clkbuf_1 output137 (.A(net702),
    .X(net968));
 sky130_fd_sc_hd__clkbuf_1 output138 (.A(net703),
    .X(net969));
 sky130_fd_sc_hd__clkbuf_1 output139 (.A(net704),
    .X(net970));
 sky130_fd_sc_hd__clkbuf_1 output140 (.A(net705),
    .X(net971));
 sky130_fd_sc_hd__clkbuf_1 output141 (.A(net706),
    .X(net972));
 sky130_fd_sc_hd__clkbuf_1 output142 (.A(net1026),
    .X(net973));
 sky130_fd_sc_hd__clkbuf_1 output143 (.A(net708),
    .X(net974));
 sky130_fd_sc_hd__clkbuf_1 output144 (.A(net709),
    .X(net975));
 sky130_fd_sc_hd__clkbuf_1 output145 (.A(net710),
    .X(net976));
 sky130_fd_sc_hd__clkbuf_1 output146 (.A(net1048),
    .X(net977));
 sky130_fd_sc_hd__clkbuf_1 output147 (.A(net712),
    .X(net978));
 sky130_fd_sc_hd__clkbuf_1 output148 (.A(net1088),
    .X(net979));
 sky130_fd_sc_hd__clkbuf_1 output149 (.A(net714),
    .X(net980));
 sky130_fd_sc_hd__clkbuf_1 output150 (.A(net715),
    .X(net981));
 sky130_fd_sc_hd__clkbuf_1 output151 (.A(net716),
    .X(net982));
 sky130_fd_sc_hd__clkbuf_1 output152 (.A(net717),
    .X(net983));
 sky130_fd_sc_hd__clkbuf_1 output153 (.A(net718),
    .X(net984));
 sky130_fd_sc_hd__clkbuf_1 output154 (.A(net719),
    .X(net985));
 sky130_fd_sc_hd__clkbuf_1 output155 (.A(net720),
    .X(net986));
 sky130_fd_sc_hd__clkbuf_1 output156 (.A(net721),
    .X(net987));
 sky130_fd_sc_hd__clkbuf_1 output157 (.A(net722),
    .X(net988));
 sky130_fd_sc_hd__clkbuf_1 output158 (.A(net1020),
    .X(net989));
 sky130_fd_sc_hd__clkbuf_1 output159 (.A(net724),
    .X(net990));
 sky130_fd_sc_hd__clkbuf_1 output160 (.A(net725),
    .X(net991));
 sky130_fd_sc_hd__clkbuf_1 output161 (.A(net1087),
    .X(net992));
 sky130_fd_sc_hd__clkbuf_1 output162 (.A(net727),
    .X(net993));
 sky130_fd_sc_hd__clkbuf_1 output163 (.A(net728),
    .X(net994));
 sky130_fd_sc_hd__clkbuf_1 output164 (.A(net729),
    .X(net995));
 sky130_fd_sc_hd__clkbuf_1 output165 (.A(net730),
    .X(net996));
 sky130_fd_sc_hd__clkbuf_1 output166 (.A(net731),
    .X(net997));
 sky130_fd_sc_hd__clkbuf_1 output167 (.A(net1066),
    .X(net998));
 sky130_fd_sc_hd__clkbuf_1 output168 (.A(net733),
    .X(net999));
 sky130_fd_sc_hd__clkbuf_1 output169 (.A(net822),
    .X(net1000));
 sky130_fd_sc_hd__clkbuf_1 output170 (.A(net735),
    .X(net1001));
 sky130_fd_sc_hd__clkbuf_1 output171 (.A(net736),
    .X(net1002));
 sky130_fd_sc_hd__clkbuf_1 output172 (.A(net737),
    .X(net1003));
 sky130_fd_sc_hd__clkbuf_1 output173 (.A(net765),
    .X(net1004));
 sky130_fd_sc_hd__clkbuf_1 output174 (.A(net739),
    .X(net1005));
 sky130_fd_sc_hd__clkbuf_2 rebuffer1 (.A(net738),
    .X(net770));
 sky130_fd_sc_hd__buf_1 rebuffer10 (.A(net778),
    .X(net779));
 sky130_fd_sc_hd__buf_1 rebuffer11 (.A(net778),
    .X(net780));
 sky130_fd_sc_hd__clkbuf_2 rebuffer12 (.A(net817),
    .X(net781));
 sky130_fd_sc_hd__clkbuf_1 rebuffer13 (.A(net59),
    .X(net782));
 sky130_fd_sc_hd__clkbuf_1 rebuffer14 (.A(net59),
    .X(net783));
 sky130_fd_sc_hd__buf_1 rebuffer15 (.A(net23),
    .X(net784));
 sky130_fd_sc_hd__buf_1 rebuffer16 (.A(net76),
    .X(net785));
 sky130_fd_sc_hd__buf_1 rebuffer17 (.A(net76),
    .X(net786));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer18 (.A(net786),
    .X(net787));
 sky130_fd_sc_hd__clkbuf_1 rebuffer19 (.A(net787),
    .X(net788));
 sky130_fd_sc_hd__buf_1 rebuffer2 (.A(net738),
    .X(net771));
 sky130_fd_sc_hd__buf_2 rebuffer20 (.A(net43),
    .X(net789));
 sky130_fd_sc_hd__clkbuf_1 rebuffer21 (.A(net789),
    .X(net790));
 sky130_fd_sc_hd__buf_1 rebuffer23 (.A(net804),
    .X(net792));
 sky130_fd_sc_hd__clkbuf_1 rebuffer24 (.A(net1135),
    .X(net793));
 sky130_fd_sc_hd__clkbuf_1 rebuffer25 (.A(net793),
    .X(net794));
 sky130_fd_sc_hd__clkbuf_1 rebuffer26 (.A(net247),
    .X(net795));
 sky130_fd_sc_hd__buf_2 rebuffer27 (.A(net742),
    .X(net796));
 sky130_fd_sc_hd__clkbuf_1 rebuffer28 (.A(net796),
    .X(net797));
 sky130_fd_sc_hd__buf_2 rebuffer29 (.A(net201),
    .X(net798));
 sky130_fd_sc_hd__buf_4 rebuffer3 (.A(net14),
    .X(net772));
 sky130_fd_sc_hd__clkbuf_1 rebuffer30 (.A(net798),
    .X(net799));
 sky130_fd_sc_hd__buf_1 rebuffer31 (.A(net63),
    .X(net800));
 sky130_fd_sc_hd__clkbuf_1 rebuffer32 (.A(net800),
    .X(net801));
 sky130_fd_sc_hd__clkbuf_1 rebuffer33 (.A(net1009),
    .X(net802));
 sky130_fd_sc_hd__buf_1 rebuffer34 (.A(net1009),
    .X(net803));
 sky130_fd_sc_hd__clkbuf_1 rebuffer35 (.A(net805),
    .X(net804));
 sky130_fd_sc_hd__clkbuf_1 rebuffer36 (.A(net806),
    .X(net805));
 sky130_fd_sc_hd__clkbuf_1 rebuffer37 (.A(net807),
    .X(net806));
 sky130_fd_sc_hd__clkbuf_1 rebuffer38 (.A(net808),
    .X(net807));
 sky130_fd_sc_hd__clkbuf_1 rebuffer39 (.A(net809),
    .X(net808));
 sky130_fd_sc_hd__buf_1 rebuffer4 (.A(net1157),
    .X(net773));
 sky130_fd_sc_hd__clkbuf_1 rebuffer40 (.A(net810),
    .X(net809));
 sky130_fd_sc_hd__clkbuf_1 rebuffer41 (.A(net811),
    .X(net810));
 sky130_fd_sc_hd__clkbuf_1 rebuffer42 (.A(net812),
    .X(net811));
 sky130_fd_sc_hd__buf_1 rebuffer43 (.A(net1150),
    .X(net812));
 sky130_fd_sc_hd__clkbuf_1 rebuffer44 (.A(net1142),
    .X(net813));
 sky130_fd_sc_hd__buf_1 rebuffer45 (.A(net1161),
    .X(net814));
 sky130_fd_sc_hd__clkbuf_1 rebuffer46 (.A(net1161),
    .X(net815));
 sky130_fd_sc_hd__clkbuf_1 rebuffer47 (.A(net283),
    .X(net816));
 sky130_fd_sc_hd__clkbuf_1 rebuffer48 (.A(net818),
    .X(net817));
 sky130_fd_sc_hd__clkbuf_1 rebuffer49 (.A(net819),
    .X(net818));
 sky130_fd_sc_hd__clkbuf_1 rebuffer50 (.A(net820),
    .X(net819));
 sky130_fd_sc_hd__clkbuf_1 rebuffer51 (.A(net821),
    .X(net820));
 sky130_fd_sc_hd__clkbuf_1 rebuffer52 (.A(net1149),
    .X(net821));
 sky130_fd_sc_hd__buf_1 rebuffer53 (.A(net734),
    .X(net822));
 sky130_fd_sc_hd__clkbuf_1 rebuffer54 (.A(net160),
    .X(net823));
 sky130_fd_sc_hd__buf_1 rebuffer55 (.A(net49),
    .X(net824));
 sky130_fd_sc_hd__clkdlybuf4s25_2 rebuffer56 (.A(net1034),
    .X(net825));
 sky130_fd_sc_hd__clkbuf_1 rebuffer57 (.A(net127),
    .X(net826));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer6 (.A(net698),
    .X(net775));
 sky130_fd_sc_hd__clkbuf_1 rebuffer7 (.A(net1011),
    .X(net776));
 sky130_fd_sc_hd__clkbuf_1 rebuffer8 (.A(net775),
    .X(net777));
 sky130_fd_sc_hd__dlygate4sd2_1 rebuffer9 (.A(net119),
    .X(net778));
 sky130_fd_sc_hd__dfxbp_1 s818 (.CLK(clknet_2_2__leaf_clk),
    .D(net375),
    .Q(net557),
    .Q_N(net556));
 sky130_fd_sc_hd__dfxbp_1 s819 (.CLK(clknet_2_2__leaf_clk),
    .D(net401),
    .Q(net558));
 sky130_fd_sc_hd__dfxtp_2 s820 (.CLK(clknet_2_0__leaf_clk),
    .D(net463),
    .Q(net559));
 sky130_fd_sc_hd__dfxtp_2 s821 (.CLK(clknet_2_0__leaf_clk),
    .D(net467),
    .Q(net716));
 sky130_fd_sc_hd__dfxtp_1 s822 (.CLK(clknet_2_3__leaf_clk),
    .D(net484),
    .Q(net560));
 sky130_fd_sc_hd__dlclkp_1 s823 (.CLK(clknet_2_3__leaf_clk),
    .GATE(net496),
    .GCLK(net561));
 sky130_fd_sc_hd__dlclkp_2 s824 (.CLK(clknet_2_3__leaf_clk),
    .GATE(net497),
    .GCLK(net562));
 sky130_fd_sc_hd__dlclkp_4 s825 (.CLK(clknet_2_3__leaf_clk),
    .GATE(net503),
    .GCLK(net563));
 sky130_fd_sc_hd__dlxbn_1 s826 (.D(net527),
    .GATE_N(clknet_2_0__leaf_clk),
    .Q(net565),
    .Q_N(net564));
 sky130_fd_sc_hd__dlxbn_1 s827 (.D(net528),
    .GATE_N(clknet_2_0__leaf_clk),
    .Q(net567),
    .Q_N(net566));
 sky130_fd_sc_hd__buf_6 wire189 (.A(net26),
    .X(net754));
 sky130_fd_sc_hd__buf_4 wire191 (.A(net23),
    .X(net756));
 sky130_fd_sc_hd__clkbuf_1 input100 (.A(in0),
    .X(net832));
 sky130_fd_sc_hd__clkbuf_1 input101 (.A(in1),
    .X(net833));
 sky130_fd_sc_hd__buf_1 input102 (.A(in10),
    .X(net834));
 sky130_fd_sc_hd__clkbuf_1 input103 (.A(in11),
    .X(net835));
 sky130_fd_sc_hd__clkbuf_1 input104 (.A(in12),
    .X(net836));
 sky130_fd_sc_hd__clkbuf_1 input105 (.A(in13),
    .X(net837));
 sky130_fd_sc_hd__clkbuf_1 input106 (.A(in14),
    .X(net838));
 sky130_fd_sc_hd__buf_1 input107 (.A(in15),
    .X(net839));
 sky130_fd_sc_hd__buf_1 input108 (.A(in16),
    .X(net840));
 sky130_fd_sc_hd__clkbuf_1 input109 (.A(in17),
    .X(net841));
 sky130_fd_sc_hd__buf_1 input110 (.A(in18),
    .X(net842));
 sky130_fd_sc_hd__clkbuf_1 input111 (.A(in19),
    .X(net843));
 sky130_fd_sc_hd__clkbuf_1 input112 (.A(in2),
    .X(net844));
 sky130_fd_sc_hd__clkbuf_1 input113 (.A(in20),
    .X(net845));
 sky130_fd_sc_hd__clkbuf_1 input114 (.A(in21),
    .X(net846));
 sky130_fd_sc_hd__clkbuf_1 input115 (.A(in22),
    .X(net847));
 sky130_fd_sc_hd__clkbuf_1 input116 (.A(in23),
    .X(net848));
 sky130_fd_sc_hd__clkbuf_1 input117 (.A(in24),
    .X(net849));
 sky130_fd_sc_hd__clkbuf_1 input118 (.A(in25),
    .X(net850));
 sky130_fd_sc_hd__buf_1 input119 (.A(in26),
    .X(net851));
 sky130_fd_sc_hd__clkbuf_1 input120 (.A(in27),
    .X(net852));
 sky130_fd_sc_hd__clkbuf_1 input121 (.A(in28),
    .X(net853));
 sky130_fd_sc_hd__clkbuf_1 input122 (.A(in29),
    .X(net854));
 sky130_fd_sc_hd__clkbuf_1 input123 (.A(in3),
    .X(net855));
 sky130_fd_sc_hd__clkbuf_1 input124 (.A(in30),
    .X(net856));
 sky130_fd_sc_hd__clkbuf_1 input125 (.A(in31),
    .X(net857));
 sky130_fd_sc_hd__clkbuf_1 input126 (.A(in32),
    .X(net858));
 sky130_fd_sc_hd__clkbuf_1 input127 (.A(in33),
    .X(net859));
 sky130_fd_sc_hd__clkbuf_1 input128 (.A(in34),
    .X(net860));
 sky130_fd_sc_hd__clkbuf_1 input129 (.A(in35),
    .X(net861));
 sky130_fd_sc_hd__clkbuf_1 input130 (.A(in36),
    .X(net862));
 sky130_fd_sc_hd__clkbuf_1 input131 (.A(in37),
    .X(net863));
 sky130_fd_sc_hd__clkbuf_1 input132 (.A(in38),
    .X(net864));
 sky130_fd_sc_hd__clkbuf_1 input133 (.A(in39),
    .X(net865));
 sky130_fd_sc_hd__buf_6 input134 (.A(in4),
    .X(net866));
 sky130_fd_sc_hd__clkbuf_1 input135 (.A(in40),
    .X(net867));
 sky130_fd_sc_hd__clkbuf_1 input136 (.A(in41),
    .X(net868));
 sky130_fd_sc_hd__clkbuf_1 input137 (.A(in42),
    .X(net869));
 sky130_fd_sc_hd__clkbuf_1 input138 (.A(in43),
    .X(net870));
 sky130_fd_sc_hd__clkbuf_1 input139 (.A(in44),
    .X(net871));
 sky130_fd_sc_hd__clkbuf_1 input140 (.A(in45),
    .X(net872));
 sky130_fd_sc_hd__clkbuf_1 input141 (.A(in46),
    .X(net873));
 sky130_fd_sc_hd__clkbuf_1 input142 (.A(in47),
    .X(net874));
 sky130_fd_sc_hd__clkbuf_1 input143 (.A(in48),
    .X(net875));
 sky130_fd_sc_hd__clkbuf_1 input144 (.A(in49),
    .X(net876));
 sky130_fd_sc_hd__clkbuf_1 input145 (.A(in5),
    .X(net877));
 sky130_fd_sc_hd__clkbuf_1 input146 (.A(in50),
    .X(net878));
 sky130_fd_sc_hd__clkbuf_1 input147 (.A(in51),
    .X(net879));
 sky130_fd_sc_hd__clkbuf_1 input148 (.A(in52),
    .X(net880));
 sky130_fd_sc_hd__clkbuf_1 input149 (.A(in53),
    .X(net881));
 sky130_fd_sc_hd__clkbuf_1 input150 (.A(in54),
    .X(net882));
 sky130_fd_sc_hd__clkbuf_1 input151 (.A(in55),
    .X(net883));
 sky130_fd_sc_hd__clkbuf_1 input152 (.A(in56),
    .X(net884));
 sky130_fd_sc_hd__clkbuf_1 input153 (.A(in57),
    .X(net885));
 sky130_fd_sc_hd__clkbuf_1 input154 (.A(in58),
    .X(net886));
 sky130_fd_sc_hd__clkbuf_1 input155 (.A(in59),
    .X(net887));
 sky130_fd_sc_hd__clkbuf_1 input156 (.A(in6),
    .X(net888));
 sky130_fd_sc_hd__clkbuf_1 input157 (.A(in60),
    .X(net889));
 sky130_fd_sc_hd__clkbuf_1 input158 (.A(in61),
    .X(net890));
 sky130_fd_sc_hd__clkbuf_1 input159 (.A(in62),
    .X(net891));
 sky130_fd_sc_hd__clkbuf_1 input160 (.A(in63),
    .X(net892));
 sky130_fd_sc_hd__clkbuf_1 input161 (.A(in64),
    .X(net893));
 sky130_fd_sc_hd__clkbuf_1 input162 (.A(in65),
    .X(net894));
 sky130_fd_sc_hd__clkbuf_1 input163 (.A(in66),
    .X(net895));
 sky130_fd_sc_hd__clkbuf_1 input164 (.A(in67),
    .X(net896));
 sky130_fd_sc_hd__clkbuf_1 input165 (.A(in68),
    .X(net897));
 sky130_fd_sc_hd__clkbuf_1 input166 (.A(in69),
    .X(net898));
 sky130_fd_sc_hd__clkbuf_1 input167 (.A(in7),
    .X(net899));
 sky130_fd_sc_hd__clkbuf_1 input168 (.A(in70),
    .X(net900));
 sky130_fd_sc_hd__clkbuf_1 input169 (.A(in71),
    .X(net901));
 sky130_fd_sc_hd__clkbuf_1 input170 (.A(in72),
    .X(net902));
 sky130_fd_sc_hd__clkbuf_1 input171 (.A(in73),
    .X(net903));
 sky130_fd_sc_hd__buf_1 input172 (.A(in74),
    .X(net904));
 sky130_fd_sc_hd__clkbuf_1 input173 (.A(in75),
    .X(net905));
 sky130_fd_sc_hd__clkbuf_1 input174 (.A(in76),
    .X(net906));
 sky130_fd_sc_hd__clkbuf_1 input175 (.A(in77),
    .X(net907));
 sky130_fd_sc_hd__clkbuf_1 input176 (.A(in78),
    .X(net908));
 sky130_fd_sc_hd__clkbuf_1 input177 (.A(in79),
    .X(net909));
 sky130_fd_sc_hd__clkbuf_1 input178 (.A(in8),
    .X(net910));
 sky130_fd_sc_hd__clkbuf_1 input179 (.A(in80),
    .X(net911));
 sky130_fd_sc_hd__clkbuf_1 input180 (.A(in81),
    .X(net912));
 sky130_fd_sc_hd__clkbuf_1 input181 (.A(in82),
    .X(net913));
 sky130_fd_sc_hd__clkbuf_1 input182 (.A(in83),
    .X(net914));
 sky130_fd_sc_hd__clkbuf_1 input183 (.A(in84),
    .X(net915));
 sky130_fd_sc_hd__clkbuf_1 input184 (.A(in85),
    .X(net916));
 sky130_fd_sc_hd__clkbuf_1 input185 (.A(in86),
    .X(net917));
 sky130_fd_sc_hd__clkbuf_1 input186 (.A(in87),
    .X(net918));
 sky130_fd_sc_hd__clkbuf_1 input187 (.A(in88),
    .X(net919));
 sky130_fd_sc_hd__clkbuf_1 input188 (.A(in89),
    .X(net920));
 sky130_fd_sc_hd__clkbuf_1 input189 (.A(in9),
    .X(net921));
 sky130_fd_sc_hd__clkbuf_1 input190 (.A(in90),
    .X(net922));
 sky130_fd_sc_hd__clkbuf_1 input191 (.A(in91),
    .X(net923));
 sky130_fd_sc_hd__clkbuf_1 input192 (.A(in92),
    .X(net924));
 sky130_fd_sc_hd__clkbuf_1 input193 (.A(in93),
    .X(net925));
 sky130_fd_sc_hd__clkbuf_1 input194 (.A(in94),
    .X(net926));
 sky130_fd_sc_hd__buf_1 input195 (.A(in95),
    .X(net927));
 sky130_fd_sc_hd__clkbuf_1 input196 (.A(in97),
    .X(net928));
 sky130_fd_sc_hd__clkbuf_1 input197 (.A(in98),
    .X(net929));
 sky130_fd_sc_hd__clkbuf_1 input198 (.A(in99),
    .X(net930));
 sky130_fd_sc_hd__clkbuf_4 output199 (.A(net931),
    .X(out0));
 sky130_fd_sc_hd__clkbuf_4 output200 (.A(net932),
    .X(out1));
 sky130_fd_sc_hd__buf_2 output201 (.A(net933),
    .X(out10));
 sky130_fd_sc_hd__buf_2 output202 (.A(net934),
    .X(out11));
 sky130_fd_sc_hd__buf_2 output203 (.A(net935),
    .X(out13));
 sky130_fd_sc_hd__buf_2 output204 (.A(net936),
    .X(out15));
 sky130_fd_sc_hd__clkbuf_4 output205 (.A(net937),
    .X(out16));
 sky130_fd_sc_hd__buf_2 output206 (.A(net938),
    .X(out17));
 sky130_fd_sc_hd__buf_2 output207 (.A(net939),
    .X(out18));
 sky130_fd_sc_hd__clkbuf_4 output208 (.A(net940),
    .X(out19));
 sky130_fd_sc_hd__buf_2 output209 (.A(net941),
    .X(out2));
 sky130_fd_sc_hd__buf_2 output210 (.A(net942),
    .X(out20));
 sky130_fd_sc_hd__clkbuf_4 output211 (.A(net943),
    .X(out21));
 sky130_fd_sc_hd__buf_2 output212 (.A(net944),
    .X(out22));
 sky130_fd_sc_hd__buf_2 output213 (.A(net945),
    .X(out26));
 sky130_fd_sc_hd__buf_2 output214 (.A(net946),
    .X(out28));
 sky130_fd_sc_hd__buf_2 output215 (.A(net947),
    .X(out3));
 sky130_fd_sc_hd__clkbuf_4 output216 (.A(net948),
    .X(out30));
 sky130_fd_sc_hd__clkbuf_4 output217 (.A(net949),
    .X(out32));
 sky130_fd_sc_hd__buf_2 output218 (.A(net950),
    .X(out33));
 sky130_fd_sc_hd__buf_2 output219 (.A(net951),
    .X(out34));
 sky130_fd_sc_hd__buf_2 output220 (.A(net952),
    .X(out35));
 sky130_fd_sc_hd__buf_2 output221 (.A(net953),
    .X(out36));
 sky130_fd_sc_hd__buf_2 output222 (.A(net954),
    .X(out38));
 sky130_fd_sc_hd__buf_2 output223 (.A(net955),
    .X(out39));
 sky130_fd_sc_hd__clkbuf_4 output224 (.A(net956),
    .X(out4));
 sky130_fd_sc_hd__buf_2 output225 (.A(net957),
    .X(out40));
 sky130_fd_sc_hd__buf_2 output226 (.A(net958),
    .X(out42));
 sky130_fd_sc_hd__buf_2 output227 (.A(net959),
    .X(out45));
 sky130_fd_sc_hd__buf_2 output228 (.A(net960),
    .X(out46));
 sky130_fd_sc_hd__buf_2 output229 (.A(net961),
    .X(out47));
 sky130_fd_sc_hd__buf_2 output230 (.A(net962),
    .X(out49));
 sky130_fd_sc_hd__buf_2 output231 (.A(net963),
    .X(out5));
 sky130_fd_sc_hd__buf_2 output232 (.A(net964),
    .X(out50));
 sky130_fd_sc_hd__buf_2 output233 (.A(net965),
    .X(out51));
 sky130_fd_sc_hd__buf_2 output234 (.A(net966),
    .X(out52));
 sky130_fd_sc_hd__buf_2 output235 (.A(net967),
    .X(out53));
 sky130_fd_sc_hd__buf_2 output236 (.A(net968),
    .X(out54));
 sky130_fd_sc_hd__buf_2 output237 (.A(net969),
    .X(out55));
 sky130_fd_sc_hd__buf_2 output238 (.A(net970),
    .X(out57));
 sky130_fd_sc_hd__buf_2 output239 (.A(net971),
    .X(out58));
 sky130_fd_sc_hd__buf_2 output240 (.A(net972),
    .X(out59));
 sky130_fd_sc_hd__buf_2 output241 (.A(net973),
    .X(out6));
 sky130_fd_sc_hd__buf_2 output242 (.A(net974),
    .X(out60));
 sky130_fd_sc_hd__buf_2 output243 (.A(net975),
    .X(out61));
 sky130_fd_sc_hd__buf_2 output244 (.A(net976),
    .X(out62));
 sky130_fd_sc_hd__buf_2 output245 (.A(net977),
    .X(out63));
 sky130_fd_sc_hd__buf_2 output246 (.A(net978),
    .X(out65));
 sky130_fd_sc_hd__buf_2 output247 (.A(net979),
    .X(out67));
 sky130_fd_sc_hd__buf_2 output248 (.A(net980),
    .X(out68));
 sky130_fd_sc_hd__buf_2 output249 (.A(net981),
    .X(out69));
 sky130_fd_sc_hd__clkbuf_4 output250 (.A(net982),
    .X(out7));
 sky130_fd_sc_hd__buf_2 output251 (.A(net983),
    .X(out71));
 sky130_fd_sc_hd__buf_2 output252 (.A(net984),
    .X(out72));
 sky130_fd_sc_hd__buf_2 output253 (.A(net985),
    .X(out73));
 sky130_fd_sc_hd__buf_2 output254 (.A(net986),
    .X(out75));
 sky130_fd_sc_hd__buf_2 output255 (.A(net987),
    .X(out76));
 sky130_fd_sc_hd__buf_2 output256 (.A(net988),
    .X(out79));
 sky130_fd_sc_hd__buf_2 output257 (.A(net989),
    .X(out8));
 sky130_fd_sc_hd__buf_2 output258 (.A(net990),
    .X(out81));
 sky130_fd_sc_hd__buf_2 output259 (.A(net991),
    .X(out82));
 sky130_fd_sc_hd__buf_2 output260 (.A(net992),
    .X(out83));
 sky130_fd_sc_hd__buf_2 output261 (.A(net993),
    .X(out84));
 sky130_fd_sc_hd__buf_2 output262 (.A(net994),
    .X(out85));
 sky130_fd_sc_hd__buf_2 output263 (.A(net995),
    .X(out86));
 sky130_fd_sc_hd__buf_2 output264 (.A(net996),
    .X(out88));
 sky130_fd_sc_hd__buf_2 output265 (.A(net997),
    .X(out89));
 sky130_fd_sc_hd__buf_2 output266 (.A(net998),
    .X(out9));
 sky130_fd_sc_hd__buf_2 output267 (.A(net999),
    .X(out91));
 sky130_fd_sc_hd__buf_2 output268 (.A(net1000),
    .X(out92));
 sky130_fd_sc_hd__buf_2 output269 (.A(net1001),
    .X(out93));
 sky130_fd_sc_hd__buf_2 output270 (.A(net1002),
    .X(out94));
 sky130_fd_sc_hd__buf_2 output271 (.A(net1003),
    .X(out95));
 sky130_fd_sc_hd__buf_2 output272 (.A(net1004),
    .X(out96));
 sky130_fd_sc_hd__buf_2 output273 (.A(net1005),
    .X(out98));
 sky130_fd_sc_hd__buf_6 fanout274 (.A(net349),
    .X(net1006));
 sky130_fd_sc_hd__buf_6 fanout275 (.A(net540),
    .X(net1007));
 sky130_fd_sc_hd__clkbuf_2 fanout276 (.A(net255),
    .X(net1008));
 sky130_fd_sc_hd__buf_6 fanout277 (.A(net255),
    .X(net1009));
 sky130_fd_sc_hd__clkbuf_2 fanout278 (.A(net355),
    .X(net1010));
 sky130_fd_sc_hd__clkbuf_4 fanout279 (.A(net775),
    .X(net1011));
 sky130_fd_sc_hd__clkbuf_4 fanout280 (.A(net307),
    .X(net1012));
 sky130_fd_sc_hd__buf_2 fanout281 (.A(net188),
    .X(net1013));
 sky130_fd_sc_hd__buf_1 fanout282 (.A(net1015),
    .X(net1014));
 sky130_fd_sc_hd__clkbuf_2 fanout283 (.A(net1016),
    .X(net1015));
 sky130_fd_sc_hd__buf_2 fanout284 (.A(net740),
    .X(net1016));
 sky130_fd_sc_hd__buf_2 fanout285 (.A(net305),
    .X(net1017));
 sky130_fd_sc_hd__buf_1 fanout286 (.A(net1019),
    .X(net1018));
 sky130_fd_sc_hd__buf_4 fanout287 (.A(net151),
    .X(net1019));
 sky130_fd_sc_hd__clkbuf_4 fanout288 (.A(net723),
    .X(net1020));
 sky130_fd_sc_hd__clkbuf_2 fanout289 (.A(net744),
    .X(net1021));
 sky130_fd_sc_hd__buf_1 fanout290 (.A(net1023),
    .X(net1022));
 sky130_fd_sc_hd__clkbuf_2 fanout291 (.A(net1024),
    .X(net1023));
 sky130_fd_sc_hd__clkbuf_2 fanout292 (.A(net743),
    .X(net1024));
 sky130_fd_sc_hd__buf_1 fanout293 (.A(net1026),
    .X(net1025));
 sky130_fd_sc_hd__buf_4 fanout294 (.A(net741),
    .X(net1026));
 sky130_fd_sc_hd__buf_2 fanout295 (.A(net227),
    .X(net1027));
 sky130_fd_sc_hd__clkbuf_4 fanout296 (.A(net226),
    .X(net1028));
 sky130_fd_sc_hd__clkbuf_2 fanout297 (.A(net1030),
    .X(net1029));
 sky130_fd_sc_hd__buf_6 fanout298 (.A(net139),
    .X(net1030));
 sky130_fd_sc_hd__clkbuf_2 fanout299 (.A(net745),
    .X(net1031));
 sky130_fd_sc_hd__buf_4 max_cap300 (.A(net296),
    .X(net1032));
 sky130_fd_sc_hd__buf_2 fanout301 (.A(net774),
    .X(net1033));
 sky130_fd_sc_hd__buf_1 fanout302 (.A(net1035),
    .X(net1034));
 sky130_fd_sc_hd__buf_8 fanout303 (.A(net746),
    .X(net1035));
 sky130_fd_sc_hd__buf_4 fanout304 (.A(net147),
    .X(net1036));
 sky130_fd_sc_hd__buf_6 fanout305 (.A(net61),
    .X(net1037));
 sky130_fd_sc_hd__buf_8 fanout306 (.A(net747),
    .X(net1038));
 sky130_fd_sc_hd__clkbuf_2 fanout307 (.A(net364),
    .X(net1039));
 sky130_fd_sc_hd__clkbuf_2 fanout308 (.A(net364),
    .X(net1040));
 sky130_fd_sc_hd__buf_2 fanout309 (.A(net129),
    .X(net1041));
 sky130_fd_sc_hd__clkbuf_4 fanout310 (.A(net116),
    .X(net1042));
 sky130_fd_sc_hd__buf_4 max_cap311 (.A(net113),
    .X(net1043));
 sky130_fd_sc_hd__buf_2 fanout312 (.A(net1045),
    .X(net1044));
 sky130_fd_sc_hd__buf_4 fanout313 (.A(net112),
    .X(net1045));
 sky130_fd_sc_hd__clkbuf_2 fanout314 (.A(net1047),
    .X(net1046));
 sky130_fd_sc_hd__buf_6 fanout315 (.A(net110),
    .X(net1047));
 sky130_fd_sc_hd__clkbuf_4 fanout316 (.A(net711),
    .X(net1048));
 sky130_fd_sc_hd__clkbuf_4 fanout317 (.A(net682),
    .X(net1049));
 sky130_fd_sc_hd__clkbuf_2 fanout318 (.A(net126),
    .X(net1050));
 sky130_fd_sc_hd__buf_6 max_cap319 (.A(net107),
    .X(net1051));
 sky130_fd_sc_hd__buf_4 fanout320 (.A(net45),
    .X(net1052));
 sky130_fd_sc_hd__clkbuf_4 fanout321 (.A(net28),
    .X(net1053));
 sky130_fd_sc_hd__clkbuf_4 fanout322 (.A(net685),
    .X(net1054));
 sky130_fd_sc_hd__buf_2 fanout323 (.A(net757),
    .X(net1055));
 sky130_fd_sc_hd__buf_2 fanout324 (.A(net57),
    .X(net1056));
 sky130_fd_sc_hd__buf_4 fanout325 (.A(net29),
    .X(net1057));
 sky130_fd_sc_hd__buf_2 fanout326 (.A(net681),
    .X(net1058));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout327 (.A(net1060),
    .X(net1059));
 sky130_fd_sc_hd__clkbuf_2 fanout328 (.A(net1061),
    .X(net1060));
 sky130_fd_sc_hd__clkbuf_4 fanout329 (.A(net44),
    .X(net1061));
 sky130_fd_sc_hd__buf_2 fanout330 (.A(net42),
    .X(net1062));
 sky130_fd_sc_hd__clkbuf_2 fanout331 (.A(net1064),
    .X(net1063));
 sky130_fd_sc_hd__buf_4 fanout332 (.A(net20),
    .X(net1064));
 sky130_fd_sc_hd__buf_2 fanout333 (.A(net36),
    .X(net1065));
 sky130_fd_sc_hd__buf_6 fanout334 (.A(net732),
    .X(net1066));
 sky130_fd_sc_hd__buf_4 fanout335 (.A(net18),
    .X(net1067));
 sky130_fd_sc_hd__clkbuf_4 fanout336 (.A(net108),
    .X(net1068));
 sky130_fd_sc_hd__buf_2 fanout337 (.A(net40),
    .X(net1069));
 sky130_fd_sc_hd__clkbuf_2 fanout338 (.A(net40),
    .X(net1070));
 sky130_fd_sc_hd__buf_4 fanout339 (.A(net697),
    .X(net1071));
 sky130_fd_sc_hd__clkbuf_4 fanout340 (.A(net60),
    .X(net1072));
 sky130_fd_sc_hd__clkbuf_4 fanout341 (.A(net53),
    .X(net1073));
 sky130_fd_sc_hd__clkbuf_2 fanout342 (.A(net34),
    .X(net1074));
 sky130_fd_sc_hd__clkbuf_2 fanout343 (.A(net34),
    .X(net1075));
 sky130_fd_sc_hd__buf_2 fanout344 (.A(net19),
    .X(net1076));
 sky130_fd_sc_hd__buf_2 fanout345 (.A(net19),
    .X(net1077));
 sky130_fd_sc_hd__buf_2 fanout346 (.A(net17),
    .X(net1078));
 sky130_fd_sc_hd__clkbuf_2 fanout347 (.A(net17),
    .X(net1079));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout348 (.A(net1081),
    .X(net1080));
 sky130_fd_sc_hd__clkbuf_2 fanout349 (.A(net559),
    .X(net1081));
 sky130_fd_sc_hd__clkbuf_2 fanout350 (.A(net714),
    .X(net1082));
 sky130_fd_sc_hd__buf_2 fanout351 (.A(net767),
    .X(net1083));
 sky130_fd_sc_hd__buf_1 fanout352 (.A(net1085),
    .X(net1084));
 sky130_fd_sc_hd__clkbuf_4 fanout353 (.A(net1086),
    .X(net1085));
 sky130_fd_sc_hd__clkbuf_4 fanout354 (.A(net768),
    .X(net1086));
 sky130_fd_sc_hd__buf_2 fanout355 (.A(net726),
    .X(net1087));
 sky130_fd_sc_hd__buf_2 fanout356 (.A(net713),
    .X(net1088));
 sky130_fd_sc_hd__clkbuf_2 fanout357 (.A(net1090),
    .X(net1089));
 sky130_fd_sc_hd__buf_2 fanout358 (.A(net769),
    .X(net1090));
 sky130_fd_sc_hd__buf_2 fanout359 (.A(net104),
    .X(net1091));
 sky130_fd_sc_hd__clkbuf_2 fanout360 (.A(net30),
    .X(net1092));
 sky130_fd_sc_hd__clkbuf_4 fanout361 (.A(net15),
    .X(net1093));
 sky130_fd_sc_hd__clkbuf_4 fanout362 (.A(net660),
    .X(net1094));
 sky130_fd_sc_hd__buf_4 fanout363 (.A(net655),
    .X(net1095));
 sky130_fd_sc_hd__buf_4 fanout364 (.A(net574),
    .X(net1096));
 sky130_fd_sc_hd__clkbuf_8 fanout365 (.A(net573),
    .X(net1097));
 sky130_fd_sc_hd__buf_4 fanout366 (.A(net644),
    .X(net1098));
 sky130_fd_sc_hd__clkbuf_4 fanout367 (.A(net572),
    .X(net1099));
 sky130_fd_sc_hd__buf_4 fanout368 (.A(net571),
    .X(net1100));
 sky130_fd_sc_hd__buf_4 fanout369 (.A(net1102),
    .X(net1101));
 sky130_fd_sc_hd__buf_2 fanout370 (.A(net622),
    .X(net1102));
 sky130_fd_sc_hd__buf_2 fanout371 (.A(net1104),
    .X(net1103));
 sky130_fd_sc_hd__clkbuf_4 fanout372 (.A(net617),
    .X(net1104));
 sky130_fd_sc_hd__clkbuf_2 fanout373 (.A(net1106),
    .X(net1105));
 sky130_fd_sc_hd__clkbuf_4 fanout374 (.A(net612),
    .X(net1106));
 sky130_fd_sc_hd__clkbuf_4 fanout375 (.A(net611),
    .X(net1107));
 sky130_fd_sc_hd__buf_2 fanout376 (.A(net1109),
    .X(net1108));
 sky130_fd_sc_hd__clkbuf_4 fanout377 (.A(net569),
    .X(net1109));
 sky130_fd_sc_hd__buf_12 fanout378 (.A(net600),
    .X(net1110));
 sky130_fd_sc_hd__buf_4 fanout379 (.A(net598),
    .X(net1111));
 sky130_fd_sc_hd__buf_2 fanout380 (.A(net596),
    .X(net1112));
 sky130_fd_sc_hd__buf_12 fanout381 (.A(net568),
    .X(net1113));
 sky130_fd_sc_hd__clkbuf_2 fanout382 (.A(net1115),
    .X(net1114));
 sky130_fd_sc_hd__clkbuf_8 fanout383 (.A(net592),
    .X(net1115));
 sky130_fd_sc_hd__buf_4 fanout384 (.A(net589),
    .X(net1116));
 sky130_fd_sc_hd__buf_1 fanout385 (.A(net1118),
    .X(net1117));
 sky130_fd_sc_hd__buf_8 fanout386 (.A(net585),
    .X(net1118));
 sky130_fd_sc_hd__buf_2 fanout387 (.A(net1120),
    .X(net1119));
 sky130_fd_sc_hd__buf_4 fanout388 (.A(net550),
    .X(net1120));
 sky130_fd_sc_hd__buf_4 fanout389 (.A(net580),
    .X(net1121));
 sky130_fd_sc_hd__clkbuf_4 fanout390 (.A(net578),
    .X(net1122));
 sky130_fd_sc_hd__buf_4 fanout391 (.A(net576),
    .X(net1123));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer5 (.A(net16),
    .X(net1124));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer22 (.A(net1157),
    .X(net1125));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer58 (.A(net351),
    .X(net1126));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer59 (.A(net204),
    .X(net1127));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer60 (.A(net1007),
    .X(net1128));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer61 (.A(net1130),
    .X(net1129));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer62 (.A(net56),
    .X(net1130));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer63 (.A(net682),
    .X(net1131));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer64 (.A(net1131),
    .X(net1132));
 sky130_fd_sc_hd__clkbuf_1 rebuffer65 (.A(net201),
    .X(net1133));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer66 (.A(net1133),
    .X(net1134));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer67 (.A(net1136),
    .X(net1135));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer68 (.A(net1137),
    .X(net1136));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer69 (.A(net1138),
    .X(net1137));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer70 (.A(net1139),
    .X(net1138));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer71 (.A(net1140),
    .X(net1139));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer72 (.A(net247),
    .X(net1140));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer73 (.A(net540),
    .X(net1141));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer74 (.A(net249),
    .X(net1142));
 sky130_fd_sc_hd__clkbuf_1 clone75 (.A(net600),
    .X(net1143));
 sky130_fd_sc_hd__clkbuf_1 clone76 (.A(net747),
    .X(net1144));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer77 (.A(net204),
    .X(net1145));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer78 (.A(net1145),
    .X(net1146));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer79 (.A(net224),
    .X(net1147));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer80 (.A(net1147),
    .X(net1148));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer81 (.A(net172),
    .X(net1149));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer82 (.A(net234),
    .X(net1150));
 sky130_fd_sc_hd__clkbuf_1 clone83 (.A(net568),
    .X(net1151));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer84 (.A(net1035),
    .X(net1152));
 sky130_fd_sc_hd__clkbuf_1 clone85 (.A(net349),
    .X(net1153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(net559),
    .X(net1154));
 sky130_fd_sc_hd__diode_2 ANTENNA_input100_A (.DIODE(in0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input101_A (.DIODE(in1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input102_A (.DIODE(in10));
 sky130_fd_sc_hd__diode_2 ANTENNA_input103_A (.DIODE(in11));
 sky130_fd_sc_hd__diode_2 ANTENNA_input104_A (.DIODE(in12));
 sky130_fd_sc_hd__diode_2 ANTENNA_input105_A (.DIODE(in13));
 sky130_fd_sc_hd__diode_2 ANTENNA_input106_A (.DIODE(in14));
 sky130_fd_sc_hd__diode_2 ANTENNA_input107_A (.DIODE(in15));
 sky130_fd_sc_hd__diode_2 ANTENNA_input108_A (.DIODE(in16));
 sky130_fd_sc_hd__diode_2 ANTENNA_input109_A (.DIODE(in17));
 sky130_fd_sc_hd__diode_2 ANTENNA_input110_A (.DIODE(in18));
 sky130_fd_sc_hd__diode_2 ANTENNA_input111_A (.DIODE(in19));
 sky130_fd_sc_hd__diode_2 ANTENNA_input112_A (.DIODE(in2));
 sky130_fd_sc_hd__diode_2 ANTENNA_input113_A (.DIODE(in20));
 sky130_fd_sc_hd__diode_2 ANTENNA_input114_A (.DIODE(in21));
 sky130_fd_sc_hd__diode_2 ANTENNA_input115_A (.DIODE(in22));
 sky130_fd_sc_hd__diode_2 ANTENNA_input116_A (.DIODE(in23));
 sky130_fd_sc_hd__diode_2 ANTENNA_input117_A (.DIODE(in24));
 sky130_fd_sc_hd__diode_2 ANTENNA_input118_A (.DIODE(in25));
 sky130_fd_sc_hd__diode_2 ANTENNA_input119_A (.DIODE(in26));
 sky130_fd_sc_hd__diode_2 ANTENNA_input120_A (.DIODE(in27));
 sky130_fd_sc_hd__diode_2 ANTENNA_input121_A (.DIODE(in28));
 sky130_fd_sc_hd__diode_2 ANTENNA_input122_A (.DIODE(in29));
 sky130_fd_sc_hd__diode_2 ANTENNA_input123_A (.DIODE(in3));
 sky130_fd_sc_hd__diode_2 ANTENNA_input124_A (.DIODE(in30));
 sky130_fd_sc_hd__diode_2 ANTENNA_input125_A (.DIODE(in31));
 sky130_fd_sc_hd__diode_2 ANTENNA_input126_A (.DIODE(in32));
 sky130_fd_sc_hd__diode_2 ANTENNA_input127_A (.DIODE(in33));
 sky130_fd_sc_hd__diode_2 ANTENNA_input128_A (.DIODE(in34));
 sky130_fd_sc_hd__diode_2 ANTENNA_input129_A (.DIODE(in35));
 sky130_fd_sc_hd__diode_2 ANTENNA_input130_A (.DIODE(in36));
 sky130_fd_sc_hd__diode_2 ANTENNA_input131_A (.DIODE(in37));
 sky130_fd_sc_hd__diode_2 ANTENNA_input132_A (.DIODE(in38));
 sky130_fd_sc_hd__diode_2 ANTENNA_input133_A (.DIODE(in39));
 sky130_fd_sc_hd__diode_2 ANTENNA_input134_A (.DIODE(in4));
 sky130_fd_sc_hd__diode_2 ANTENNA_input135_A (.DIODE(in40));
 sky130_fd_sc_hd__diode_2 ANTENNA_input136_A (.DIODE(in41));
 sky130_fd_sc_hd__diode_2 ANTENNA_input137_A (.DIODE(in42));
 sky130_fd_sc_hd__diode_2 ANTENNA_input138_A (.DIODE(in43));
 sky130_fd_sc_hd__diode_2 ANTENNA_input139_A (.DIODE(in44));
 sky130_fd_sc_hd__diode_2 ANTENNA_input140_A (.DIODE(in45));
 sky130_fd_sc_hd__diode_2 ANTENNA_input141_A (.DIODE(in46));
 sky130_fd_sc_hd__diode_2 ANTENNA_input142_A (.DIODE(in47));
 sky130_fd_sc_hd__diode_2 ANTENNA_input143_A (.DIODE(in48));
 sky130_fd_sc_hd__diode_2 ANTENNA_input144_A (.DIODE(in49));
 sky130_fd_sc_hd__diode_2 ANTENNA_input145_A (.DIODE(in5));
 sky130_fd_sc_hd__diode_2 ANTENNA_input146_A (.DIODE(in50));
 sky130_fd_sc_hd__diode_2 ANTENNA_input147_A (.DIODE(in51));
 sky130_fd_sc_hd__diode_2 ANTENNA_input148_A (.DIODE(in52));
 sky130_fd_sc_hd__diode_2 ANTENNA_input149_A (.DIODE(in53));
 sky130_fd_sc_hd__diode_2 ANTENNA_input150_A (.DIODE(in54));
 sky130_fd_sc_hd__diode_2 ANTENNA_input151_A (.DIODE(in55));
 sky130_fd_sc_hd__diode_2 ANTENNA_input152_A (.DIODE(in56));
 sky130_fd_sc_hd__diode_2 ANTENNA_input153_A (.DIODE(in57));
 sky130_fd_sc_hd__diode_2 ANTENNA_input154_A (.DIODE(in58));
 sky130_fd_sc_hd__diode_2 ANTENNA_input155_A (.DIODE(in59));
 sky130_fd_sc_hd__diode_2 ANTENNA_input156_A (.DIODE(in6));
 sky130_fd_sc_hd__diode_2 ANTENNA_input157_A (.DIODE(in60));
 sky130_fd_sc_hd__diode_2 ANTENNA_input158_A (.DIODE(in61));
 sky130_fd_sc_hd__diode_2 ANTENNA_input159_A (.DIODE(in62));
 sky130_fd_sc_hd__diode_2 ANTENNA_input160_A (.DIODE(in63));
 sky130_fd_sc_hd__diode_2 ANTENNA_input161_A (.DIODE(in64));
 sky130_fd_sc_hd__diode_2 ANTENNA_input162_A (.DIODE(in65));
 sky130_fd_sc_hd__diode_2 ANTENNA_input163_A (.DIODE(in66));
 sky130_fd_sc_hd__diode_2 ANTENNA_input164_A (.DIODE(in67));
 sky130_fd_sc_hd__diode_2 ANTENNA_input165_A (.DIODE(in68));
 sky130_fd_sc_hd__diode_2 ANTENNA_input166_A (.DIODE(in69));
 sky130_fd_sc_hd__diode_2 ANTENNA_input167_A (.DIODE(in7));
 sky130_fd_sc_hd__diode_2 ANTENNA_input168_A (.DIODE(in70));
 sky130_fd_sc_hd__diode_2 ANTENNA_input169_A (.DIODE(in71));
 sky130_fd_sc_hd__diode_2 ANTENNA_input170_A (.DIODE(in72));
 sky130_fd_sc_hd__diode_2 ANTENNA_input171_A (.DIODE(in73));
 sky130_fd_sc_hd__diode_2 ANTENNA_input172_A (.DIODE(in74));
 sky130_fd_sc_hd__diode_2 ANTENNA_input173_A (.DIODE(in75));
 sky130_fd_sc_hd__diode_2 ANTENNA_input174_A (.DIODE(in76));
 sky130_fd_sc_hd__diode_2 ANTENNA_input175_A (.DIODE(in77));
 sky130_fd_sc_hd__diode_2 ANTENNA_input176_A (.DIODE(in78));
 sky130_fd_sc_hd__diode_2 ANTENNA_input177_A (.DIODE(in79));
 sky130_fd_sc_hd__diode_2 ANTENNA_input178_A (.DIODE(in8));
 sky130_fd_sc_hd__diode_2 ANTENNA_input179_A (.DIODE(in80));
 sky130_fd_sc_hd__diode_2 ANTENNA_input180_A (.DIODE(in81));
 sky130_fd_sc_hd__diode_2 ANTENNA_input181_A (.DIODE(in82));
 sky130_fd_sc_hd__diode_2 ANTENNA_input182_A (.DIODE(in83));
 sky130_fd_sc_hd__diode_2 ANTENNA_input183_A (.DIODE(in84));
 sky130_fd_sc_hd__diode_2 ANTENNA_input184_A (.DIODE(in85));
 sky130_fd_sc_hd__diode_2 ANTENNA_input185_A (.DIODE(in86));
 sky130_fd_sc_hd__diode_2 ANTENNA_input186_A (.DIODE(in87));
 sky130_fd_sc_hd__diode_2 ANTENNA_input187_A (.DIODE(in88));
 sky130_fd_sc_hd__diode_2 ANTENNA_input188_A (.DIODE(in89));
 sky130_fd_sc_hd__diode_2 ANTENNA_input189_A (.DIODE(in9));
 sky130_fd_sc_hd__diode_2 ANTENNA_input190_A (.DIODE(in90));
 sky130_fd_sc_hd__diode_2 ANTENNA_input191_A (.DIODE(in91));
 sky130_fd_sc_hd__diode_2 ANTENNA_input192_A (.DIODE(in92));
 sky130_fd_sc_hd__diode_2 ANTENNA_input193_A (.DIODE(in93));
 sky130_fd_sc_hd__diode_2 ANTENNA_input194_A (.DIODE(in94));
 sky130_fd_sc_hd__diode_2 ANTENNA_input195_A (.DIODE(in95));
 sky130_fd_sc_hd__diode_2 ANTENNA_input196_A (.DIODE(in97));
 sky130_fd_sc_hd__diode_2 ANTENNA_input197_A (.DIODE(in98));
 sky130_fd_sc_hd__diode_2 ANTENNA_input198_A (.DIODE(in99));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_A1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_A2 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c446_A2 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c277_A (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_Y (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout359_A (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_A3_1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_A2_1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_B1_N_1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c272_Y_1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout336_A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_A2_1 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA_c276_Y_1 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap311_A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c416_B_1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_Y_1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout310_A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_A2_1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_X_1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout318_A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_A0_1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_c295_Y_1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout309_A (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_A2_1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_Y_1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap201_A (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_A2 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c159_A (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_Y (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_A1 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_A2 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_Y (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout361_A (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_A1_1 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_A2_1 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_c398_B1_N_1 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_Y_1 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_A0 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_A3 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_X (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout347_A (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout346_A (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_Y_1 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout345_A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout344_A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_Y_1 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_A1 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_c678_B1 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_B (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_A2 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_c406_X (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_A1 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_c531_B (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_X (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_B1_N (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_A (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_B (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA_c428_B (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_X (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_A2 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA_c611_A2 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_A1 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_A3 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_B (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_Y (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_A1 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_B1_N (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_Y (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout321_A (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c764_A0_1 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_X_1 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout325_A (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_c239_A0_1 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_A1_1 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_A4_1 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_X_1 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_A1 (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA_c563_B (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA_c541_A2 (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA_c535_A (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA_c534_B (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA_c530_Y (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_A (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout360_A (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_A3_1 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_A2_1 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_Y_1 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_A (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA_c678_A3 (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA_c562_B (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA_c535_B (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA_c533_B (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA_c532_Y (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout285_A (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA_c545_B_1 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA_c537_Y_1 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA_c701_A2 (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_A2 (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_A2 (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA_c558_A1 (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA_c554_B1 (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_B1_N (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_Y (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_A1 (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA_c564_Y (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout343_A (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout342_A (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_Y_1 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout333_A (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c763_S0_1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_Y_1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout308_A (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout307_A (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_Y_1 (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout338_A (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout337_A (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_X_1 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout330_A (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_A1_1 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_X_1 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_c286_B_1 (.DIODE(net1158));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout320_A (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_A2_1 (.DIODE(net1158));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_B1_N_1 (.DIODE(net1158));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_X_1 (.DIODE(net1158));
 sky130_fd_sc_hd__diode_2 ANTENNA_c428_A (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_A2 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_B (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_B1_N (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_X (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_A2 (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA_c720_B1_N (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_A0 (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_X (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_A1 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_c183_A (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_c180_X (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold86_A (.DIODE(net559));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout349_A (.DIODE(net559));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_B1_1 (.DIODE(net559));
 sky130_fd_sc_hd__diode_2 ANTENNA_c767_S1_1 (.DIODE(net559));
 sky130_fd_sc_hd__diode_2 ANTENNA_s820_Q_1 (.DIODE(net559));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone83_A (.DIODE(net568));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout381_A (.DIODE(net568));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_S0_1 (.DIODE(net568));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_X_1 (.DIODE(net568));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_A2 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout324_A (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_A3_1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_B1_N_1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_X_1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout368_A (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA_c116_A_1 (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_X_1 (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout364_A (.DIODE(net574));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_X_1 (.DIODE(net574));
 sky130_fd_sc_hd__diode_2 ANTENNA_c765_S1_1 (.DIODE(net574));
 sky130_fd_sc_hd__diode_2 ANTENNA_c743_A4_1 (.DIODE(net574));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_S0_1 (.DIODE(net574));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout391_A (.DIODE(net576));
 sky130_fd_sc_hd__diode_2 ANTENNA_c235_B_1 (.DIODE(net576));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_X_1 (.DIODE(net576));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_A1 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_B (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_A4 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA_c203_B (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_Y (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout389_A (.DIODE(net580));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_A3_1 (.DIODE(net580));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_B_1 (.DIODE(net580));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_A3_1 (.DIODE(net580));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_X_1 (.DIODE(net580));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout384_A (.DIODE(net589));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge791_S1_1 (.DIODE(net589));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_X_1 (.DIODE(net589));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer14_A (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer13_A (.DIODE(net1155));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_B (.DIODE(net1155));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_A2 (.DIODE(net1155));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_B1 (.DIODE(net1155));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_A1 (.DIODE(net1155));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_S0 (.DIODE(net1155));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_X (.DIODE(net1155));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout340_A (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA_c765_A2_1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_S0_1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_A2_1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA_c190_X_1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout305_A (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA_c373_A3_1 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA_c191_Y_1 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout375_A (.DIODE(net611));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_A1_1 (.DIODE(net611));
 sky130_fd_sc_hd__diode_2 ANTENNA_input46_X_1 (.DIODE(net611));
 sky130_fd_sc_hd__diode_2 ANTENNA_c744_A1_1 (.DIODE(net611));
 sky130_fd_sc_hd__diode_2 ANTENNA_c610_A2_1 (.DIODE(net611));
 sky130_fd_sc_hd__diode_2 ANTENNA_input65_X (.DIODE(net630));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_A (.DIODE(net630));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout363_A (.DIODE(net655));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_A2_1 (.DIODE(net655));
 sky130_fd_sc_hd__diode_2 ANTENNA_input90_X_1 (.DIODE(net655));
 sky130_fd_sc_hd__diode_2 ANTENNA_output100_A (.DIODE(net665));
 sky130_fd_sc_hd__diode_2 ANTENNA_c743_X (.DIODE(net665));
 sky130_fd_sc_hd__diode_2 ANTENNA_output119_A (.DIODE(net684));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_X (.DIODE(net684));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout322_A (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA_c232_B1_N_1 (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA_c611_A1_1 (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA_c762_A1_1 (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_X_1 (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA_output122_A (.DIODE(net687));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_B1_N (.DIODE(net687));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_B1_N (.DIODE(net687));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_X (.DIODE(net687));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout339_A (.DIODE(net697));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_B1_1 (.DIODE(net697));
 sky130_fd_sc_hd__diode_2 ANTENNA_c267_X_1 (.DIODE(net697));
 sky130_fd_sc_hd__diode_2 ANTENNA_output144_A (.DIODE(net709));
 sky130_fd_sc_hd__diode_2 ANTENNA_c206_B (.DIODE(net709));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_B1_N (.DIODE(net709));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_B (.DIODE(net709));
 sky130_fd_sc_hd__diode_2 ANTENNA_c198_Y (.DIODE(net709));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout356_A (.DIODE(net713));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_A1_1 (.DIODE(net713));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_Y_1 (.DIODE(net713));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout350_A (.DIODE(net714));
 sky130_fd_sc_hd__diode_2 ANTENNA_output149_A_1 (.DIODE(net714));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge807_Q_1 (.DIODE(net714));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout288_A (.DIODE(net723));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A2_1 (.DIODE(net723));
 sky130_fd_sc_hd__diode_2 ANTENNA_c236_X_1 (.DIODE(net723));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout355_A (.DIODE(net726));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_A3_1 (.DIODE(net726));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_A1_1 (.DIODE(net726));
 sky130_fd_sc_hd__diode_2 ANTENNA_c240_B1_N_1 (.DIODE(net726));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_X_1 (.DIODE(net726));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout334_A (.DIODE(net732));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_A3_1 (.DIODE(net732));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_Y_1 (.DIODE(net732));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone76_A (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout306_A (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_A3_1 (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout182_X_1 (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap188_X (.DIODE(net753));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_A (.DIODE(net753));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_A2 (.DIODE(net753));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_A1 (.DIODE(net753));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout323_A (.DIODE(net757));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_A3_1 (.DIODE(net757));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap192_X_1 (.DIODE(net757));
 sky130_fd_sc_hd__diode_2 ANTENNA_c273_A (.DIODE(net764));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap199_X (.DIODE(net764));
 sky130_fd_sc_hd__diode_2 ANTENNA_c398_A2 (.DIODE(net764));
 sky130_fd_sc_hd__diode_2 ANTENNA_c271_B (.DIODE(net764));
 sky130_fd_sc_hd__diode_2 ANTENNA_c269_A (.DIODE(net764));
 sky130_fd_sc_hd__diode_2 ANTENNA_c267_B1_N (.DIODE(net764));
 sky130_fd_sc_hd__diode_2 ANTENNA_c270_A (.DIODE(net766));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap201_X (.DIODE(net766));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_A3 (.DIODE(net766));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_A (.DIODE(net766));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout351_A (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap202_X_1 (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_B1_1 (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_B1_N_1 (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_S1_1 (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout301_A (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_c760_S0_1 (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone5_X_1 (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer19_A (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer18_X (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c611_S0 (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer21_A (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer20_X (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_A2 (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_A1 (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_c191_B (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer30_A (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer29_X (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA_c536_A (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout284_X (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout283_A (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_B1_1 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_B1_1 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_A2_1 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c340_B1_N_1 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_B1_1 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_B1_N_1 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout294_X (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_output142_A_1 (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout293_A (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout175_A_1 (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_S0_1 (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_A3_1 (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_B1_1 (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_B1_N_1 (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_S1_1 (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c767_A3_1 (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_A3_1 (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout298_X (.DIODE(net1030));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_A2_1 (.DIODE(net1160));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_B_1 (.DIODE(net1160));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_A4_1 (.DIODE(net1160));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_B1_N_1 (.DIODE(net1030));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_B1_N_1 (.DIODE(net1160));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_S0_1 (.DIODE(net1030));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout297_A (.DIODE(net1030));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_A2_1 (.DIODE(net1030));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout308_X (.DIODE(net1040));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_S0_1 (.DIODE(net1040));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_B1_N_1 (.DIODE(net1040));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_A3_1 (.DIODE(net1040));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_A1_1 (.DIODE(net1040));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_B1_1 (.DIODE(net1040));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_A1 (.DIODE(net1047));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout315_X (.DIODE(net1047));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_A2_1 (.DIODE(net1047));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout314_A (.DIODE(net1047));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_A2_1 (.DIODE(net1047));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_S1_1 (.DIODE(net1047));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_B1_N_1 (.DIODE(net1047));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout329_X (.DIODE(net1061));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout328_A (.DIODE(net1061));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_B1_1 (.DIODE(net1061));
 sky130_fd_sc_hd__diode_2 ANTENNA_c691_B_1 (.DIODE(net1061));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_S1_1 (.DIODE(net1061));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_A3_1 (.DIODE(net1061));
 sky130_fd_sc_hd__diode_2 ANTENNA_c720_A2_1 (.DIODE(net1061));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout332_X (.DIODE(net1064));
 sky130_fd_sc_hd__diode_2 ANTENNA_c698_A2_1 (.DIODE(net1064));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A1_1 (.DIODE(net1064));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_A3_1 (.DIODE(net1064));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_A_1 (.DIODE(net1064));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout331_A (.DIODE(net1064));
 sky130_fd_sc_hd__diode_2 ANTENNA_c678_A2_1 (.DIODE(net1064));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout343_X (.DIODE(net1075));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_S1_1 (.DIODE(net1075));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_A3_1 (.DIODE(net1075));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_A3_1 (.DIODE(net1075));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_B1_1 (.DIODE(net1075));
 sky130_fd_sc_hd__diode_2 ANTENNA_c685_B1_N_1 (.DIODE(net1075));
 sky130_fd_sc_hd__diode_2 ANTENNA_c587_A0_1 (.DIODE(net1075));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_A2_1 (.DIODE(net1075));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout345_X (.DIODE(net1077));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_A1_1 (.DIODE(net1077));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_B1_N_1 (.DIODE(net1077));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_B_1 (.DIODE(net1077));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_B1_N_1 (.DIODE(net1077));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_A2_1 (.DIODE(net1077));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout354_X (.DIODE(net1086));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_B1_N_1 (.DIODE(net1086));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_S1_1 (.DIODE(net1086));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_B1_N_1 (.DIODE(net1086));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_A3_1 (.DIODE(net1086));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_S1_1 (.DIODE(net1086));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout353_A (.DIODE(net1086));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_B1_1 (.DIODE(net1086));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_B_1 (.DIODE(net1086));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout358_X (.DIODE(net1090));
 sky130_fd_sc_hd__diode_2 ANTENNA_c104_S1_1 (.DIODE(net1090));
 sky130_fd_sc_hd__diode_2 ANTENNA_c100_A3_1 (.DIODE(net1090));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout357_A (.DIODE(net1090));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout203_A_1 (.DIODE(net1090));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_B1_1 (.DIODE(net1090));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_A4_1 (.DIODE(net1090));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout374_X (.DIODE(net1106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_A2_1 (.DIODE(net1106));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout373_A (.DIODE(net1106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_A1_1 (.DIODE(net1106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c582_B1_N_1 (.DIODE(net1106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_A2_1 (.DIODE(net1106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A3_1 (.DIODE(net1106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_B1_1 (.DIODE(net1106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_S1_1 (.DIODE(net1106));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout377_X (.DIODE(net1109));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_A2_1 (.DIODE(net1109));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_A3_1 (.DIODE(net1109));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_A0_1 (.DIODE(net1109));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_A3_1 (.DIODE(net1109));
 sky130_fd_sc_hd__diode_2 ANTENNA_c110_A_1 (.DIODE(net1109));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout376_A (.DIODE(net1109));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_B_1 (.DIODE(net1110));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout378_X (.DIODE(net1110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c662_A_1 (.DIODE(net1110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_B1_N_1 (.DIODE(net1110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_A_1 (.DIODE(net1110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_A_1 (.DIODE(net1110));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout383_X (.DIODE(net1115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c496_B1_N_1 (.DIODE(net1115));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout382_A (.DIODE(net1115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c102_B1_N_1 (.DIODE(net1115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_B_1 (.DIODE(net1115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_A3_1 (.DIODE(net1115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_A2_1 (.DIODE(net1115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_B1_N_1 (.DIODE(net1115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_B_1 (.DIODE(net1115));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout386_X (.DIODE(net1118));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_A3_1 (.DIODE(net1118));
 sky130_fd_sc_hd__diode_2 ANTENNA_c208_B1_N_1 (.DIODE(net1118));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_B1_N_1 (.DIODE(net1118));
 sky130_fd_sc_hd__diode_2 ANTENNA_c373_A1_1 (.DIODE(net1118));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_A2_1 (.DIODE(net1118));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_B1_1 (.DIODE(net1118));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge792_S1_1 (.DIODE(net1118));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_B_1 (.DIODE(net1118));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_B_1 (.DIODE(net1118));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout385_A (.DIODE(net1118));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout388_X (.DIODE(net1120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_S0_1 (.DIODE(net1120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_A3_1 (.DIODE(net1120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_A3_1 (.DIODE(net1120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c669_A2_1 (.DIODE(net1120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c540_A_1 (.DIODE(net1120));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout387_A (.DIODE(net1120));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer64_A (.DIODE(net1131));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_B_1 (.DIODE(net1131));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer63_X (.DIODE(net1131));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_A_1 (.DIODE(net1141));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone22_A_1 (.DIODE(net1141));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer73_X (.DIODE(net1141));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(net686));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(net1054));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(net1055));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(net1100));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(net1104));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(net1105));
 sky130_fd_sc_hd__a31o_1 clone1 (.A1(net55),
    .A2(net22),
    .A3(net1056),
    .B1(net1107),
    .X(net1155));
 sky130_fd_sc_hd__clkbuf_1 clone2 (.A(net732),
    .X(net1156));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer75 (.A(net230),
    .X(net1157));
 sky130_fd_sc_hd__a21bo_1 clone77 (.A1(net31),
    .A2(net594),
    .B1_N(net43),
    .X(net1158));
 sky130_fd_sc_hd__xnor2_1 clone78 (.A(net750),
    .B(net764),
    .Y(net1159));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer83 (.A(net1030),
    .X(net1160));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer85 (.A(net344),
    .X(net1161));
 sky130_fd_sc_hd__a21bo_1 clone86 (.A1(net577),
    .A2(net1097),
    .B1_N(net21),
    .X(net1162));
 sky130_fd_sc_hd__clkbuf_1 clone87 (.A(net61),
    .X(net1163));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_594 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_328 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_255 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_189 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_384 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_438 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_456 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_583 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_403 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_494 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_609 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_443 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_303 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_331 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_592 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_609 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_415 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_490 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_311 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_47 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_239 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_609 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_219 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_424 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_392 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_275 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_594 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_606 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_606 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_578 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_611 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_618 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_308 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_413 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_244 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_273 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_301 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_368 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_599 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_283 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_423 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_42 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_355 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_469 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_311 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_382 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_12 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_142 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_594 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_64 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_163 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_619 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_400 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_619 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_23 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_32 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_591 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_272 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_394 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_443 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_484 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_540 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_609 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_272 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_382 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_270 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_512 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_133 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_239 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_459 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_59 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_609 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_469 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_114 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_60 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_609 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_619 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_367 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_20 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_431 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_191 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_242 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_413 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_25 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_328 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_8 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_112 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_387 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_435 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_395 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_239 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_426 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_422 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_143 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_303 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_617 ();
endmodule
