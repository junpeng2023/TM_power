module netlist_0 (clk,
    in0,
    in1,
    in10,
    in11,
    in12,
    in13,
    in14,
    in15,
    in16,
    in17,
    in18,
    in19,
    in2,
    in20,
    in21,
    in22,
    in23,
    in24,
    in25,
    in26,
    in27,
    in28,
    in29,
    in3,
    in30,
    in31,
    in32,
    in33,
    in34,
    in35,
    in36,
    in37,
    in38,
    in39,
    in4,
    in40,
    in41,
    in42,
    in43,
    in44,
    in45,
    in46,
    in47,
    in48,
    in49,
    in5,
    in50,
    in51,
    in52,
    in53,
    in54,
    in55,
    in56,
    in57,
    in58,
    in59,
    in6,
    in60,
    in61,
    in7,
    in8,
    in9,
    out0,
    out1,
    out10,
    out11,
    out12,
    out13,
    out14,
    out15,
    out16,
    out17,
    out18,
    out19,
    out2,
    out20,
    out21,
    out22,
    out23,
    out24,
    out25,
    out26,
    out27,
    out28,
    out29,
    out3,
    out30,
    out31,
    out32,
    out33,
    out34,
    out35,
    out36,
    out37,
    out38,
    out39,
    out4,
    out40,
    out41,
    out42,
    out43,
    out44,
    out45,
    out46,
    out47,
    out48,
    out49,
    out5,
    out50,
    out51,
    out52,
    out53,
    out54,
    out55,
    out56,
    out57,
    out58,
    out59,
    out6,
    out60,
    out61,
    out7,
    out8,
    out9,
    rst);
 input clk;
 input in0;
 input in1;
 input in10;
 input in11;
 input in12;
 input in13;
 input in14;
 input in15;
 input in16;
 input in17;
 input in18;
 input in19;
 input in2;
 input in20;
 input in21;
 input in22;
 input in23;
 input in24;
 input in25;
 input in26;
 input in27;
 input in28;
 input in29;
 input in3;
 input in30;
 input in31;
 input in32;
 input in33;
 input in34;
 input in35;
 input in36;
 input in37;
 input in38;
 input in39;
 input in4;
 input in40;
 input in41;
 input in42;
 input in43;
 input in44;
 input in45;
 input in46;
 input in47;
 input in48;
 input in49;
 input in5;
 input in50;
 input in51;
 input in52;
 input in53;
 input in54;
 input in55;
 input in56;
 input in57;
 input in58;
 input in59;
 input in6;
 input in60;
 input in61;
 input in7;
 input in8;
 input in9;
 output out0;
 output out1;
 output out10;
 output out11;
 output out12;
 output out13;
 output out14;
 output out15;
 output out16;
 output out17;
 output out18;
 output out19;
 output out2;
 output out20;
 output out21;
 output out22;
 output out23;
 output out24;
 output out25;
 output out26;
 output out27;
 output out28;
 output out29;
 output out3;
 output out30;
 output out31;
 output out32;
 output out33;
 output out34;
 output out35;
 output out36;
 output out37;
 output out38;
 output out39;
 output out4;
 output out40;
 output out41;
 output out42;
 output out43;
 output out44;
 output out45;
 output out46;
 output out47;
 output out48;
 output out49;
 output out5;
 output out50;
 output out51;
 output out52;
 output out53;
 output out54;
 output out55;
 output out56;
 output out57;
 output out58;
 output out59;
 output out6;
 output out60;
 output out61;
 output out7;
 output out8;
 output out9;
 input rst;

 wire net0;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net63;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net64;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net65;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net66;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net67;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net68;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net69;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net7;
 wire net70;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net71;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net72;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net73;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net74;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net75;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net76;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net77;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net78;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net79;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net8;
 wire net80;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net81;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net82;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net83;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net84;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net85;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net86;
 wire net860;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net133;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_0_net854;
 wire clknet_1_0__leaf_net854;
 wire clknet_1_1__leaf_net854;
 wire clknet_0_net706;
 wire clknet_1_0__leaf_net706;
 wire clknet_1_1__leaf_net706;
 wire clknet_0_net623;
 wire clknet_1_0__leaf_net623;
 wire clknet_1_1__leaf_net623;
 wire clknet_0_net585;
 wire clknet_1_0__leaf_net585;
 wire clknet_1_1__leaf_net585;
 wire clknet_0_net425;
 wire clknet_1_0__leaf_net425;
 wire clknet_1_1__leaf_net425;
 wire clknet_0_net433;
 wire clknet_1_0__leaf_net433;
 wire clknet_1_1__leaf_net433;
 wire clknet_0_net423;
 wire clknet_1_0__leaf_net423;
 wire clknet_1_1__leaf_net423;
 wire clknet_0_net934;
 wire clknet_1_0__leaf_net934;
 wire clknet_1_1__leaf_net934;
 wire clknet_0_net517;
 wire clknet_1_0__leaf_net517;
 wire clknet_1_1__leaf_net517;
 wire clknet_0_net490;
 wire clknet_1_0__leaf_net490;
 wire clknet_1_1__leaf_net490;
 wire clknet_0_net493;
 wire clknet_1_0__leaf_net493;
 wire clknet_1_1__leaf_net493;
 wire clknet_0_net835;
 wire clknet_1_0__leaf_net835;
 wire clknet_1_1__leaf_net835;
 wire clknet_0_net499;
 wire clknet_1_0__leaf_net499;
 wire clknet_1_1__leaf_net499;
 wire clknet_0_net498;
 wire clknet_1_0__leaf_net498;
 wire clknet_1_1__leaf_net498;
 wire clknet_0_net833;
 wire clknet_1_0__leaf_net833;
 wire clknet_1_1__leaf_net833;
 wire clknet_0_net973;
 wire clknet_1_0__leaf_net973;
 wire clknet_1_1__leaf_net973;
 wire clknet_0_net922;
 wire clknet_1_0__leaf_net922;
 wire clknet_1_1__leaf_net922;
 wire clknet_0_net522;
 wire clknet_1_0__leaf_net522;
 wire clknet_1_1__leaf_net522;
 wire clknet_0_net617;
 wire clknet_1_0__leaf_net617;
 wire clknet_1_1__leaf_net617;
 wire clknet_0_net834;
 wire clknet_1_0__leaf_net834;
 wire clknet_1_1__leaf_net834;
 wire clknet_0_net508;
 wire clknet_1_0__leaf_net508;
 wire clknet_1_1__leaf_net508;
 wire clknet_0_net510;
 wire clknet_1_0__leaf_net510;
 wire clknet_1_1__leaf_net510;
 wire clknet_0_net515;
 wire clknet_1_0__leaf_net515;
 wire clknet_1_1__leaf_net515;
 wire clknet_0_net483;
 wire clknet_1_0__leaf_net483;
 wire clknet_1_1__leaf_net483;
 wire clknet_0_net606;
 wire clknet_1_0__leaf_net606;
 wire clknet_1_1__leaf_net606;
 wire clknet_0_net465;
 wire clknet_1_0__leaf_net465;
 wire clknet_1_1__leaf_net465;
 wire clknet_0_net471;
 wire clknet_1_0__leaf_net471;
 wire clknet_1_1__leaf_net471;
 wire clknet_0_net461;
 wire clknet_1_0__leaf_net461;
 wire clknet_1_1__leaf_net461;
 wire clknet_0_net474;
 wire clknet_1_0__leaf_net474;
 wire clknet_1_1__leaf_net474;
 wire clknet_0_net853;
 wire clknet_1_0__leaf_net853;
 wire clknet_1_1__leaf_net853;
 wire clknet_0_net604;
 wire clknet_1_0__leaf_net604;
 wire clknet_1_1__leaf_net604;
 wire clknet_0_net591;
 wire clknet_1_0__leaf_net591;
 wire clknet_1_1__leaf_net591;
 wire clknet_0_net469;
 wire clknet_1_0__leaf_net469;
 wire clknet_1_1__leaf_net469;
 wire clknet_0_net852;
 wire clknet_1_0__leaf_net852;
 wire clknet_1_1__leaf_net852;
 wire clknet_0_net595;
 wire clknet_1_0__leaf_net595;
 wire clknet_1_1__leaf_net595;
 wire clknet_0_net924;
 wire clknet_1_0__leaf_net924;
 wire clknet_1_1__leaf_net924;
 wire clknet_0_net815;
 wire clknet_1_0__leaf_net815;
 wire clknet_1_1__leaf_net815;
 wire clknet_0_net927;
 wire clknet_1_0__leaf_net927;
 wire clknet_1_1__leaf_net927;
 wire clknet_0_net506;
 wire clknet_1_0__leaf_net506;
 wire clknet_1_1__leaf_net506;
 wire clknet_0_net954;
 wire clknet_1_0__leaf_net954;
 wire clknet_1_1__leaf_net954;
 wire clknet_0_net938;
 wire clknet_1_0__leaf_net938;
 wire clknet_1_1__leaf_net938;
 wire clknet_0_net977;
 wire clknet_1_0__leaf_net977;
 wire clknet_1_1__leaf_net977;
 wire clknet_0_net799;
 wire clknet_1_0__leaf_net799;
 wire clknet_1_1__leaf_net799;
 wire clknet_0_net330;
 wire clknet_1_0__leaf_net330;
 wire clknet_1_1__leaf_net330;
 wire clknet_0_net798;
 wire clknet_1_0__leaf_net798;
 wire clknet_1_1__leaf_net798;
 wire clknet_0_net303;
 wire clknet_1_0__leaf_net303;
 wire clknet_1_1__leaf_net303;
 wire clknet_0_net705;
 wire clknet_1_0__leaf_net705;
 wire clknet_1_1__leaf_net705;
 wire clknet_0_net302;
 wire clknet_1_0__leaf_net302;
 wire clknet_1_1__leaf_net302;
 wire clknet_0_net946;
 wire clknet_1_0__leaf_net946;
 wire clknet_1_1__leaf_net946;
 wire clknet_0_net397;
 wire clknet_1_0__leaf_net397;
 wire clknet_1_1__leaf_net397;
 wire clknet_0_net386;
 wire clknet_1_0__leaf_net386;
 wire clknet_1_1__leaf_net386;
 wire clknet_0_net952;
 wire clknet_1_0__leaf_net952;
 wire clknet_1_1__leaf_net952;
 wire clknet_0_net282;
 wire clknet_1_0__leaf_net282;
 wire clknet_1_1__leaf_net282;
 wire clknet_0_net761;
 wire clknet_1_0__leaf_net761;
 wire clknet_1_1__leaf_net761;
 wire clknet_0_net191;
 wire clknet_1_0__leaf_net191;
 wire clknet_1_1__leaf_net191;
 wire clknet_0_net743;
 wire clknet_1_0__leaf_net743;
 wire clknet_1_1__leaf_net743;
 wire clknet_0_net49;
 wire clknet_1_0__leaf_net49;
 wire clknet_1_1__leaf_net49;
 wire clknet_0_net971;
 wire clknet_1_0__leaf_net971;
 wire clknet_1_1__leaf_net971;
 wire clknet_0_net52;
 wire clknet_1_0__leaf_net52;
 wire clknet_1_1__leaf_net52;
 wire clknet_0_net57;
 wire clknet_1_0__leaf_net57;
 wire clknet_1_1__leaf_net57;
 wire clknet_0_net744;
 wire clknet_1_0__leaf_net744;
 wire clknet_1_1__leaf_net744;
 wire clknet_0_net179;
 wire clknet_1_0__leaf_net179;
 wire clknet_1_1__leaf_net179;
 wire clknet_0_net181;
 wire clknet_1_0__leaf_net181;
 wire clknet_1_1__leaf_net181;
 wire clknet_0_net937;
 wire clknet_1_0__leaf_net937;
 wire clknet_1_1__leaf_net937;
 wire clknet_0_net972;
 wire clknet_1_0__leaf_net972;
 wire clknet_1_1__leaf_net972;
 wire clknet_0_net153;
 wire clknet_1_0__leaf_net153;
 wire clknet_1_1__leaf_net153;
 wire clknet_0_net797;
 wire clknet_1_0__leaf_net797;
 wire clknet_1_1__leaf_net797;
 wire clknet_0_net947;
 wire clknet_1_0__leaf_net947;
 wire clknet_1_1__leaf_net947;
 wire clknet_0_net401;
 wire clknet_1_0__leaf_net401;
 wire clknet_1_1__leaf_net401;
 wire clknet_0_net945;
 wire clknet_1_0__leaf_net945;
 wire clknet_1_1__leaf_net945;
 wire clknet_0_net403;
 wire clknet_1_0__leaf_net403;
 wire clknet_1_1__leaf_net403;
 wire clknet_0_net300;
 wire clknet_1_0__leaf_net300;
 wire clknet_1_1__leaf_net300;
 wire clknet_0_net145;
 wire clknet_1_0__leaf_net145;
 wire clknet_1_1__leaf_net145;
 wire clknet_0_net62;
 wire clknet_1_0__leaf_net62;
 wire clknet_1_1__leaf_net62;
 wire clknet_0_net182;
 wire clknet_1_0__leaf_net182;
 wire clknet_1_1__leaf_net182;
 wire clknet_0_net188;
 wire clknet_1_0__leaf_net188;
 wire clknet_1_1__leaf_net188;
 wire clknet_0_net185;
 wire clknet_1_0__leaf_net185;
 wire clknet_1_1__leaf_net185;
 wire clknet_0_net184;
 wire clknet_1_0__leaf_net184;
 wire clknet_1_1__leaf_net184;
 wire clknet_0_net67;
 wire clknet_1_0__leaf_net67;
 wire clknet_1_1__leaf_net67;
 wire clknet_0_net959;
 wire clknet_1_0__leaf_net959;
 wire clknet_1_1__leaf_net959;
 wire clknet_0_net974;
 wire clknet_1_0__leaf_net974;
 wire clknet_1_1__leaf_net974;
 wire clknet_0_net177;
 wire clknet_1_0__leaf_net177;
 wire clknet_1_1__leaf_net177;
 wire clknet_0_net60;
 wire clknet_1_0__leaf_net60;
 wire clknet_1_1__leaf_net60;
 wire clknet_0_net56;
 wire clknet_1_0__leaf_net56;
 wire clknet_1_1__leaf_net56;
 wire clknet_0_net965;
 wire clknet_1_0__leaf_net965;
 wire clknet_1_1__leaf_net965;
 wire clknet_0_net54;
 wire clknet_1_0__leaf_net54;
 wire clknet_1_1__leaf_net54;
 wire clknet_0_net48;
 wire clknet_1_0__leaf_net48;
 wire clknet_1_1__leaf_net48;
 wire clknet_0_net50;
 wire clknet_1_0__leaf_net50;
 wire clknet_1_1__leaf_net50;
 wire clknet_0_net171;
 wire clknet_1_0__leaf_net171;
 wire clknet_1_1__leaf_net171;
 wire clknet_0_net957;
 wire clknet_1_0__leaf_net957;
 wire clknet_1_1__leaf_net957;
 wire clknet_0_net762;
 wire clknet_1_0__leaf_net762;
 wire clknet_1_1__leaf_net762;
 wire clknet_0_net780;
 wire clknet_1_0__leaf_net780;
 wire clknet_1_1__leaf_net780;
 wire clknet_0_net273;
 wire clknet_1_0__leaf_net273;
 wire clknet_1_1__leaf_net273;
 wire clknet_0_net275;
 wire clknet_1_0__leaf_net275;
 wire clknet_1_1__leaf_net275;
 wire clknet_0_net251;
 wire clknet_1_0__leaf_net251;
 wire clknet_1_1__leaf_net251;
 wire clknet_0_net257;
 wire clknet_1_0__leaf_net257;
 wire clknet_1_1__leaf_net257;
 wire clknet_0_net253;
 wire clknet_1_0__leaf_net253;
 wire clknet_1_1__leaf_net253;
 wire clknet_0_net246;
 wire clknet_1_0__leaf_net246;
 wire clknet_1_1__leaf_net246;
 wire clknet_0_net475;
 wire clknet_1_0__leaf_net475;
 wire clknet_1_1__leaf_net475;
 wire clknet_0_net462;
 wire clknet_1_0__leaf_net462;
 wire clknet_1_1__leaf_net462;
 wire clknet_0_net369;
 wire clknet_1_0__leaf_net369;
 wire clknet_1_1__leaf_net369;
 wire clknet_0_net245;
 wire clknet_1_0__leaf_net245;
 wire clknet_1_1__leaf_net245;
 wire clknet_0_net396;
 wire clknet_1_0__leaf_net396;
 wire clknet_1_1__leaf_net396;
 wire clknet_0_net779;
 wire clknet_1_0__leaf_net779;
 wire clknet_1_1__leaf_net779;
 wire clknet_0_net250;
 wire clknet_1_0__leaf_net250;
 wire clknet_1_1__leaf_net250;
 wire clknet_0_net778;
 wire clknet_1_0__leaf_net778;
 wire clknet_1_1__leaf_net778;
 wire clknet_0_net238;
 wire clknet_1_0__leaf_net238;
 wire clknet_1_1__leaf_net238;
 wire clknet_0_net332;
 wire clknet_1_0__leaf_net332;
 wire clknet_1_1__leaf_net332;
 wire clknet_0_net331;
 wire clknet_1_0__leaf_net331;
 wire clknet_1_1__leaf_net331;
 wire clknet_0_net760;
 wire clknet_1_0__leaf_net760;
 wire clknet_1_1__leaf_net760;
 wire clknet_0_net742;
 wire clknet_1_0__leaf_net742;
 wire clknet_1_1__leaf_net742;
 wire clknet_0_net562;
 wire clknet_1_0__leaf_net562;
 wire clknet_1_1__leaf_net562;
 wire clknet_0_net560;
 wire clknet_1_0__leaf_net560;
 wire clknet_1_1__leaf_net560;
 wire clknet_0_net568;
 wire clknet_1_0__leaf_net568;
 wire clknet_1_1__leaf_net568;
 wire clknet_0_net542;
 wire clknet_1_0__leaf_net542;
 wire clknet_1_1__leaf_net542;
 wire clknet_0_net592;
 wire clknet_1_0__leaf_net592;
 wire clknet_1_1__leaf_net592;
 wire clknet_0_net552;
 wire clknet_1_0__leaf_net552;
 wire clknet_1_1__leaf_net552;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;

 sky130_fd_sc_hd__a41o_2 c100 (.A1(net28),
    .A2(net15),
    .A3(net26),
    .A4(net35),
    .B1(net1009),
    .X(net38));
 sky130_fd_sc_hd__a21bo_1 c101 (.A1(net38),
    .A2(net29),
    .B1_N(net1009),
    .X(net39));
 sky130_fd_sc_hd__sdfbbn_2 c102 (.CLK_N(clknet_4_14_0_clk),
    .D(net37),
    .RESET_B(net39),
    .SCD(net38),
    .SCE(net998),
    .SET_B(net1009),
    .Q(net969),
    .Q_N(net40));
 sky130_fd_sc_hd__a41o_1 c103 (.A1(net39),
    .A2(net31),
    .A3(net969),
    .A4(net38),
    .B1(net1009),
    .X(net41));
 sky130_fd_sc_hd__a41o_1 c104 (.A1(net33),
    .A2(net969),
    .A3(net38),
    .A4(net943),
    .B1(net873),
    .X(net42));
 sky130_fd_sc_hd__mux4_1 c105 (.A0(net32),
    .A1(net4),
    .A2(net39),
    .A3(net40),
    .S0(net33),
    .S1(net1044),
    .X(net43));
 sky130_fd_sc_hd__sdfbbn_1 c106 (.CLK_N(clknet_4_14_0_clk),
    .D(net31),
    .RESET_B(net1085),
    .SCD(net42),
    .SCE(net38),
    .SET_B(net37),
    .Q(net45),
    .Q_N(net44));
 sky130_fd_sc_hd__a41o_1 c107 (.A1(net900),
    .A2(net969),
    .A3(net1009),
    .A4(net702),
    .B1(net755),
    .X(net46));
 sky130_fd_sc_hd__mux4_2 c108 (.A0(net45),
    .A1(net969),
    .A2(net46),
    .A3(net29),
    .S0(net1009),
    .S1(net702),
    .X(net967));
 sky130_fd_sc_hd__mux4_1 c109 (.A0(net42),
    .A1(net46),
    .A2(net967),
    .A3(net44),
    .S0(net40),
    .S1(net702),
    .X(net47));
 sky130_fd_sc_hd__buf_1 c110 (.A(clknet_1_1__leaf_net743),
    .X(net48));
 sky130_fd_sc_hd__buf_1 c111 (.A(clknet_1_1__leaf_net743),
    .X(net49));
 sky130_fd_sc_hd__a21bo_1 c112 (.A1(net22),
    .A2(clknet_1_0__leaf_net48),
    .B1_N(net40),
    .X(net50));
 sky130_fd_sc_hd__dfbbn_2 c113 (.CLK_N(clknet_4_15_0_clk),
    .D(clknet_1_1__leaf_net48),
    .RESET_B(net967),
    .SET_B(net943),
    .Q(net942),
    .Q_N(net51));
 sky130_fd_sc_hd__a21bo_1 c114 (.A1(net15),
    .A2(clknet_1_0__leaf_net48),
    .B1_N(net1044),
    .X(net958));
 sky130_fd_sc_hd__a21bo_1 c115 (.A1(net1035),
    .A2(clknet_1_1__leaf_net48),
    .B1_N(clknet_1_1__leaf_net49),
    .X(net52));
 sky130_fd_sc_hd__a21bo_1 c116 (.A1(net45),
    .A2(net1032),
    .B1_N(clknet_1_1__leaf_net52),
    .X(net959));
 sky130_fd_sc_hd__mux4_1 c117 (.A0(net32),
    .A1(net1044),
    .A2(net942),
    .A3(clknet_1_1__leaf_net959),
    .S0(clknet_1_1__leaf_net48),
    .S1(net31),
    .X(net53));
 sky130_fd_sc_hd__a31o_1 c118 (.A1(net1032),
    .A2(clknet_1_1__leaf_net959),
    .A3(net51),
    .B1(net756),
    .X(net54));
 sky130_fd_sc_hd__a41o_1 c119 (.A1(clknet_1_0__leaf_net959),
    .A2(net1040),
    .A3(net1032),
    .A4(clknet_1_1__leaf_net48),
    .B1(net949),
    .X(net965));
 sky130_fd_sc_hd__a41o_1 c120 (.A1(clknet_1_1__leaf_net50),
    .A2(clknet_1_0__leaf_net48),
    .A3(net1035),
    .A4(clknet_1_1__leaf_net959),
    .B1(net942),
    .X(net55));
 sky130_fd_sc_hd__a21bo_1 c121 (.A1(clknet_1_1__leaf_net54),
    .A2(clknet_1_1__leaf_net959),
    .B1_N(net943),
    .X(net56));
 sky130_fd_sc_hd__a41o_1 c122 (.A1(clknet_1_0__leaf_net52),
    .A2(net5),
    .A3(net942),
    .A4(clknet_1_0__leaf_net56),
    .B1(clknet_1_1__leaf_net48),
    .X(net57));
 sky130_fd_sc_hd__a21bo_1 c123 (.A1(clknet_1_1__leaf_net48),
    .A2(clknet_1_1__leaf_net959),
    .B1_N(net17),
    .X(net58));
 sky130_fd_sc_hd__mux4_1 c124 (.A0(net55),
    .A1(net32),
    .A2(clknet_1_0__leaf_net52),
    .A3(clknet_1_1__leaf_net56),
    .S0(clknet_1_0__leaf_net54),
    .S1(clknet_1_1__leaf_net959),
    .X(net59));
 sky130_fd_sc_hd__a41o_1 c125 (.A1(net10),
    .A2(net942),
    .A3(clknet_1_0__leaf_net48),
    .A4(clknet_1_1__leaf_net959),
    .B1(clknet_1_0__leaf_net50),
    .X(net60));
 sky130_fd_sc_hd__a31o_1 c126 (.A1(clknet_1_0__leaf_net60),
    .A2(clknet_1_1__leaf_net959),
    .A3(net1055),
    .B1(net17),
    .X(net61));
 sky130_fd_sc_hd__mux4_1 c127 (.A0(clknet_1_0__leaf_net57),
    .A1(net22),
    .A2(net15),
    .A3(clknet_1_0__leaf_net48),
    .S0(clknet_1_0__leaf_net60),
    .S1(net1040),
    .X(net62));
 sky130_fd_sc_hd__a41o_1 c128 (.A1(net58),
    .A2(net51),
    .A3(clknet_1_0__leaf_net62),
    .A4(clknet_1_1__leaf_net57),
    .B1(net967),
    .X(net63));
 sky130_fd_sc_hd__sdfbbp_1 c129 (.CLK(clknet_4_15_0_clk),
    .D(net61),
    .RESET_B(clknet_1_0__leaf_net62),
    .SCD(net31),
    .SCE(clknet_1_0__leaf_net959),
    .SET_B(clknet_1_1__leaf_net744),
    .Q(net65),
    .Q_N(net64));
 sky130_fd_sc_hd__a31o_1 c130 (.A1(clknet_1_0__leaf_net56),
    .A2(clknet_1_0__leaf_net62),
    .A3(clknet_1_1__leaf_net959),
    .B1(net64),
    .X(net66));
 sky130_fd_sc_hd__mux4_1 c131 (.A0(net66),
    .A1(net1040),
    .A2(clknet_1_0__leaf_net62),
    .A3(clknet_1_0__leaf_net965),
    .S0(clknet_1_1__leaf_net60),
    .S1(clknet_1_0__leaf_net959),
    .X(net67));
 sky130_fd_sc_hd__a21bo_4 c132 (.A1(net916),
    .A2(net861),
    .B1_N(net1049),
    .X(net68));
 sky130_fd_sc_hd__a21bo_4 c133 (.A1(net916),
    .A2(net920),
    .B1_N(net1034),
    .X(net69));
 sky130_fd_sc_hd__a41o_4 c134 (.A1(net1034),
    .A2(net921),
    .A3(net871),
    .A4(net1042),
    .B1(net920),
    .X(net70));
 sky130_fd_sc_hd__a21bo_1 c135 (.A1(net905),
    .A2(net862),
    .B1_N(net1049),
    .X(net71));
 sky130_fd_sc_hd__a41o_4 c136 (.A1(net863),
    .A2(net69),
    .A3(net71),
    .A4(net1049),
    .B1(net1020),
    .X(net72));
 sky130_fd_sc_hd__a41o_4 c137 (.A1(net864),
    .A2(net1049),
    .A3(net883),
    .A4(net1020),
    .B1(net1006),
    .X(net73));
 sky130_fd_sc_hd__a21bo_4 c138 (.A1(net1034),
    .A2(net69),
    .B1_N(net1006),
    .X(net74));
 sky130_fd_sc_hd__a41o_1 c139 (.A1(net74),
    .A2(net866),
    .A3(net861),
    .A4(net1034),
    .B1(net1058),
    .X(net75));
 sky130_fd_sc_hd__a31o_4 c140 (.A1(net73),
    .A2(net69),
    .A3(net866),
    .B1(net1049),
    .X(net76));
 sky130_fd_sc_hd__mux4_2 c141 (.A0(net862),
    .A1(net71),
    .A2(net868),
    .A3(net76),
    .S0(net74),
    .S1(net1006),
    .X(net77));
 sky130_fd_sc_hd__a41o_4 c142 (.A1(net73),
    .A2(net74),
    .A3(net861),
    .A4(net1042),
    .B1(net1058),
    .X(net78));
 sky130_fd_sc_hd__a41o_1 c143 (.A1(net71),
    .A2(net74),
    .A3(net920),
    .A4(net69),
    .B1(net1058),
    .X(net79));
 sky130_fd_sc_hd__a41o_4 c144 (.A1(net861),
    .A2(net1006),
    .A3(net1020),
    .A4(net1034),
    .B1(net74),
    .X(net80));
 sky130_fd_sc_hd__a41o_4 c145 (.A1(net75),
    .A2(net73),
    .A3(net80),
    .A4(net79),
    .B1(net1004),
    .X(net81));
 sky130_fd_sc_hd__a41o_4 c146 (.A1(net79),
    .A2(net867),
    .A3(net1004),
    .A4(net74),
    .B1(net1001),
    .X(net82));
 sky130_fd_sc_hd__a41o_2 c147 (.A1(net867),
    .A2(net874),
    .A3(net1020),
    .A4(net1035),
    .B1(net80),
    .X(net83));
 sky130_fd_sc_hd__a41o_4 c148 (.A1(net82),
    .A2(net920),
    .A3(net80),
    .A4(net866),
    .B1(net905),
    .X(net84));
 sky130_fd_sc_hd__mux4_2 c149 (.A0(net69),
    .A1(net76),
    .A2(net79),
    .A3(net1004),
    .S0(net1064),
    .S1(net74),
    .X(net85));
 sky130_fd_sc_hd__a41o_1 c150 (.A1(net921),
    .A2(net871),
    .A3(net1064),
    .A4(net1004),
    .B1(net80),
    .X(net86));
 sky130_fd_sc_hd__a41o_1 c151 (.A1(net86),
    .A2(net864),
    .A3(net1050),
    .A4(net1001),
    .B1(net1004),
    .X(net87));
 sky130_fd_sc_hd__mux4_2 c152 (.A0(net83),
    .A1(net87),
    .A2(net80),
    .A3(net86),
    .S0(net1006),
    .S1(net69),
    .X(net88));
 sky130_fd_sc_hd__mux4_2 c153 (.A0(net88),
    .A1(net920),
    .A2(net87),
    .A3(net1063),
    .S0(net69),
    .S1(net86),
    .X(net89));
 sky130_fd_sc_hd__a41o_4 c154 (.A1(net84),
    .A2(net884),
    .A3(net85),
    .A4(net1050),
    .B1(net1045),
    .X(net90));
 sky130_fd_sc_hd__a31o_1 c155 (.A1(net874),
    .A2(net889),
    .A3(net996),
    .B1(net1071),
    .X(net91));
 sky130_fd_sc_hd__a41o_2 c156 (.A1(net869),
    .A2(net87),
    .A3(net80),
    .A4(net1044),
    .B1(net875),
    .X(net92));
 sky130_fd_sc_hd__a31o_1 c157 (.A1(net895),
    .A2(net896),
    .A3(net1042),
    .B1(net882),
    .X(net93));
 sky130_fd_sc_hd__mux4_2 c158 (.A0(net893),
    .A1(net875),
    .A2(net996),
    .A3(net1071),
    .S0(net93),
    .S1(net880),
    .X(net94));
 sky130_fd_sc_hd__mux4_2 c159 (.A0(net91),
    .A1(net94),
    .A2(net996),
    .A3(net93),
    .S0(net76),
    .S1(net1064),
    .X(net95));
 sky130_fd_sc_hd__a41o_2 c160 (.A1(net877),
    .A2(net879),
    .A3(net92),
    .A4(net1064),
    .B1(net897),
    .X(net96));
 sky130_fd_sc_hd__a31o_2 c161 (.A1(net870),
    .A2(net876),
    .A3(net886),
    .B1(net69),
    .X(net97));
 sky130_fd_sc_hd__a31o_4 c162 (.A1(net97),
    .A2(net879),
    .A3(net1051),
    .B1(net877),
    .X(net98));
 sky130_fd_sc_hd__a41o_2 c163 (.A1(net1044),
    .A2(net876),
    .A3(net80),
    .A4(net1042),
    .B1(net98),
    .X(net99));
 sky130_fd_sc_hd__a41o_1 c164 (.A1(net94),
    .A2(net93),
    .A3(net85),
    .A4(net1066),
    .B1(net878),
    .X(net100));
 sky130_fd_sc_hd__a21bo_1 c165 (.A1(net100),
    .A2(net877),
    .B1_N(net95),
    .X(net101));
 sky130_fd_sc_hd__mux4_1 c166 (.A0(net898),
    .A1(net1005),
    .A2(net92),
    .A3(net1042),
    .S0(net94),
    .S1(net100),
    .X(net102));
 sky130_fd_sc_hd__mux4_1 c167 (.A0(net102),
    .A1(net100),
    .A2(net91),
    .A3(net879),
    .S0(net87),
    .S1(net80),
    .X(net103));
 sky130_fd_sc_hd__a41o_2 c168 (.A1(net883),
    .A2(net91),
    .A3(net101),
    .A4(net1044),
    .B1(net96),
    .X(net104));
 sky130_fd_sc_hd__mux4_2 c169 (.A0(net101),
    .A1(net870),
    .A2(net879),
    .A3(net98),
    .S0(net988),
    .S1(net893),
    .X(net105));
 sky130_fd_sc_hd__mux4_2 c170 (.A0(net87),
    .A1(net102),
    .A2(net103),
    .A3(net94),
    .S0(net893),
    .S1(net101),
    .X(net106));
 sky130_fd_sc_hd__a41o_1 c171 (.A1(net92),
    .A2(net106),
    .A3(net988),
    .A4(net99),
    .B1(net101),
    .X(net107));
 sky130_fd_sc_hd__mux4_1 c172 (.A0(net875),
    .A1(net105),
    .A2(net99),
    .A3(net106),
    .S0(net94),
    .S1(net107),
    .X(net108));
 sky130_fd_sc_hd__mux4_1 c173 (.A0(net103),
    .A1(net105),
    .A2(net102),
    .A3(net107),
    .S0(net96),
    .S1(net106),
    .X(net109));
 sky130_fd_sc_hd__mux4_1 c174 (.A0(net106),
    .A1(net1064),
    .A2(net996),
    .A3(net107),
    .S0(net1030),
    .S1(net758),
    .X(net110));
 sky130_fd_sc_hd__mux4_1 c175 (.A0(net93),
    .A1(net101),
    .A2(net103),
    .A3(net107),
    .S0(net98),
    .S1(net105),
    .X(net111));
 sky130_fd_sc_hd__a21bo_2 c176 (.A1(net1),
    .A2(net99),
    .B1_N(net886),
    .X(net112));
 sky130_fd_sc_hd__a31o_4 c177 (.A1(net1071),
    .A2(net996),
    .A3(net1038),
    .B1(net757),
    .X(net113));
 sky130_fd_sc_hd__a31o_1 c178 (.A1(net879),
    .A2(net107),
    .A3(net113),
    .B1(net909),
    .X(net114));
 sky130_fd_sc_hd__a41o_2 c179 (.A1(net98),
    .A2(net1),
    .A3(net1040),
    .A4(net1038),
    .B1(net1028),
    .X(net115));
 sky130_fd_sc_hd__mux4_2 c180 (.A0(net868),
    .A1(net92),
    .A2(net1038),
    .A3(net99),
    .S0(net1003),
    .S1(net1028),
    .X(net116));
 sky130_fd_sc_hd__mux4_2 c181 (.A0(net911),
    .A1(net878),
    .A2(net89),
    .A3(net1036),
    .S0(net1003),
    .S1(net750),
    .X(net117));
 sky130_fd_sc_hd__a31o_1 c182 (.A1(net105),
    .A2(net98),
    .A3(net85),
    .B1(net1050),
    .X(net118));
 sky130_fd_sc_hd__mux4_2 c183 (.A0(net1042),
    .A1(net115),
    .A2(net1036),
    .A3(net112),
    .S0(net92),
    .S1(net1028),
    .X(net119));
 sky130_fd_sc_hd__mux4_1 c184 (.A0(net119),
    .A1(net116),
    .A2(net118),
    .A3(net1003),
    .S0(net117),
    .S1(net1019),
    .X(net120));
 sky130_fd_sc_hd__mux4_2 c185 (.A0(net89),
    .A1(net112),
    .A2(net3),
    .A3(net106),
    .S0(net911),
    .S1(net119),
    .X(net121));
 sky130_fd_sc_hd__a41o_1 c186 (.A1(net886),
    .A2(net894),
    .A3(net99),
    .A4(net1002),
    .B1(net1027),
    .X(net122));
 sky130_fd_sc_hd__a21bo_2 c187 (.A1(net113),
    .A2(net112),
    .B1_N(net1043),
    .X(net123));
 sky130_fd_sc_hd__mux4_2 c188 (.A0(net906),
    .A1(net1005),
    .A2(net123),
    .A3(net879),
    .S0(net1000),
    .S1(net1027),
    .X(net124));
 sky130_fd_sc_hd__a41o_1 c189 (.A1(net107),
    .A2(net121),
    .A3(net894),
    .A4(net116),
    .B1(net123),
    .X(net125));
 sky130_fd_sc_hd__a31o_1 c190 (.A1(net123),
    .A2(net124),
    .A3(net878),
    .B1(net118),
    .X(net126));
 sky130_fd_sc_hd__mux4_2 c191 (.A0(net123),
    .A1(net124),
    .A2(net113),
    .A3(net1000),
    .S0(net643),
    .S1(net1027),
    .X(net127));
 sky130_fd_sc_hd__a41o_1 c192 (.A1(net116),
    .A2(net117),
    .A3(net127),
    .A4(net112),
    .B1(net643),
    .X(net128));
 sky130_fd_sc_hd__mux4_2 c193 (.A0(net123),
    .A1(net124),
    .A2(net119),
    .A3(net1005),
    .S0(net643),
    .S1(net1028),
    .X(net129));
 sky130_fd_sc_hd__mux4_2 c194 (.A0(net1000),
    .A1(net906),
    .A2(net1045),
    .A3(net117),
    .S0(net127),
    .S1(net644),
    .X(net130));
 sky130_fd_sc_hd__mux4_2 c195 (.A0(net128),
    .A1(net95),
    .A2(net129),
    .A3(net106),
    .S0(net123),
    .S1(net124),
    .X(net131));
 sky130_fd_sc_hd__mux4_1 c196 (.A0(net121),
    .A1(net131),
    .A2(net129),
    .A3(net119),
    .S0(net105),
    .S1(net643),
    .X(net132));
 sky130_fd_sc_hd__mux4_2 c197 (.A0(net130),
    .A1(net129),
    .A2(net128),
    .A3(net118),
    .S0(net116),
    .X(net709));
 sky130_fd_sc_hd__a41o_1 c198 (.A1(net20),
    .A2(net14),
    .A3(net0),
    .A4(net130),
    .B1(net1019),
    .X(net134));
 sky130_fd_sc_hd__mux4_1 c199 (.A0(net6),
    .A1(net1019),
    .A2(net889),
    .A3(net122),
    .S0(net1039),
    .S1(net85),
    .X(net135));
 sky130_fd_sc_hd__a41o_1 c200 (.A1(net909),
    .A2(net23),
    .A3(net996),
    .A4(net68),
    .B1(net708),
    .X(net136));
 sky130_fd_sc_hd__sdfbbn_1 c201 (.CLK_N(clknet_4_11_0_clk),
    .D(net134),
    .RESET_B(net20),
    .SCD(net1043),
    .SCE(net130),
    .SET_B(net878),
    .Q(net138),
    .Q_N(net137));
 sky130_fd_sc_hd__mux4_1 c202 (.A0(net121),
    .A1(net1043),
    .A2(net112),
    .A3(net21),
    .S0(net119),
    .S1(net1055),
    .X(net139));
 sky130_fd_sc_hd__a41o_2 c203 (.A1(net1036),
    .A2(net127),
    .A3(net998),
    .A4(net7),
    .B1(net130),
    .X(net140));
 sky130_fd_sc_hd__a41o_1 c204 (.A1(net138),
    .A2(net913),
    .A3(net14),
    .A4(net1031),
    .B1(net708),
    .X(net141));
 sky130_fd_sc_hd__mux4_1 c205 (.A0(net909),
    .A1(net138),
    .A2(net140),
    .A3(net996),
    .S0(net1019),
    .S1(net708),
    .X(net142));
 sky130_fd_sc_hd__a41o_1 c206 (.A1(net23),
    .A2(net121),
    .A3(net138),
    .A4(net106),
    .B1(net136),
    .X(net143));
 sky130_fd_sc_hd__mux4_1 c207 (.A0(net140),
    .A1(net119),
    .A2(net98),
    .A3(net137),
    .S0(clknet_1_0__leaf_net705),
    .S1(net1027),
    .X(net144));
 sky130_fd_sc_hd__mux4_1 c208 (.A0(net136),
    .A1(net909),
    .A2(net21),
    .A3(net20),
    .S0(clknet_1_0__leaf_net744),
    .S1(net759),
    .X(net145));
 sky130_fd_sc_hd__sdfbbn_1 c209 (.CLK_N(clknet_4_11_0_clk),
    .D(net127),
    .RESET_B(net135),
    .SCD(net913),
    .SCE(net137),
    .SET_B(net140),
    .Q(net147),
    .Q_N(net146));
 sky130_fd_sc_hd__mux4_1 c210 (.A0(net140),
    .A1(net1043),
    .A2(net6),
    .A3(net146),
    .S0(net996),
    .S1(net759),
    .X(net148));
 sky130_fd_sc_hd__a41o_2 c211 (.A1(net138),
    .A2(net146),
    .A3(net106),
    .A4(net141),
    .B1(net759),
    .X(net149));
 sky130_fd_sc_hd__mux4_1 c212 (.A0(net135),
    .A1(net130),
    .A2(net12),
    .A3(net140),
    .S0(clknet_1_0__leaf_net743),
    .S1(net759),
    .X(net150));
 sky130_fd_sc_hd__mux4_1 c213 (.A0(clknet_1_1__leaf_net145),
    .A1(net149),
    .A2(net137),
    .A3(net92),
    .S0(net122),
    .S1(net708),
    .X(net151));
 sky130_fd_sc_hd__a41o_1 c214 (.A1(net878),
    .A2(net6),
    .A3(clknet_1_0__leaf_net145),
    .A4(clknet_1_0__leaf_net705),
    .B1(clknet_1_0__leaf_net743),
    .X(net946));
 sky130_fd_sc_hd__a41o_1 c215 (.A1(net20),
    .A2(net1039),
    .A3(clknet_1_0__leaf_net946),
    .A4(net149),
    .B1(clknet_1_0__leaf_net743),
    .X(net152));
 sky130_fd_sc_hd__a41o_1 c216 (.A1(net141),
    .A2(clknet_1_0__leaf_net946),
    .A3(net7),
    .A4(net14),
    .B1(clknet_1_0__leaf_net744),
    .X(net153));
 sky130_fd_sc_hd__mux4_1 c217 (.A0(clknet_1_0__leaf_net153),
    .A1(net146),
    .A2(clknet_1_0__leaf_net946),
    .A3(clknet_1_0__leaf_net744),
    .S0(net1027),
    .S1(net759),
    .X(net154));
 sky130_fd_sc_hd__mux4_1 c218 (.A0(net80),
    .A1(clknet_1_0__leaf_net153),
    .A2(net92),
    .A3(net680),
    .S0(clknet_1_0__leaf_net743),
    .S1(net759),
    .X(net155));
 sky130_fd_sc_hd__mux4_1 c219 (.A0(net14),
    .A1(net3),
    .A2(net140),
    .A3(net137),
    .S0(net680),
    .S1(net759),
    .X(net156));
 sky130_fd_sc_hd__mux4_1 c220 (.A0(net112),
    .A1(net998),
    .A2(net140),
    .A3(clknet_1_0__leaf_net946),
    .S0(net1019),
    .S1(net961),
    .X(net157));
 sky130_fd_sc_hd__mux4_1 c221 (.A0(net996),
    .A1(net4),
    .A2(net147),
    .A3(net140),
    .S0(net112),
    .S1(clknet_1_0__leaf_net761),
    .X(net158));
 sky130_fd_sc_hd__mux4_2 c222 (.A0(net1019),
    .A1(net36),
    .A2(net913),
    .A3(net106),
    .S0(net1009),
    .S1(net666),
    .X(net926));
 sky130_fd_sc_hd__mux4_1 c223 (.A0(clknet_1_1__leaf_net153),
    .A1(net35),
    .A2(net961),
    .A3(net755),
    .S0(net966),
    .S1(clknet_1_1__leaf_net761),
    .X(net159));
 sky130_fd_sc_hd__mux4_1 c224 (.A0(net969),
    .A1(net1056),
    .A2(clknet_1_1__leaf_net153),
    .A3(net666),
    .S0(net681),
    .S1(net764),
    .X(net160));
 sky130_fd_sc_hd__mux4_1 c225 (.A0(net147),
    .A1(net926),
    .A2(clknet_1_1__leaf_net705),
    .A3(net966),
    .S0(clknet_1_1__leaf_net762),
    .S1(net765),
    .X(net161));
 sky130_fd_sc_hd__mux4_1 c226 (.A0(net926),
    .A1(net30),
    .A2(net998),
    .A3(net1070),
    .S0(net756),
    .S1(clknet_1_0__leaf_net761),
    .X(net162));
 sky130_fd_sc_hd__mux4_1 c227 (.A0(net92),
    .A1(net1039),
    .A2(net926),
    .A3(net681),
    .S0(clknet_1_1__leaf_net762),
    .S1(net765),
    .X(net163));
 sky130_fd_sc_hd__mux4_1 c228 (.A0(net106),
    .A1(net92),
    .A2(clknet_1_1__leaf_net153),
    .A3(net1019),
    .S0(clknet_1_1__leaf_net760),
    .S1(net766),
    .X(net164));
 sky130_fd_sc_hd__mux4_1 c229 (.A0(net140),
    .A1(net908),
    .A2(net926),
    .A3(clknet_1_1__leaf_net762),
    .S0(net765),
    .S1(net766),
    .X(net165));
 sky130_fd_sc_hd__mux4_1 c230 (.A0(net1056),
    .A1(net1009),
    .A2(clknet_1_1__leaf_net153),
    .A3(clknet_1_0__leaf_net761),
    .S0(net767),
    .S1(net768),
    .X(net166));
 sky130_fd_sc_hd__mux4_1 c231 (.A0(net1043),
    .A1(net1055),
    .A2(clknet_1_1__leaf_net153),
    .A3(net1009),
    .S0(net763),
    .S1(net770),
    .X(net167));
 sky130_fd_sc_hd__mux4_1 c232 (.A0(net913),
    .A1(net996),
    .A2(net85),
    .A3(net112),
    .S0(net764),
    .S1(net767),
    .X(net168));
 sky130_fd_sc_hd__mux4_1 c233 (.A0(net147),
    .A1(clknet_1_1__leaf_net744),
    .A2(clknet_1_1__leaf_net762),
    .A3(net929),
    .S0(net768),
    .S1(net769),
    .X(net972));
 sky130_fd_sc_hd__mux4_2 c234 (.A0(net147),
    .A1(net90),
    .A2(net1038),
    .A3(net966),
    .S0(net763),
    .S1(net770),
    .X(net169));
 sky130_fd_sc_hd__mux4_1 c235 (.A0(net4),
    .A1(net140),
    .A2(net961),
    .A3(net767),
    .S0(net769),
    .S1(net770),
    .X(net170));
 sky130_fd_sc_hd__mux4_1 c236 (.A0(net40),
    .A1(net1035),
    .A2(clknet_1_0__leaf_net761),
    .A3(net764),
    .S0(net769),
    .S1(net770),
    .X(net171));
 sky130_fd_sc_hd__mux4_1 c237 (.A0(net30),
    .A1(net38),
    .A2(net168),
    .A3(net763),
    .S0(net766),
    .S1(net771),
    .X(net172));
 sky130_fd_sc_hd__mux4_1 c238 (.A0(net85),
    .A1(clknet_1_0__leaf_net171),
    .A2(net172),
    .A3(net169),
    .S0(net961),
    .S1(net771),
    .X(net173));
 sky130_fd_sc_hd__mux4_2 c239 (.A0(net169),
    .A1(net765),
    .A2(net767),
    .A3(net769),
    .S0(net771),
    .S1(net772),
    .X(net174));
 sky130_fd_sc_hd__mux4_1 c240 (.A0(net168),
    .A1(net174),
    .A2(net998),
    .A3(net960),
    .S0(net929),
    .S1(net772),
    .X(net175));
 sky130_fd_sc_hd__mux4_1 c241 (.A0(clknet_1_1__leaf_net171),
    .A1(net85),
    .A2(net169),
    .A3(net175),
    .S0(net766),
    .S1(net769),
    .X(net957));
 sky130_fd_sc_hd__mux4_1 c242 (.A0(clknet_1_0__leaf_net67),
    .A1(net65),
    .A2(clknet_1_0__leaf_net62),
    .A3(net97),
    .S0(net1055),
    .S1(net765),
    .X(net176));
 sky130_fd_sc_hd__mux4_1 c243 (.A0(net69),
    .A1(net1044),
    .A2(clknet_1_0__leaf_net959),
    .A3(net1040),
    .S0(net943),
    .S1(net1027),
    .X(net177));
 sky130_fd_sc_hd__mux4_1 c244 (.A0(clknet_1_0__leaf_net177),
    .A1(net926),
    .A2(clknet_1_0__leaf_net62),
    .A3(net969),
    .S0(clknet_1_0__leaf_net744),
    .S1(net755),
    .X(net178));
 sky130_fd_sc_hd__mux4_1 c245 (.A0(clknet_1_0__leaf_net177),
    .A1(net97),
    .A2(net51),
    .A3(clknet_1_1__leaf_net744),
    .S0(net1027),
    .S1(net966),
    .X(net179));
 sky130_fd_sc_hd__mux4_1 c246 (.A0(clknet_1_0__leaf_net179),
    .A1(net46),
    .A2(clknet_1_0__leaf_net959),
    .A3(net1045),
    .S0(clknet_1_1__leaf_net177),
    .S1(net966),
    .X(net937));
 sky130_fd_sc_hd__mux4_1 c247 (.A0(net65),
    .A1(clknet_1_0__leaf_net177),
    .A2(net967),
    .A3(net960),
    .S0(net966),
    .S1(clknet_1_0__leaf_net761),
    .X(net180));
 sky130_fd_sc_hd__mux4_1 c248 (.A0(net36),
    .A1(clknet_1_0__leaf_net177),
    .A2(clknet_1_1__leaf_net179),
    .A3(net732),
    .S0(net749),
    .S1(clknet_1_1__leaf_net761),
    .X(net181));
 sky130_fd_sc_hd__mux4_1 c249 (.A0(net46),
    .A1(clknet_1_0__leaf_net62),
    .A2(net1040),
    .A3(net732),
    .S0(net749),
    .S1(net929),
    .X(net182));
 sky130_fd_sc_hd__mux4_1 c250 (.A0(clknet_1_1__leaf_net181),
    .A1(clknet_1_1__leaf_net177),
    .A2(clknet_1_0__leaf_net182),
    .A3(net51),
    .S0(net926),
    .S1(clknet_1_0__leaf_net959),
    .X(net183));
 sky130_fd_sc_hd__mux4_1 c251 (.A0(clknet_1_0__leaf_net49),
    .A1(net1041),
    .A2(clknet_1_0__leaf_net182),
    .A3(clknet_1_1__leaf_net177),
    .S0(clknet_1_0__leaf_net181),
    .S1(net963),
    .X(net971));
 sky130_fd_sc_hd__mux4_1 c252 (.A0(net175),
    .A1(net1045),
    .A2(clknet_1_1__leaf_net177),
    .A3(clknet_1_0__leaf_net959),
    .S0(clknet_1_0__leaf_net182),
    .S1(net732),
    .X(net184));
 sky130_fd_sc_hd__mux4_1 c253 (.A0(net1044),
    .A1(net69),
    .A2(clknet_1_0__leaf_net182),
    .A3(clknet_1_0__leaf_net177),
    .S0(net65),
    .S1(net749),
    .X(net185));
 sky130_fd_sc_hd__mux4_1 c254 (.A0(clknet_1_1__leaf_net62),
    .A1(clknet_1_1__leaf_net182),
    .A2(net51),
    .A3(clknet_1_1__leaf_net177),
    .S0(clknet_1_0__leaf_net185),
    .S1(net956),
    .X(net186));
 sky130_fd_sc_hd__mux4_1 c255 (.A0(clknet_1_1__leaf_net67),
    .A1(net35),
    .A2(clknet_1_0__leaf_net184),
    .A3(net949),
    .S0(clknet_1_1__leaf_net761),
    .S1(net773),
    .X(net187));
 sky130_fd_sc_hd__mux4_1 c256 (.A0(clknet_1_0__leaf_net182),
    .A1(net1045),
    .A2(net749),
    .A3(net929),
    .S0(net956),
    .S1(net775),
    .X(net188));
 sky130_fd_sc_hd__mux4_1 c257 (.A0(clknet_1_1__leaf_net188),
    .A1(clknet_1_1__leaf_net182),
    .A2(net64),
    .A3(net756),
    .S0(net773),
    .S1(net775),
    .X(net189));
 sky130_fd_sc_hd__mux4_1 c258 (.A0(clknet_1_1__leaf_net184),
    .A1(clknet_1_1__leaf_net62),
    .A2(clknet_1_1__leaf_net744),
    .A3(net966),
    .S0(net956),
    .S1(net775),
    .X(net190));
 sky130_fd_sc_hd__mux4_1 c259 (.A0(net949),
    .A1(clknet_1_1__leaf_net761),
    .A2(net765),
    .A3(net956),
    .S0(net775),
    .S1(net776),
    .X(net191));
 sky130_fd_sc_hd__mux4_1 c260 (.A0(clknet_1_0__leaf_net191),
    .A1(clknet_1_1__leaf_net182),
    .A2(net51),
    .A3(net773),
    .S0(net774),
    .S1(net776),
    .X(net192));
 sky130_fd_sc_hd__mux4_1 c261 (.A0(net192),
    .A1(clknet_1_1__leaf_net191),
    .A2(net949),
    .A3(net773),
    .S0(net774),
    .S1(net776),
    .X(net193));
 sky130_fd_sc_hd__mux4_1 c262 (.A0(clknet_1_1__leaf_net182),
    .A1(clknet_1_1__leaf_net62),
    .A2(net949),
    .A3(clknet_1_1__leaf_net743),
    .S0(net774),
    .S1(net776),
    .X(net194));
 sky130_fd_sc_hd__mux4_1 c263 (.A0(clknet_1_1__leaf_net185),
    .A1(net194),
    .A2(clknet_1_1__leaf_net62),
    .A3(clknet_1_1__leaf_net743),
    .S0(net774),
    .S1(net776),
    .X(net195));
 sky130_fd_sc_hd__xnor2_1 c264 (.A(net1002),
    .B(net1071),
    .Y(net196));
 sky130_fd_sc_hd__a41o_4 c265 (.A1(net86),
    .A2(net866),
    .A3(net1020),
    .A4(net1058),
    .B1(net999),
    .X(net197));
 sky130_fd_sc_hd__xnor2_2 c266 (.A(net1066),
    .B(net197),
    .Y(net198));
 sky130_fd_sc_hd__a21bo_1 c267 (.A1(net89),
    .A2(net198),
    .B1_N(net1001),
    .X(net199));
 sky130_fd_sc_hd__a21bo_2 c268 (.A1(net197),
    .A2(net83),
    .B1_N(net1066),
    .X(net200));
 sky130_fd_sc_hd__a21bo_1 c269 (.A1(net199),
    .A2(net866),
    .B1_N(net200),
    .X(net201));
 sky130_fd_sc_hd__a31o_2 c270 (.A1(net199),
    .A2(net200),
    .A3(net999),
    .B1(net83),
    .X(net202));
 sky130_fd_sc_hd__a21bo_1 c271 (.A1(net200),
    .A2(net202),
    .B1_N(net198),
    .X(net203));
 sky130_fd_sc_hd__a21bo_1 c272 (.A1(net198),
    .A2(net201),
    .B1_N(net202),
    .X(net204));
 sky130_fd_sc_hd__xnor2_2 c273 (.A(net990),
    .B(net989),
    .Y(net205));
 sky130_fd_sc_hd__a21bo_1 c274 (.A1(net205),
    .A2(net999),
    .B1_N(net989),
    .X(net206));
 sky130_fd_sc_hd__a21bo_1 c275 (.A1(net205),
    .A2(net199),
    .B1_N(net989),
    .X(net207));
 sky130_fd_sc_hd__mux4_2 c276 (.A0(net71),
    .A1(net206),
    .A2(net205),
    .A3(net999),
    .S0(net1066),
    .S1(net1071),
    .X(net208));
 sky130_fd_sc_hd__mux4_2 c277 (.A0(net79),
    .A1(net207),
    .A2(net201),
    .A3(net205),
    .S0(net199),
    .S1(net1046),
    .X(net209));
 sky130_fd_sc_hd__mux4_1 c278 (.A0(net208),
    .A1(net999),
    .A2(net202),
    .A3(net989),
    .S0(net980),
    .S1(net1066),
    .X(net210));
 sky130_fd_sc_hd__a31o_1 c279 (.A1(net201),
    .A2(net199),
    .A3(net207),
    .B1(net668),
    .X(net211));
 sky130_fd_sc_hd__sdfrbp_2 c280 (.CLK(clknet_4_2_0_clk),
    .D(net211),
    .RESET_B(net205),
    .SCD(net990),
    .SCE(net668),
    .Q(net213),
    .Q_N(net212));
 sky130_fd_sc_hd__sdfbbp_1 c281 (.CLK(clknet_4_2_0_clk),
    .D(net207),
    .RESET_B(net200),
    .SCD(net211),
    .SCE(net866),
    .SET_B(net989),
    .Q(net215),
    .Q_N(net214));
 sky130_fd_sc_hd__a41o_1 c282 (.A1(net198),
    .A2(net206),
    .A3(net212),
    .A4(net208),
    .B1(net668),
    .X(net216));
 sky130_fd_sc_hd__mux4_2 c283 (.A0(net213),
    .A1(net75),
    .A2(net206),
    .A3(net198),
    .S0(net999),
    .S1(net674),
    .X(net217));
 sky130_fd_sc_hd__a41o_1 c284 (.A1(net217),
    .A2(net989),
    .A3(net75),
    .A4(net214),
    .B1(net674),
    .X(net218));
 sky130_fd_sc_hd__mux4_1 c285 (.A0(net989),
    .A1(net206),
    .A2(net217),
    .A3(net208),
    .S0(net668),
    .S1(net674),
    .X(net219));
 sky130_fd_sc_hd__a31o_1 c286 (.A1(net876),
    .A2(net1063),
    .A3(net889),
    .B1(net777),
    .X(net220));
 sky130_fd_sc_hd__a21bo_2 c287 (.A1(net1063),
    .A2(net1001),
    .B1_N(net95),
    .X(net221));
 sky130_fd_sc_hd__a21bo_2 c288 (.A1(net96),
    .A2(net1007),
    .B1_N(net1031),
    .X(net222));
 sky130_fd_sc_hd__a31o_1 c289 (.A1(net206),
    .A2(net95),
    .A3(net196),
    .B1(net1058),
    .X(net223));
 sky130_fd_sc_hd__a31o_1 c290 (.A1(net220),
    .A2(net1063),
    .A3(net880),
    .B1(net81),
    .X(net224));
 sky130_fd_sc_hd__a21bo_1 c291 (.A1(net96),
    .A2(net84),
    .B1_N(net222),
    .X(net225));
 sky130_fd_sc_hd__mux4_1 c292 (.A0(net225),
    .A1(net223),
    .A2(net222),
    .A3(net980),
    .S0(net78),
    .S1(net96),
    .X(net226));
 sky130_fd_sc_hd__mux4_1 c293 (.A0(net224),
    .A1(net222),
    .A2(net223),
    .A3(net876),
    .S0(net1031),
    .S1(net777),
    .X(net227));
 sky130_fd_sc_hd__a21bo_4 c294 (.A1(net225),
    .A2(net674),
    .B1_N(net1026),
    .X(net228));
 sky130_fd_sc_hd__a21bo_1 c295 (.A1(net657),
    .A2(net668),
    .B1_N(net1026),
    .X(net229));
 sky130_fd_sc_hd__a31o_1 c296 (.A1(net892),
    .A2(net221),
    .A3(net202),
    .B1(net98),
    .X(net230));
 sky130_fd_sc_hd__a21bo_1 c297 (.A1(net224),
    .A2(net230),
    .B1_N(net668),
    .X(net231));
 sky130_fd_sc_hd__mux4_2 c298 (.A0(net230),
    .A1(net224),
    .A2(net889),
    .A3(net990),
    .S0(net880),
    .S1(net1026),
    .X(net232));
 sky130_fd_sc_hd__mux4_1 c299 (.A0(net223),
    .A1(net98),
    .A2(net232),
    .A3(net222),
    .S1(net757),
    .X(net233));
 sky130_fd_sc_hd__a21bo_1 c300 (.A1(net1007),
    .A2(net228),
    .B1_N(net668),
    .X(net234));
 sky130_fd_sc_hd__a21bo_2 c301 (.A1(net232),
    .A2(net657),
    .B1_N(net1031),
    .X(net975));
 sky130_fd_sc_hd__mux4_1 c302 (.A0(net887),
    .A1(net232),
    .A2(net975),
    .A3(net894),
    .S0(net96),
    .S1(net657),
    .X(net235));
 sky130_fd_sc_hd__mux4_1 c303 (.A0(net89),
    .A1(net223),
    .A2(net1005),
    .A3(net1045),
    .S0(net1050),
    .S1(clknet_1_1__leaf_net778),
    .X(net236));
 sky130_fd_sc_hd__mux4_2 c304 (.A0(net221),
    .A1(net96),
    .A2(net657),
    .A3(net668),
    .S0(net674),
    .S1(net1031),
    .X(net237));
 sky130_fd_sc_hd__mux4_1 c305 (.A0(net234),
    .A1(net96),
    .A2(net228),
    .A3(net673),
    .S0(net1031),
    .S1(clknet_1_1__leaf_net778),
    .X(net238));
 sky130_fd_sc_hd__mux4_1 c306 (.A0(net234),
    .A1(net896),
    .A2(net96),
    .A3(net223),
    .S0(net232),
    .S1(net673),
    .X(net239));
 sky130_fd_sc_hd__mux4_2 c307 (.A0(net229),
    .A1(net224),
    .A2(net202),
    .A3(net232),
    .S0(net230),
    .S1(net673),
    .X(net240));
 sky130_fd_sc_hd__buf_2 c308 (.A(net738),
    .X(net950));
 sky130_fd_sc_hd__a21bo_1 c309 (.A1(net117),
    .A2(net221),
    .B1_N(net1027),
    .X(net241));
 sky130_fd_sc_hd__a41o_1 c310 (.A1(net241),
    .A2(net897),
    .A3(net644),
    .A4(net657),
    .B1(net709),
    .X(net242));
 sky130_fd_sc_hd__clkbuf_1 c311 (.A(net738),
    .X(net243));
 sky130_fd_sc_hd__mux4_1 c312 (.A0(net84),
    .A1(net241),
    .A2(net950),
    .A3(net1065),
    .S0(net975),
    .S1(net709),
    .X(net244));
 sky130_fd_sc_hd__a41o_1 c313 (.A1(net221),
    .A2(net908),
    .A3(net76),
    .A4(net644),
    .B1(clknet_1_0__leaf_net780),
    .X(net245));
 sky130_fd_sc_hd__a41o_1 c314 (.A1(net129),
    .A2(clknet_1_0__leaf_net245),
    .A3(net99),
    .A4(clknet_1_1__leaf_net778),
    .B1(clknet_1_0__leaf_net780),
    .X(net246));
 sky130_fd_sc_hd__buf_1 c315 (.A(net672),
    .X(net247));
 sky130_fd_sc_hd__mux4_1 c316 (.A0(net897),
    .A1(clknet_1_0__leaf_net245),
    .A2(net117),
    .A3(clknet_1_1__leaf_net246),
    .S0(net131),
    .S1(net95),
    .X(net248));
 sky130_fd_sc_hd__buf_1 c317 (.A(net672),
    .X(net249));
 sky130_fd_sc_hd__mux4_1 c318 (.A0(net95),
    .A1(net950),
    .A2(net673),
    .A3(net757),
    .S0(clknet_1_0__leaf_net779),
    .S1(net782),
    .X(net250));
 sky130_fd_sc_hd__mux4_1 c319 (.A0(net241),
    .A1(net0),
    .A2(net129),
    .A3(net1036),
    .S0(net758),
    .S1(clknet_1_0__leaf_net780),
    .X(net251));
 sky130_fd_sc_hd__mux4_1 c320 (.A0(net240),
    .A1(net124),
    .A2(clknet_1_1__leaf_net251),
    .A3(net1038),
    .S0(clknet_1_0__leaf_net245),
    .S1(net777),
    .X(net252));
 sky130_fd_sc_hd__mux4_1 c321 (.A0(net889),
    .A1(net247),
    .A2(clknet_1_0__leaf_net250),
    .A3(clknet_1_0__leaf_net251),
    .S0(net673),
    .S1(net709),
    .X(net253));
 sky130_fd_sc_hd__sdfbbn_1 c322 (.CLK_N(clknet_4_8_0_clk),
    .D(clknet_1_0__leaf_net253),
    .RESET_B(clknet_1_1__leaf_net246),
    .SCD(net249),
    .SCE(net1061),
    .SET_B(net1028),
    .Q(net255),
    .Q_N(net254));
 sky130_fd_sc_hd__mux4_1 c323 (.A0(net118),
    .A1(net255),
    .A2(net241),
    .A3(clknet_1_0__leaf_net251),
    .S0(net885),
    .S1(net215),
    .X(net256));
 sky130_fd_sc_hd__mux4_1 c324 (.A0(net99),
    .A1(net255),
    .A2(clknet_1_0__leaf_net251),
    .A3(net242),
    .S0(net1038),
    .S1(net1031),
    .X(net257));
 sky130_fd_sc_hd__a41o_1 c325 (.A1(net240),
    .A2(net255),
    .A3(net980),
    .A4(net1028),
    .B1(net777),
    .X(net258));
 sky130_fd_sc_hd__mux4_1 c326 (.A0(clknet_1_1__leaf_net253),
    .A1(net254),
    .A2(net0),
    .A3(net734),
    .S0(clknet_1_0__leaf_net780),
    .S1(net782),
    .X(net259));
 sky130_fd_sc_hd__mux4_1 c327 (.A0(net131),
    .A1(net255),
    .A2(net129),
    .A3(clknet_1_0__leaf_net251),
    .S0(clknet_1_1__leaf_net257),
    .S1(net976),
    .X(net260));
 sky130_fd_sc_hd__a41o_1 c328 (.A1(clknet_1_1__leaf_net246),
    .A2(net882),
    .A3(net128),
    .A4(net254),
    .B1(net1028),
    .X(net261));
 sky130_fd_sc_hd__mux4_1 c329 (.A0(net261),
    .A1(net128),
    .A2(net254),
    .A3(net657),
    .S0(net1028),
    .S1(net783),
    .X(net262));
 sky130_fd_sc_hd__mux4_1 c330 (.A0(net221),
    .A1(net7),
    .A2(clknet_1_0__leaf_net153),
    .A3(net98),
    .S0(clknet_1_0__leaf_net760),
    .S1(net777),
    .X(net263));
 sky130_fd_sc_hd__mux4_1 c331 (.A0(clknet_1_1__leaf_net251),
    .A1(net249),
    .A2(net149),
    .A3(clknet_1_0__leaf_net760),
    .S0(clknet_1_0__leaf_net779),
    .S1(net782),
    .X(net264));
 sky130_fd_sc_hd__mux4_1 c332 (.A0(net21),
    .A1(clknet_1_1__leaf_net251),
    .A2(net149),
    .A3(net138),
    .S0(net980),
    .S1(net786),
    .X(net265));
 sky130_fd_sc_hd__mux4_1 c333 (.A0(net149),
    .A1(net119),
    .A2(net221),
    .A3(net124),
    .S1(net781),
    .X(net266));
 sky130_fd_sc_hd__mux4_1 c334 (.A0(net896),
    .A1(net1019),
    .A2(net137),
    .A3(clknet_1_0__leaf_net153),
    .S0(net966),
    .S1(clknet_1_1__leaf_net780),
    .X(net267));
 sky130_fd_sc_hd__mux4_1 c335 (.A0(net128),
    .A1(net130),
    .A2(clknet_1_0__leaf_net153),
    .A3(net237),
    .S0(net966),
    .S1(net1024),
    .X(net268));
 sky130_fd_sc_hd__mux4_1 c336 (.A0(net0),
    .A1(net149),
    .A2(net21),
    .A3(net1055),
    .S0(net781),
    .S1(net1024),
    .X(net269));
 sky130_fd_sc_hd__mux4_1 c337 (.A0(net12),
    .A1(net18),
    .A2(net1040),
    .A3(net149),
    .S0(net746),
    .S1(net777),
    .X(net270));
 sky130_fd_sc_hd__mux4_1 c338 (.A0(net3),
    .A1(net975),
    .A2(net989),
    .A3(net1088),
    .S0(net786),
    .S1(net1076),
    .X(net271));
 sky130_fd_sc_hd__a41o_1 c339 (.A1(net130),
    .A2(net221),
    .A3(net740),
    .A4(net1025),
    .B1(net789),
    .X(net272));
 sky130_fd_sc_hd__mux4_1 c340 (.A0(clknet_1_0__leaf_net250),
    .A1(clknet_1_0__leaf_net760),
    .A2(clknet_1_1__leaf_net780),
    .A3(net784),
    .S0(net1025),
    .S1(net790),
    .X(net273));
 sky130_fd_sc_hd__mux4_1 c341 (.A0(net272),
    .A1(clknet_1_1__leaf_net250),
    .A2(net21),
    .A3(net661),
    .S0(net746),
    .S1(clknet_1_0__leaf_net779),
    .X(net274));
 sky130_fd_sc_hd__mux4_1 c342 (.A0(clknet_1_0__leaf_net273),
    .A1(net130),
    .A2(net247),
    .A3(net661),
    .S0(net781),
    .S1(net785),
    .X(net275));
 sky130_fd_sc_hd__mux4_1 c343 (.A0(net7),
    .A1(net149),
    .A2(net662),
    .A3(net777),
    .S0(net786),
    .S1(net790),
    .X(net276));
 sky130_fd_sc_hd__mux4_1 c344 (.A0(clknet_1_1__leaf_net273),
    .A1(net975),
    .A2(net1003),
    .A3(clknet_1_0__leaf_net275),
    .S0(net746),
    .S1(net970),
    .X(net277));
 sky130_fd_sc_hd__mux4_1 c345 (.A0(clknet_1_0__leaf_net273),
    .A1(clknet_1_0__leaf_net153),
    .A2(net882),
    .A3(net1051),
    .S0(net1025),
    .S1(net794),
    .X(net278));
 sky130_fd_sc_hd__mux4_1 c346 (.A0(net272),
    .A1(net119),
    .A2(net733),
    .A3(net739),
    .S0(clknet_1_1__leaf_net780),
    .S1(net794),
    .X(net279));
 sky130_fd_sc_hd__mux4_1 c347 (.A0(clknet_1_1__leaf_net245),
    .A1(net272),
    .A2(net7),
    .A3(net1018),
    .S0(net1028),
    .S1(net970),
    .X(net280));
 sky130_fd_sc_hd__mux4_2 c348 (.A0(net727),
    .A1(net733),
    .A2(net790),
    .A3(net791),
    .S0(net794),
    .S1(net795),
    .X(net281));
 sky130_fd_sc_hd__mux4_1 c349 (.A0(clknet_1_1__leaf_net946),
    .A1(net733),
    .A2(net739),
    .A3(net786),
    .S0(net1025),
    .S1(net795),
    .X(net282));
 sky130_fd_sc_hd__mux4_1 c350 (.A0(clknet_1_0__leaf_net282),
    .A1(net12),
    .A2(net281),
    .A3(net727),
    .S0(net787),
    .S1(net794),
    .X(net283));
 sky130_fd_sc_hd__mux4_2 c351 (.A0(net281),
    .A1(net4),
    .A2(net662),
    .A3(net727),
    .S0(net733),
    .S1(net795),
    .X(net284));
 sky130_fd_sc_hd__mux4_1 c352 (.A0(net4),
    .A1(net1059),
    .A2(net119),
    .A3(net40),
    .S0(net865),
    .S1(net1003),
    .X(net285));
 sky130_fd_sc_hd__mux4_1 c353 (.A0(clknet_1_0__leaf_net275),
    .A1(net1019),
    .A2(net740),
    .A3(clknet_1_1__leaf_net760),
    .S0(net765),
    .S1(net769),
    .X(net286));
 sky130_fd_sc_hd__mux4_1 c354 (.A0(net98),
    .A1(clknet_1_0__leaf_net282),
    .A2(clknet_1_1__leaf_net760),
    .A3(net782),
    .S0(net1025),
    .S1(net791),
    .X(net287));
 sky130_fd_sc_hd__sdfbbn_1 c355 (.CLK_N(clknet_4_13_0_clk),
    .D(net967),
    .RESET_B(net740),
    .SCD(net1086),
    .SCE(net772),
    .SET_B(net1078),
    .Q(net289),
    .Q_N(net288));
 sky130_fd_sc_hd__mux4_2 c356 (.A0(net40),
    .A1(net908),
    .A2(net963),
    .A3(net771),
    .S0(net782),
    .S1(net786),
    .X(net930));
 sky130_fd_sc_hd__mux4_1 c357 (.A0(clknet_1_1__leaf_net282),
    .A1(net980),
    .A2(net1018),
    .A3(net1008),
    .S0(net772),
    .S1(net796),
    .X(net290));
 sky130_fd_sc_hd__mux4_1 c358 (.A0(net285),
    .A1(net1002),
    .A2(clknet_1_1__leaf_net282),
    .A3(net765),
    .S0(net770),
    .S1(net791),
    .X(net291));
 sky130_fd_sc_hd__mux4_2 c359 (.A0(net289),
    .A1(net930),
    .A2(net725),
    .A3(net740),
    .S0(net768),
    .S1(net786),
    .X(net940));
 sky130_fd_sc_hd__mux4_2 c360 (.A0(net247),
    .A1(net213),
    .A2(net1019),
    .A3(net288),
    .S0(net745),
    .S1(net765),
    .X(net292));
 sky130_fd_sc_hd__a41o_1 c361 (.A1(net292),
    .A2(clknet_1_1__leaf_net275),
    .A3(net1046),
    .A4(net40),
    .B1(net998),
    .X(net293));
 sky130_fd_sc_hd__a41o_1 c362 (.A1(net289),
    .A2(net292),
    .A3(net940),
    .A4(net284),
    .B1(clknet_1_1__leaf_net282),
    .X(net294));
 sky130_fd_sc_hd__sdfbbp_1 c363 (.CLK(clknet_4_13_0_clk),
    .D(clknet_1_1__leaf_net153),
    .RESET_B(clknet_1_0__leaf_net957),
    .SCD(net975),
    .SCE(net962),
    .SET_B(clknet_1_1__leaf_net779),
    .Q(net296),
    .Q_N(net295));
 sky130_fd_sc_hd__mux4_1 c364 (.A0(net292),
    .A1(clknet_1_0__leaf_net705),
    .A2(net961),
    .A3(net745),
    .S0(net772),
    .S1(net787),
    .X(net297));
 sky130_fd_sc_hd__mux4_1 c365 (.A0(net1008),
    .A1(net930),
    .A2(clknet_1_1__leaf_net153),
    .A3(net668),
    .S0(net745),
    .S1(clknet_1_1__leaf_net762),
    .X(net298));
 sky130_fd_sc_hd__mux4_1 c366 (.A0(net172),
    .A1(net1038),
    .A2(net1010),
    .A3(clknet_1_0__leaf_net946),
    .S0(net288),
    .S1(net961),
    .X(net299));
 sky130_fd_sc_hd__mux4_2 c367 (.A0(net174),
    .A1(net296),
    .A2(net284),
    .A3(net1008),
    .S0(net734),
    .S1(clknet_1_1__leaf_net797),
    .X(net300));
 sky130_fd_sc_hd__mux4_2 c368 (.A0(net1000),
    .A1(net1040),
    .A2(net4),
    .A3(net212),
    .S0(clknet_1_1__leaf_net300),
    .S1(clknet_1_1__leaf_net797),
    .X(net947));
 sky130_fd_sc_hd__mux4_1 c369 (.A0(net872),
    .A1(clknet_1_1__leaf_net153),
    .A2(clknet_1_1__leaf_net300),
    .A3(net292),
    .S0(net745),
    .S1(net796),
    .X(net301));
 sky130_fd_sc_hd__mux4_1 c370 (.A0(net297),
    .A1(net292),
    .A2(net1008),
    .A3(net961),
    .S0(net772),
    .S1(clknet_1_0__leaf_net797),
    .X(net302));
 sky130_fd_sc_hd__mux4_1 c371 (.A0(net296),
    .A1(clknet_1_1__leaf_net302),
    .A2(net734),
    .A3(net768),
    .S0(net781),
    .S1(clknet_1_1__leaf_net798),
    .X(net303));
 sky130_fd_sc_hd__mux4_1 c372 (.A0(clknet_1_1__leaf_net275),
    .A1(net1003),
    .A2(clknet_1_1__leaf_net303),
    .A3(net1036),
    .S0(clknet_1_0__leaf_net946),
    .S1(clknet_1_0__leaf_net797),
    .X(net304));
 sky130_fd_sc_hd__mux4_1 c373 (.A0(net295),
    .A1(clknet_1_0__leaf_net947),
    .A2(clknet_1_1__leaf_net705),
    .A3(net725),
    .S0(net796),
    .S1(clknet_1_1__leaf_net797),
    .X(net964));
 sky130_fd_sc_hd__mux4_1 c392 (.A0(net942),
    .A1(clknet_1_0__leaf_net972),
    .A2(clknet_1_0__leaf_net965),
    .A3(clknet_1_0__leaf_net971),
    .S0(net960),
    .S1(clknet_1_1__leaf_net779),
    .X(net305));
 sky130_fd_sc_hd__mux4_1 c393 (.A0(net36),
    .A1(net215),
    .A2(clknet_1_0__leaf_net959),
    .A3(net968),
    .S0(net702),
    .S1(net963),
    .X(net974));
 sky130_fd_sc_hd__mux4_1 c394 (.A0(clknet_1_0__leaf_net188),
    .A1(clknet_1_0__leaf_net974),
    .A2(clknet_1_0__leaf_net937),
    .S0(net702),
    .S1(clknet_1_1__leaf_net779),
    .X(net306));
 sky130_fd_sc_hd__a41o_1 c395 (.A1(net17),
    .A2(clknet_1_0__leaf_net974),
    .A3(net968),
    .A4(net702),
    .B1(clknet_1_1__leaf_net779),
    .X(net941));
 sky130_fd_sc_hd__xnor2_1 c396 (.A(net197),
    .B(net1035),
    .Y(net307));
 sky130_fd_sc_hd__buf_1 c397 (.A(net675),
    .X(net308));
 sky130_fd_sc_hd__buf_1 c398 (.A(net675),
    .X(net309));
 sky130_fd_sc_hd__a21bo_2 c399 (.A1(net309),
    .A2(net197),
    .B1_N(net1007),
    .X(net310));
 sky130_fd_sc_hd__xnor2_2 c400 (.A(net995),
    .B(net999),
    .Y(net311));
 sky130_fd_sc_hd__a21bo_4 c401 (.A1(net73),
    .A2(net866),
    .B1_N(net311),
    .X(net312));
 sky130_fd_sc_hd__a41o_1 c402 (.A1(net994),
    .A2(net1054),
    .A3(net211),
    .A4(net1065),
    .B1(net990),
    .X(net313));
 sky130_fd_sc_hd__mux4_1 c403 (.A0(net75),
    .A1(net88),
    .A2(net1063),
    .A3(net77),
    .S0(net309),
    .S1(net866),
    .X(net314));
 sky130_fd_sc_hd__a31o_4 c404 (.A1(net307),
    .A2(net994),
    .A3(net314),
    .B1(net202),
    .X(net315));
 sky130_fd_sc_hd__a21bo_1 c405 (.A1(net314),
    .A2(net307),
    .B1_N(net214),
    .X(net316));
 sky130_fd_sc_hd__a21bo_2 c406 (.A1(net82),
    .A2(net311),
    .B1_N(net312),
    .X(net317));
 sky130_fd_sc_hd__a21bo_1 c407 (.A1(net317),
    .A2(net308),
    .B1_N(net1047),
    .X(net318));
 sky130_fd_sc_hd__a31o_1 c408 (.A1(net314),
    .A2(net211),
    .A3(net317),
    .B1(net986),
    .X(net319));
 sky130_fd_sc_hd__a21bo_1 c409 (.A1(net986),
    .A2(net315),
    .B1_N(net649),
    .X(net320));
 sky130_fd_sc_hd__a41o_4 c410 (.A1(net316),
    .A2(net986),
    .A3(net1001),
    .A4(net317),
    .B1(net714),
    .X(net321));
 sky130_fd_sc_hd__a41o_1 c411 (.A1(net311),
    .A2(net1033),
    .A3(net321),
    .A4(net982),
    .B1(net866),
    .X(net322));
 sky130_fd_sc_hd__mux4_1 c412 (.A0(net989),
    .A1(net322),
    .A2(net987),
    .A3(net315),
    .S0(net994),
    .S1(net982),
    .X(net323));
 sky130_fd_sc_hd__a41o_1 c413 (.A1(net315),
    .A2(net321),
    .A3(net995),
    .A4(net994),
    .B1(net1074),
    .X(net324));
 sky130_fd_sc_hd__mux4_1 c414 (.A0(net866),
    .A1(net324),
    .A2(net987),
    .A3(net995),
    .S0(net312),
    .S1(net649),
    .X(net325));
 sky130_fd_sc_hd__mux4_1 c415 (.A0(net322),
    .A1(net197),
    .A2(net312),
    .A3(net982),
    .S0(net316),
    .S1(net714),
    .X(net326));
 sky130_fd_sc_hd__mux4_1 c416 (.A0(net317),
    .A1(net324),
    .A2(net987),
    .A3(net989),
    .S0(net982),
    .S1(net648),
    .X(net327));
 sky130_fd_sc_hd__mux4_2 c417 (.A0(net312),
    .A1(net1007),
    .A2(net987),
    .A3(net714),
    .S0(net800),
    .S1(net803),
    .X(net328));
 sky130_fd_sc_hd__a21bo_2 c418 (.A1(net315),
    .A2(net200),
    .B1_N(net803),
    .X(net329));
 sky130_fd_sc_hd__a21bo_1 c419 (.A1(net232),
    .A2(clknet_1_1__leaf_net778),
    .B1_N(clknet_1_0__leaf_net799),
    .X(net330));
 sky130_fd_sc_hd__a21bo_1 c420 (.A1(clknet_1_0__leaf_net238),
    .A2(net317),
    .B1_N(net232),
    .X(net331));
 sky130_fd_sc_hd__a21bo_1 c421 (.A1(clknet_1_1__leaf_net238),
    .A2(net865),
    .B1_N(net657),
    .X(net332));
 sky130_fd_sc_hd__sdfrtn_1 c422 (.CLK_N(clknet_4_2_0_clk),
    .D(net1079),
    .RESET_B(clknet_1_0__leaf_net331),
    .SCD(net657),
    .SCE(net1083),
    .Q(net333));
 sky130_fd_sc_hd__sdfbbn_2 c423 (.CLK_N(clknet_4_2_0_clk),
    .D(net200),
    .RESET_B(clknet_1_0__leaf_net332),
    .SCD(net999),
    .SCE(net987),
    .SET_B(net1079),
    .Q(net335),
    .Q_N(net334));
 sky130_fd_sc_hd__mux4_1 c424 (.A0(net880),
    .A1(clknet_1_0__leaf_net330),
    .A2(net335),
    .A3(clknet_1_0__leaf_net331),
    .S0(net317),
    .S1(net329),
    .X(net336));
 sky130_fd_sc_hd__a41o_1 c425 (.A1(net220),
    .A2(net880),
    .A3(clknet_1_0__leaf_net331),
    .A4(net882),
    .B1(net804),
    .X(net337));
 sky130_fd_sc_hd__a41o_1 c426 (.A1(clknet_1_0__leaf_net332),
    .A2(net999),
    .A3(net214),
    .A4(net1084),
    .B1(net805),
    .X(net338));
 sky130_fd_sc_hd__sdfbbn_2 c427 (.CLK_N(clknet_4_3_0_clk),
    .D(net329),
    .RESET_B(net990),
    .SCD(clknet_1_0__leaf_net331),
    .SCE(clknet_1_0__leaf_net330),
    .SET_B(net220),
    .Q(net340),
    .Q_N(net339));
 sky130_fd_sc_hd__sdfbbp_1 c428 (.CLK(clknet_4_2_0_clk),
    .D(net333),
    .RESET_B(net980),
    .SCD(net987),
    .SCE(net334),
    .SET_B(net200),
    .Q(net342),
    .Q_N(net341));
 sky130_fd_sc_hd__sdfrtp_2 c429 (.CLK(clknet_4_2_0_clk),
    .D(net340),
    .RESET_B(net324),
    .SCD(net333),
    .SCE(net650),
    .Q(net343));
 sky130_fd_sc_hd__mux4_1 c430 (.A0(net343),
    .A1(net315),
    .A2(net896),
    .A3(net341),
    .S0(net1026),
    .S1(net802),
    .X(net344));
 sky130_fd_sc_hd__mux4_2 c431 (.A0(net999),
    .A1(net232),
    .A2(net343),
    .A3(net333),
    .S0(net985),
    .S1(net804),
    .X(net345));
 sky130_fd_sc_hd__sdfbbn_1 c432 (.CLK_N(clknet_4_3_0_clk),
    .D(net342),
    .RESET_B(clknet_1_0__leaf_net331),
    .SCD(net980),
    .SCE(net343),
    .SET_B(net1084),
    .Q(net347),
    .Q_N(net346));
 sky130_fd_sc_hd__mux4_1 c433 (.A0(net316),
    .A1(net321),
    .A2(net347),
    .A3(net339),
    .S0(net343),
    .S1(net802),
    .X(net348));
 sky130_fd_sc_hd__mux4_1 c434 (.A0(net202),
    .A1(clknet_1_0__leaf_net332),
    .A2(net340),
    .A3(net980),
    .S0(net985),
    .S1(net650),
    .X(net349));
 sky130_fd_sc_hd__mux4_1 c435 (.A0(net324),
    .A1(net232),
    .A2(net229),
    .A3(net342),
    .S0(net321),
    .S1(net806),
    .X(net350));
 sky130_fd_sc_hd__mux4_1 c436 (.A0(net1069),
    .A1(net339),
    .A2(net329),
    .A3(net315),
    .S0(net805),
    .S1(net1023),
    .X(net351));
 sky130_fd_sc_hd__mux4_1 c437 (.A0(net351),
    .A1(net345),
    .A2(net333),
    .A3(net220),
    .S0(net343),
    .S1(net1023),
    .X(net352));
 sky130_fd_sc_hd__mux4_1 c438 (.A0(net222),
    .A1(clknet_1_0__leaf_net332),
    .A2(net990),
    .A3(net650),
    .S0(net800),
    .S1(net804),
    .X(net353));
 sky130_fd_sc_hd__mux4_1 c439 (.A0(net348),
    .A1(net228),
    .A2(net346),
    .A3(net232),
    .S0(net351),
    .S1(net807),
    .X(net354));
 sky130_fd_sc_hd__mux4_1 c440 (.A0(net231),
    .A1(clknet_1_1__leaf_net331),
    .A2(clknet_1_1__leaf_net332),
    .A3(net204),
    .S0(net913),
    .S1(net676),
    .X(net355));
 sky130_fd_sc_hd__a41o_1 c441 (.A1(net342),
    .A2(net1035),
    .A3(net908),
    .A4(net1047),
    .B1(clknet_1_0__leaf_net799),
    .X(net356));
 sky130_fd_sc_hd__sdfbbn_2 c442 (.CLK_N(clknet_4_3_0_clk),
    .D(net356),
    .RESET_B(net237),
    .SCD(clknet_1_0__leaf_net331),
    .SCE(net214),
    .SET_B(net1047),
    .Q(net932),
    .Q_N(net357));
 sky130_fd_sc_hd__a21bo_1 c443 (.A1(net913),
    .A2(net908),
    .B1_N(net249),
    .X(net358));
 sky130_fd_sc_hd__sdfbbp_1 c444 (.CLK(clknet_4_6_0_clk),
    .D(net358),
    .RESET_B(net950),
    .SCD(net124),
    .SCE(clknet_1_0__leaf_net257),
    .SET_B(net1073),
    .Q(net360),
    .Q_N(net359));
 sky130_fd_sc_hd__a31o_1 c445 (.A1(clknet_1_0__leaf_net245),
    .A2(net345),
    .A3(net358),
    .B1(net913),
    .X(net361));
 sky130_fd_sc_hd__a31o_1 c446 (.A1(net345),
    .A2(net734),
    .A3(net1028),
    .B1(net758),
    .X(net362));
 sky130_fd_sc_hd__sdfbbn_1 c447 (.CLK_N(clknet_4_3_0_clk),
    .D(net360),
    .RESET_B(clknet_1_1__leaf_net332),
    .SCD(net882),
    .SCE(net1018),
    .SET_B(net808),
    .Q(net364),
    .Q_N(net363));
 sky130_fd_sc_hd__a21bo_1 c448 (.A1(net360),
    .A2(net341),
    .B1_N(net1023),
    .X(net365));
 sky130_fd_sc_hd__a31o_1 c449 (.A1(net365),
    .A2(net1048),
    .A3(net1029),
    .B1(net783),
    .X(net366));
 sky130_fd_sc_hd__mux4_1 c450 (.A0(clknet_1_0__leaf_net257),
    .A1(net359),
    .A2(net365),
    .A3(net204),
    .S0(net346),
    .S1(net1026),
    .X(net367));
 sky130_fd_sc_hd__mux4_2 c451 (.A0(net124),
    .A1(net364),
    .A2(net991),
    .A3(net1005),
    .S0(net784),
    .S1(net808),
    .X(net368));
 sky130_fd_sc_hd__mux4_1 c452 (.A0(net368),
    .A1(net889),
    .A2(net363),
    .A3(clknet_1_0__leaf_net246),
    .S0(net113),
    .S1(net684),
    .X(net369));
 sky130_fd_sc_hd__mux4_1 c453 (.A0(net365),
    .A1(net359),
    .A2(clknet_1_1__leaf_net369),
    .A3(net341),
    .S0(net212),
    .S1(net676),
    .X(net370));
 sky130_fd_sc_hd__mux4_1 c454 (.A0(net347),
    .A1(net342),
    .A2(net366),
    .A3(net896),
    .S0(net995),
    .S1(net953),
    .X(net371));
 sky130_fd_sc_hd__a31o_1 c455 (.A1(net357),
    .A2(net113),
    .A3(net953),
    .B1(net785),
    .X(net372));
 sky130_fd_sc_hd__mux4_2 c456 (.A0(net1038),
    .A1(net346),
    .A2(net992),
    .A3(net1029),
    .S0(net758),
    .S1(net807),
    .X(net373));
 sky130_fd_sc_hd__a41o_1 c457 (.A1(net366),
    .A2(net371),
    .A3(net992),
    .A4(clknet_1_1__leaf_net332),
    .B1(net713),
    .X(net374));
 sky130_fd_sc_hd__a41o_1 c458 (.A1(net347),
    .A2(net357),
    .A3(net684),
    .A4(net713),
    .B1(net1027),
    .X(net375));
 sky130_fd_sc_hd__a41o_2 c459 (.A1(net371),
    .A2(net373),
    .A3(net672),
    .A4(net1026),
    .B1(net807),
    .X(net376));
 sky130_fd_sc_hd__mux4_2 c460 (.A0(net375),
    .A1(net1046),
    .A2(net363),
    .A3(net993),
    .S0(net376),
    .S1(net672),
    .X(net377));
 sky130_fd_sc_hd__a41o_4 c461 (.A1(net242),
    .A2(net377),
    .A3(net376),
    .A4(net368),
    .B1(net375),
    .X(net378));
 sky130_fd_sc_hd__mux4_1 c462 (.A0(net315),
    .A1(net377),
    .A2(clknet_1_1__leaf_net946),
    .A3(net12),
    .S0(net284),
    .S1(net807),
    .X(net952));
 sky130_fd_sc_hd__mux4_1 c463 (.A0(net12),
    .A1(net932),
    .A2(net209),
    .A3(net378),
    .S0(net792),
    .S1(net800),
    .X(net379));
 sky130_fd_sc_hd__mux4_1 c464 (.A0(clknet_1_0__leaf_net952),
    .A1(net1042),
    .A2(net992),
    .A3(clknet_1_0__leaf_net778),
    .S0(net795),
    .S1(net808),
    .X(net380));
 sky130_fd_sc_hd__mux4_1 c465 (.A0(net377),
    .A1(clknet_1_0__leaf_net330),
    .A2(clknet_1_1__leaf_net331),
    .A3(net992),
    .S0(net738),
    .S1(net787),
    .X(net381));
 sky130_fd_sc_hd__mux4_1 c466 (.A0(net281),
    .A1(net1045),
    .A2(net1005),
    .A3(net378),
    .S0(net808),
    .S1(net810),
    .X(net382));
 sky130_fd_sc_hd__mux4_1 c467 (.A0(clknet_1_0__leaf_net369),
    .A1(net377),
    .A2(net793),
    .A3(net795),
    .S0(clknet_1_1__leaf_net799),
    .S1(net1023),
    .X(net383));
 sky130_fd_sc_hd__mux4_1 c468 (.A0(clknet_1_0__leaf_net369),
    .A1(clknet_1_1__leaf_net952),
    .A2(net738),
    .A3(net793),
    .S0(net807),
    .S1(net810),
    .X(net384));
 sky130_fd_sc_hd__mux4_1 c469 (.A0(clknet_1_1__leaf_net330),
    .A1(net329),
    .A2(net962),
    .A3(net793),
    .S0(net1022),
    .S1(net809),
    .X(net385));
 sky130_fd_sc_hd__mux4_1 c470 (.A0(clknet_1_1__leaf_net946),
    .A1(net1052),
    .A2(net955),
    .A3(net1023),
    .S0(net1022),
    .S1(net810),
    .X(net386));
 sky130_fd_sc_hd__mux4_1 c471 (.A0(net378),
    .A1(net955),
    .A2(net801),
    .A3(net807),
    .S0(net1022),
    .S1(net809),
    .X(net387));
 sky130_fd_sc_hd__mux4_1 c472 (.A0(clknet_1_1__leaf_net330),
    .A1(clknet_1_1__leaf_net952),
    .A2(net738),
    .A3(net1025),
    .S0(net808),
    .S1(net1022),
    .X(net388));
 sky130_fd_sc_hd__mux4_1 c473 (.A0(clknet_1_1__leaf_net331),
    .A1(clknet_1_1__leaf_net369),
    .A2(net997),
    .A3(net738),
    .S0(net792),
    .S1(clknet_1_1__leaf_net799),
    .X(net389));
 sky130_fd_sc_hd__mux4_1 c474 (.A0(net950),
    .A1(net19),
    .A2(net738),
    .A3(net976),
    .S0(net1022),
    .S1(net812),
    .X(net390));
 sky130_fd_sc_hd__mux4_2 c475 (.A0(net950),
    .A1(net962),
    .A2(net1026),
    .A3(net785),
    .S0(net1022),
    .S1(net809),
    .X(net391));
 sky130_fd_sc_hd__mux4_1 c476 (.A0(net329),
    .A1(net391),
    .A2(net281),
    .A3(clknet_1_1__leaf_net386),
    .S0(net787),
    .S1(net810),
    .X(net392));
 sky130_fd_sc_hd__mux4_1 c477 (.A0(net7),
    .A1(net391),
    .A2(net12),
    .A3(net955),
    .S0(net812),
    .S1(net978),
    .X(net393));
 sky130_fd_sc_hd__mux4_2 c478 (.A0(net391),
    .A1(net393),
    .A2(net1038),
    .A3(net801),
    .S0(net811),
    .S1(net978),
    .X(net394));
 sky130_fd_sc_hd__mux4_1 c479 (.A0(net393),
    .A1(clknet_1_1__leaf_net952),
    .A2(clknet_1_1__leaf_net330),
    .A3(clknet_1_1__leaf_net799),
    .S0(net807),
    .S1(net812),
    .X(net395));
 sky130_fd_sc_hd__mux4_1 c480 (.A0(net390),
    .A1(net391),
    .A2(clknet_1_1__leaf_net245),
    .A3(net281),
    .S0(net1022),
    .S1(net811),
    .X(net396));
 sky130_fd_sc_hd__mux4_1 c481 (.A0(clknet_1_1__leaf_net396),
    .A1(net1040),
    .A2(net391),
    .A3(clknet_1_1__leaf_net946),
    .S0(net784),
    .S1(net795),
    .X(net397));
 sky130_fd_sc_hd__mux4_1 c482 (.A0(clknet_1_0__leaf_net397),
    .A1(net1040),
    .A2(clknet_1_1__leaf_net946),
    .A3(net738),
    .S0(net978),
    .S1(net813),
    .X(net398));
 sky130_fd_sc_hd__mux4_1 c483 (.A0(net391),
    .A1(clknet_1_0__leaf_net396),
    .A2(clknet_1_1__leaf_net397),
    .A3(net962),
    .S0(net978),
    .S1(net813),
    .X(net399));
 sky130_fd_sc_hd__mux4_1 c484 (.A0(net932),
    .A1(clknet_1_0__leaf_net300),
    .A2(net771),
    .A3(net796),
    .S0(clknet_1_1__leaf_net798),
    .S1(net939),
    .X(net400));
 sky130_fd_sc_hd__mux4_2 c485 (.A0(net1038),
    .A1(clknet_1_1__leaf_net300),
    .A2(clknet_1_0__leaf_net947),
    .A3(net940),
    .S0(net1008),
    .S1(net1022),
    .X(net401));
 sky130_fd_sc_hd__mux4_1 c486 (.A0(net377),
    .A1(net329),
    .A2(net295),
    .A3(net926),
    .S0(net768),
    .S1(net951),
    .X(net402));
 sky130_fd_sc_hd__mux4_2 c487 (.A0(clknet_1_0__leaf_net401),
    .A1(net339),
    .A2(net764),
    .A3(net768),
    .S0(net769),
    .S1(net770),
    .X(net403));
 sky130_fd_sc_hd__mux4_1 c488 (.A0(net119),
    .A1(net340),
    .A2(net1036),
    .A3(clknet_1_0__leaf_net403),
    .S0(net1010),
    .S1(net787),
    .X(net404));
 sky130_fd_sc_hd__mux4_1 c489 (.A0(clknet_1_0__leaf_net403),
    .A1(net997),
    .A2(net113),
    .A3(clknet_1_1__leaf_net946),
    .S0(clknet_1_0__leaf_net401),
    .S1(clknet_1_0__leaf_net300),
    .X(net405));
 sky130_fd_sc_hd__mux4_1 c490 (.A0(clknet_1_1__leaf_net401),
    .A1(net296),
    .A2(clknet_1_1__leaf_net300),
    .A3(clknet_1_1__leaf_net403),
    .S0(net1030),
    .S1(net735),
    .X(net406));
 sky130_fd_sc_hd__mux4_2 c491 (.A0(net908),
    .A1(clknet_1_1__leaf_net946),
    .A2(clknet_1_1__leaf_net401),
    .A3(clknet_1_1__leaf_net945),
    .S0(clknet_1_0__leaf_net762),
    .S1(clknet_1_1__leaf_net927),
    .X(net977));
 sky130_fd_sc_hd__mux4_1 c492 (.A0(net400),
    .A1(clknet_1_1__leaf_net403),
    .A2(net930),
    .A3(net988),
    .S0(clknet_1_0__leaf_net945),
    .S1(net951),
    .X(net407));
 sky130_fd_sc_hd__mux4_1 c493 (.A0(clknet_1_1__leaf_net403),
    .A1(net943),
    .A2(net735),
    .A3(net929),
    .S0(net768),
    .S1(clknet_1_1__leaf_net815),
    .X(net408));
 sky130_fd_sc_hd__mux4_1 c494 (.A0(clknet_1_0__leaf_net302),
    .A1(clknet_1_0__leaf_net403),
    .A2(clknet_1_0__leaf_net401),
    .A3(net814),
    .S0(clknet_1_0__leaf_net815),
    .S1(clknet_1_0__leaf_net924),
    .X(net409));
 sky130_fd_sc_hd__mux4_1 c495 (.A0(net940),
    .A1(clknet_1_0__leaf_net977),
    .A2(net950),
    .A3(net735),
    .S0(clknet_1_1__leaf_net798),
    .S1(net816),
    .X(net410));
 sky130_fd_sc_hd__mux4_1 c496 (.A0(clknet_1_0__leaf_net303),
    .A1(net209),
    .A2(net943),
    .A3(clknet_1_0__leaf_net403),
    .S0(clknet_1_0__leaf_net945),
    .S1(net763),
    .X(net411));
 sky130_fd_sc_hd__mux4_1 c497 (.A0(net329),
    .A1(clknet_1_1__leaf_net977),
    .A2(clknet_1_1__leaf_net403),
    .A3(net929),
    .S0(net796),
    .S1(clknet_1_1__leaf_net815),
    .X(net412));
 sky130_fd_sc_hd__mux4_2 c498 (.A0(net340),
    .A1(clknet_1_0__leaf_net977),
    .A2(net962),
    .A3(net770),
    .S0(clknet_1_1__leaf_net798),
    .S1(net818),
    .X(net413));
 sky130_fd_sc_hd__mux4_1 c499 (.A0(clknet_1_0__leaf_net947),
    .A1(clknet_1_1__leaf_net403),
    .A2(net768),
    .A3(net771),
    .S0(net787),
    .S1(net819),
    .X(net414));
 sky130_fd_sc_hd__mux4_1 c500 (.A0(net115),
    .A1(net213),
    .A2(net940),
    .A3(net926),
    .S0(net735),
    .S1(clknet_1_1__leaf_net815),
    .X(net415));
 sky130_fd_sc_hd__mux4_2 c501 (.A0(clknet_1_0__leaf_net947),
    .A1(net735),
    .A2(net787),
    .A3(clknet_1_1__leaf_net927),
    .S0(net819),
    .S1(net821),
    .X(net954));
 sky130_fd_sc_hd__mux4_2 c502 (.A0(net1008),
    .A1(net1003),
    .A2(net735),
    .A3(net770),
    .S0(net814),
    .S1(net820),
    .X(net948));
 sky130_fd_sc_hd__mux4_2 c503 (.A0(net993),
    .A1(net948),
    .A2(clknet_1_1__leaf_net401),
    .A3(clknet_1_0__leaf_net954),
    .S0(net953),
    .S1(net820),
    .X(net938));
 sky130_fd_sc_hd__mux4_1 c504 (.A0(net948),
    .A1(clknet_1_0__leaf_net938),
    .A2(clknet_1_0__leaf_net954),
    .A3(clknet_1_1__leaf_net977),
    .S0(net962),
    .S1(net818),
    .X(net416));
 sky130_fd_sc_hd__mux4_2 c505 (.A0(net104),
    .A1(net948),
    .A2(clknet_1_0__leaf_net938),
    .A3(net943),
    .S0(clknet_1_1__leaf_net403),
    .S1(net725),
    .X(net417));
 sky130_fd_sc_hd__a21bo_2 c528 (.A1(net207),
    .A2(net994),
    .B1_N(net982),
    .X(net418));
 sky130_fd_sc_hd__a21bo_2 c529 (.A1(net1065),
    .A2(net320),
    .B1_N(net1048),
    .X(net419));
 sky130_fd_sc_hd__a21bo_1 c530 (.A1(net981),
    .A2(net201),
    .B1_N(net1048),
    .X(net420));
 sky130_fd_sc_hd__clkbuf_4 c531 (.A(net737),
    .X(net928));
 sky130_fd_sc_hd__a41o_1 c532 (.A1(net201),
    .A2(net981),
    .A3(net990),
    .A4(net321),
    .B1(net803),
    .X(net421));
 sky130_fd_sc_hd__buf_1 c533 (.A(net737),
    .X(net422));
 sky130_fd_sc_hd__buf_1 c534 (.A(clknet_1_0__leaf_net706),
    .X(net423));
 sky130_fd_sc_hd__buf_2 c535 (.A(net737),
    .X(net424));
 sky130_fd_sc_hd__a21bo_1 c536 (.A1(net424),
    .A2(net1017),
    .B1_N(clknet_1_0__leaf_net423),
    .X(net934));
 sky130_fd_sc_hd__buf_1 c537 (.A(clknet_1_0__leaf_net706),
    .X(net425));
 sky130_fd_sc_hd__sdfrtp_1 c538 (.CLK(clknet_4_0_0_clk),
    .D(clknet_1_0__leaf_net423),
    .RESET_B(net994),
    .SCD(net981),
    .SCE(net419),
    .Q(net426));
 sky130_fd_sc_hd__a41o_1 c539 (.A1(net208),
    .A2(clknet_1_1__leaf_net425),
    .A3(net420),
    .A4(net1017),
    .B1(net1048),
    .X(net427));
 sky130_fd_sc_hd__sdfbbn_1 c540 (.CLK_N(clknet_4_0_0_clk),
    .D(net419),
    .RESET_B(clknet_1_1__leaf_net425),
    .SCD(net995),
    .SCE(net217),
    .SET_B(net426),
    .Q(net429),
    .Q_N(net428));
 sky130_fd_sc_hd__clkbuf_1 c541 (.A(net737),
    .X(net430));
 sky130_fd_sc_hd__a21bo_1 c542 (.A1(net429),
    .A2(net430),
    .B1_N(net426),
    .X(net431));
 sky130_fd_sc_hd__mux4_1 c543 (.A0(net426),
    .A1(net428),
    .A2(clknet_1_1__leaf_net425),
    .A3(net928),
    .S0(net207),
    .S1(net418),
    .X(net432));
 sky130_fd_sc_hd__mux4_1 c544 (.A0(net1017),
    .A1(clknet_1_0__leaf_net934),
    .A2(clknet_1_1__leaf_net425),
    .A3(net321),
    .S0(net986),
    .S1(net803),
    .X(net433));
 sky130_fd_sc_hd__mux4_1 c545 (.A0(clknet_1_1__leaf_net423),
    .A1(net426),
    .A2(net321),
    .A3(net419),
    .S0(net1042),
    .S1(net424),
    .X(net434));
 sky130_fd_sc_hd__mux4_1 c546 (.A0(net217),
    .A1(net424),
    .A2(clknet_1_0__leaf_net433),
    .A3(net723),
    .S0(net726),
    .S1(net822),
    .X(net435));
 sky130_fd_sc_hd__mux4_1 c547 (.A0(clknet_1_0__leaf_net433),
    .A1(net431),
    .A2(net424),
    .A3(clknet_1_0__leaf_net425),
    .S0(net321),
    .S1(net822),
    .X(net436));
 sky130_fd_sc_hd__mux4_1 c548 (.A0(clknet_1_1__leaf_net433),
    .A1(net428),
    .A2(net419),
    .A3(net723),
    .S0(net730),
    .S1(net823),
    .X(net437));
 sky130_fd_sc_hd__mux4_1 c549 (.A0(net1046),
    .A1(net986),
    .A2(net1017),
    .A3(net420),
    .S0(net730),
    .S1(net737),
    .X(net438));
 sky130_fd_sc_hd__a41o_1 c550 (.A1(net986),
    .A2(net335),
    .A3(net985),
    .A4(net1023),
    .B1(net823),
    .X(net439));
 sky130_fd_sc_hd__a31o_1 c551 (.A1(net882),
    .A2(net986),
    .A3(net1043),
    .B1(net1092),
    .X(net440));
 sky130_fd_sc_hd__a41o_2 c552 (.A1(net439),
    .A2(net986),
    .A3(net228),
    .A4(net440),
    .B1(net1075),
    .X(net441));
 sky130_fd_sc_hd__a21bo_1 c553 (.A1(net335),
    .A2(net1043),
    .B1_N(net823),
    .X(net442));
 sky130_fd_sc_hd__a41o_2 c554 (.A1(net442),
    .A2(net335),
    .A3(net1046),
    .A4(net726),
    .B1(net1023),
    .X(net443));
 sky130_fd_sc_hd__a41o_1 c555 (.A1(net237),
    .A2(net441),
    .A3(net334),
    .A4(net726),
    .B1(net804),
    .X(net444));
 sky130_fd_sc_hd__a31o_1 c556 (.A1(net443),
    .A2(net1047),
    .A3(net685),
    .B1(net757),
    .X(net445));
 sky130_fd_sc_hd__a21bo_1 c557 (.A1(net981),
    .A2(net442),
    .B1_N(net806),
    .X(net446));
 sky130_fd_sc_hd__a31o_1 c558 (.A1(net321),
    .A2(net335),
    .A3(net222),
    .B1(net822),
    .X(net447));
 sky130_fd_sc_hd__sdfrtp_4 c559 (.CLK(clknet_4_0_0_clk),
    .D(net439),
    .RESET_B(net441),
    .SCD(net237),
    .SCE(net442),
    .Q(net925));
 sky130_fd_sc_hd__mux4_2 c560 (.A0(net429),
    .A1(net228),
    .A2(net889),
    .A3(net650),
    .S0(net805),
    .S1(net806),
    .X(net448));
 sky130_fd_sc_hd__a41o_1 c561 (.A1(net446),
    .A2(net228),
    .A3(net1047),
    .A4(net979),
    .B1(net1081),
    .X(net449));
 sky130_fd_sc_hd__a41o_1 c562 (.A1(net445),
    .A2(net428),
    .A3(net439),
    .A4(net1094),
    .B1(net804),
    .X(net450));
 sky130_fd_sc_hd__sdfbbp_1 c563 (.CLK(clknet_4_1_0_clk),
    .D(net925),
    .RESET_B(net979),
    .SCD(net445),
    .SCE(net986),
    .SET_B(net685),
    .Q(net452),
    .Q_N(net451));
 sky130_fd_sc_hd__a41o_1 c564 (.A1(net429),
    .A2(net443),
    .A3(net452),
    .A4(net986),
    .B1(net448),
    .X(net453));
 sky130_fd_sc_hd__sdfbbn_2 c565 (.CLK_N(clknet_4_1_0_clk),
    .D(net453),
    .RESET_B(net421),
    .SCD(net439),
    .SCE(net979),
    .SET_B(net228),
    .Q(net455),
    .Q_N(net454));
 sky130_fd_sc_hd__a41o_2 c566 (.A1(net222),
    .A2(net454),
    .A3(net757),
    .A4(net802),
    .B1(net805),
    .X(net931));
 sky130_fd_sc_hd__mux4_1 c567 (.A0(net441),
    .A1(net452),
    .A2(net454),
    .A3(net439),
    .S0(net925),
    .S1(net979),
    .X(net456));
 sky130_fd_sc_hd__a31o_1 c568 (.A1(net447),
    .A2(net455),
    .A3(net931),
    .B1(net1080),
    .X(net457));
 sky130_fd_sc_hd__mux4_1 c569 (.A0(net450),
    .A1(net979),
    .A2(net995),
    .A3(net685),
    .S0(net726),
    .S1(net1082),
    .X(net458));
 sky130_fd_sc_hd__mux4_1 c570 (.A0(net447),
    .A1(net454),
    .A2(net451),
    .A3(net453),
    .S0(net685),
    .S1(net825),
    .X(net459));
 sky130_fd_sc_hd__mux4_1 c571 (.A0(net440),
    .A1(net231),
    .A2(net446),
    .A3(net726),
    .S0(net805),
    .S1(net936),
    .X(net460));
 sky130_fd_sc_hd__mux4_2 c572 (.A0(net376),
    .A1(clknet_1_0__leaf_net934),
    .A2(net882),
    .A3(net1018),
    .S0(net995),
    .S1(net822),
    .X(net461));
 sky130_fd_sc_hd__mux4_1 c573 (.A0(clknet_1_0__leaf_net246),
    .A1(net440),
    .A2(net1017),
    .A3(net1036),
    .S0(net448),
    .S1(net368),
    .X(net462));
 sky130_fd_sc_hd__mux4_1 c574 (.A0(net1093),
    .A1(net1090),
    .A2(clknet_1_1__leaf_net462),
    .A3(clknet_1_0__leaf_net369),
    .S0(net378),
    .S1(net992),
    .X(net463));
 sky130_fd_sc_hd__mux4_1 c575 (.A0(net368),
    .A1(net990),
    .A2(net1027),
    .A3(clknet_1_1__leaf_net778),
    .S0(net806),
    .S1(net826),
    .X(net464));
 sky130_fd_sc_hd__mux4_1 c576 (.A0(net364),
    .A1(net988),
    .A2(net995),
    .A3(clknet_1_0__leaf_net934),
    .S0(net1018),
    .S1(net783),
    .X(net465));
 sky130_fd_sc_hd__mux4_1 c577 (.A0(net440),
    .A1(clknet_1_0__leaf_net462),
    .A2(net376),
    .A3(net1046),
    .S0(clknet_1_0__leaf_net465),
    .S1(net1000),
    .X(net466));
 sky130_fd_sc_hd__mux4_1 c578 (.A0(net1089),
    .A1(net988),
    .A2(net726),
    .A3(net806),
    .S0(net936),
    .S1(net828),
    .X(net467));
 sky130_fd_sc_hd__mux4_1 c579 (.A0(net995),
    .A1(net1090),
    .A2(clknet_1_1__leaf_net465),
    .A3(net1005),
    .S0(clknet_1_0__leaf_net462),
    .S1(net376),
    .X(net468));
 sky130_fd_sc_hd__mux4_1 c580 (.A0(net452),
    .A1(net992),
    .A2(net988),
    .A3(clknet_1_0__leaf_net461),
    .S0(net806),
    .S1(net828),
    .X(net469));
 sky130_fd_sc_hd__mux4_1 c581 (.A0(net995),
    .A1(net992),
    .A2(clknet_1_0__leaf_net462),
    .A3(clknet_1_0__leaf_net465),
    .S0(net824),
    .S1(net829),
    .X(net470));
 sky130_fd_sc_hd__mux4_1 c582 (.A0(net1089),
    .A1(clknet_1_0__leaf_net465),
    .A2(net889),
    .A3(net822),
    .S0(net826),
    .S1(net830),
    .X(net471));
 sky130_fd_sc_hd__mux4_1 c583 (.A0(net464),
    .A1(net1089),
    .A2(clknet_1_0__leaf_net471),
    .A3(net1030),
    .S0(net713),
    .S1(net822),
    .X(net472));
 sky130_fd_sc_hd__mux4_1 c584 (.A0(clknet_1_1__leaf_net471),
    .A1(net213),
    .A2(net364),
    .A3(net1062),
    .S0(net1090),
    .S1(net830),
    .X(net473));
 sky130_fd_sc_hd__mux4_1 c585 (.A0(net1090),
    .A1(clknet_1_0__leaf_net461),
    .A2(net896),
    .A3(net715),
    .S0(net758),
    .S1(net830),
    .X(net474));
 sky130_fd_sc_hd__mux4_1 c586 (.A0(net928),
    .A1(clknet_1_0__leaf_net246),
    .A2(net825),
    .A3(net936),
    .S0(net830),
    .S1(net831),
    .X(net475));
 sky130_fd_sc_hd__mux4_1 c587 (.A0(clknet_1_1__leaf_net465),
    .A1(clknet_1_1__leaf_net461),
    .A2(net991),
    .A3(clknet_1_1__leaf_net475),
    .S0(clknet_1_0__leaf_net469),
    .S1(clknet_1_0__leaf_net462),
    .X(net476));
 sky130_fd_sc_hd__mux4_1 c588 (.A0(net1018),
    .A1(clknet_1_1__leaf_net474),
    .A2(clknet_1_1__leaf_net475),
    .A3(net825),
    .S0(net829),
    .S1(net831),
    .X(net477));
 sky130_fd_sc_hd__mux4_1 c589 (.A0(net932),
    .A1(net1093),
    .A2(net310),
    .A3(clknet_1_1__leaf_net465),
    .S0(clknet_1_0__leaf_net475),
    .S1(net737),
    .X(net478));
 sky130_fd_sc_hd__mux4_1 c590 (.A0(clknet_1_0__leaf_net475),
    .A1(net378),
    .A2(net1026),
    .A3(net1023),
    .S0(net829),
    .S1(net830),
    .X(net479));
 sky130_fd_sc_hd__mux4_1 c591 (.A0(clknet_1_1__leaf_net475),
    .A1(clknet_1_1__leaf_net469),
    .A2(net715),
    .A3(net724),
    .S0(net758),
    .S1(net1023),
    .X(net480));
 sky130_fd_sc_hd__mux4_2 c592 (.A0(net1003),
    .A1(net684),
    .A2(net717),
    .A3(net724),
    .S0(net737),
    .S1(net936),
    .X(net481));
 sky130_fd_sc_hd__mux4_1 c593 (.A0(clknet_1_0__leaf_net469),
    .A1(clknet_1_0__leaf_net475),
    .A2(net481),
    .A3(clknet_1_1__leaf_net465),
    .S0(net717),
    .S1(net724),
    .X(net482));
 sky130_fd_sc_hd__mux4_1 c594 (.A0(net19),
    .A1(net448),
    .A2(net928),
    .A3(clknet_1_1__leaf_net934),
    .S0(net1042),
    .S1(net1002),
    .X(net483));
 sky130_fd_sc_hd__mux4_1 c595 (.A0(net467),
    .A1(net992),
    .A2(net1018),
    .A3(net976),
    .S0(net789),
    .S1(net978),
    .X(net484));
 sky130_fd_sc_hd__mux4_1 c596 (.A0(net448),
    .A1(clknet_1_1__leaf_net934),
    .A2(net789),
    .A3(net939),
    .S0(net936),
    .S1(net827),
    .X(net485));
 sky130_fd_sc_hd__mux4_1 c597 (.A0(net19),
    .A1(net928),
    .A2(clknet_1_1__leaf_net483),
    .A3(net717),
    .S0(net1024),
    .S1(net814),
    .X(net486));
 sky130_fd_sc_hd__mux4_2 c598 (.A0(net991),
    .A1(net19),
    .A2(net684),
    .A3(net962),
    .S0(net783),
    .S1(net831),
    .X(net487));
 sky130_fd_sc_hd__mux4_1 c599 (.A0(clknet_1_1__leaf_net461),
    .A1(net394),
    .A2(net19),
    .A3(clknet_1_0__leaf_net952),
    .S0(net1002),
    .S1(net814),
    .X(net488));
 sky130_fd_sc_hd__mux4_1 c600 (.A0(net486),
    .A1(net1041),
    .A2(net992),
    .A3(net454),
    .S0(net721),
    .S1(net831),
    .X(net489));
 sky130_fd_sc_hd__mux4_2 c601 (.A0(net448),
    .A1(net985),
    .A2(clknet_1_1__leaf_net934),
    .A3(net928),
    .S0(net212),
    .S1(net831),
    .X(net490));
 sky130_fd_sc_hd__mux4_1 c602 (.A0(net484),
    .A1(net19),
    .A2(net1018),
    .A3(net481),
    .S0(net212),
    .S1(net826),
    .X(net491));
 sky130_fd_sc_hd__mux4_2 c603 (.A0(net487),
    .A1(net481),
    .A2(net1042),
    .A3(net721),
    .S0(net731),
    .S1(net978),
    .X(net492));
 sky130_fd_sc_hd__mux4_2 c604 (.A0(clknet_1_0__leaf_net490),
    .A1(net1002),
    .A2(net467),
    .A3(clknet_1_1__leaf_net483),
    .S0(net731),
    .S1(net789),
    .X(net493));
 sky130_fd_sc_hd__mux4_1 c605 (.A0(clknet_1_0__leaf_net493),
    .A1(net394),
    .A2(net284),
    .A3(net487),
    .S0(net1002),
    .S1(net721),
    .X(net494));
 sky130_fd_sc_hd__mux4_1 c606 (.A0(clknet_1_1__leaf_net493),
    .A1(net988),
    .A2(net492),
    .A3(net487),
    .S0(net993),
    .S1(net939),
    .X(net495));
 sky130_fd_sc_hd__mux4_1 c607 (.A0(net485),
    .A1(net492),
    .A2(net237),
    .A3(net378),
    .S0(net789),
    .S1(clknet_1_0__leaf_net833),
    .X(net496));
 sky130_fd_sc_hd__mux4_1 c608 (.A0(net394),
    .A1(clknet_1_0__leaf_net493),
    .A2(net683),
    .A3(net783),
    .S0(net831),
    .S1(clknet_1_0__leaf_net833),
    .X(net497));
 sky130_fd_sc_hd__mux4_1 c609 (.A0(net882),
    .A1(net487),
    .A2(net1024),
    .A3(net1022),
    .S0(clknet_1_0__leaf_net833),
    .S1(clknet_1_1__leaf_net835),
    .X(net498));
 sky130_fd_sc_hd__mux4_1 c610 (.A0(clknet_1_0__leaf_net498),
    .A1(clknet_1_1__leaf_net483),
    .A2(net19),
    .A3(net683),
    .S0(clknet_1_0__leaf_net833),
    .S1(clknet_1_1__leaf_net835),
    .X(net499));
 sky130_fd_sc_hd__mux4_1 c611 (.A0(net113),
    .A1(net1005),
    .A2(clknet_1_1__leaf_net498),
    .A3(net481),
    .S0(net731),
    .S1(net1026),
    .X(net500));
 sky130_fd_sc_hd__mux4_1 c612 (.A0(clknet_1_0__leaf_net499),
    .A1(net1018),
    .A2(clknet_1_0__leaf_net498),
    .A3(clknet_1_0__leaf_net490),
    .S0(net378),
    .S1(clknet_1_0__leaf_net835),
    .X(net501));
 sky130_fd_sc_hd__mux4_1 c613 (.A0(net378),
    .A1(net487),
    .A2(net394),
    .A3(clknet_1_1__leaf_net483),
    .S0(clknet_1_0__leaf_net834),
    .S1(net836),
    .X(net502));
 sky130_fd_sc_hd__mux4_1 c614 (.A0(net492),
    .A1(clknet_1_1__leaf_net499),
    .A2(clknet_1_1__leaf_net490),
    .A3(net682),
    .S0(net831),
    .S1(clknet_1_0__leaf_net835),
    .X(net503));
 sky130_fd_sc_hd__mux4_1 c615 (.A0(clknet_1_1__leaf_net498),
    .A1(net500),
    .A2(net487),
    .A3(clknet_1_1__leaf_net490),
    .S0(net682),
    .S1(net837),
    .X(net504));
 sky130_fd_sc_hd__mux4_1 c616 (.A0(net997),
    .A1(net1018),
    .A2(net821),
    .A3(net827),
    .S0(net933),
    .S1(net838),
    .X(net505));
 sky130_fd_sc_hd__mux4_2 c617 (.A0(net481),
    .A1(net505),
    .A2(net771),
    .A3(net1024),
    .S0(clknet_1_0__leaf_net927),
    .S1(net839),
    .X(net506));
 sky130_fd_sc_hd__mux4_1 c618 (.A0(net1008),
    .A1(clknet_1_1__leaf_net934),
    .A2(net939),
    .A3(net1022),
    .S0(net827),
    .S1(clknet_1_1__leaf_net833),
    .X(net507));
 sky130_fd_sc_hd__mux4_2 c619 (.A0(clknet_1_0__leaf_net506),
    .A1(net997),
    .A2(net357),
    .A3(net930),
    .S0(clknet_1_0__leaf_net927),
    .S1(clknet_1_1__leaf_net834),
    .X(net508));
 sky130_fd_sc_hd__mux4_2 c62 (.A0(net906),
    .A1(net913),
    .A2(net1037),
    .A3(net915),
    .S0(net914),
    .S1(net878),
    .X(net0));
 sky130_fd_sc_hd__mux4_1 c620 (.A0(net1008),
    .A1(clknet_1_0__leaf_net977),
    .A2(net769),
    .A3(clknet_1_0__leaf_net815),
    .S0(net826),
    .S1(net831),
    .X(net509));
 sky130_fd_sc_hd__mux4_2 c621 (.A0(clknet_1_0__leaf_net508),
    .A1(net993),
    .A2(net928),
    .A3(net929),
    .S0(net1024),
    .S1(net839),
    .X(net510));
 sky130_fd_sc_hd__mux4_1 c622 (.A0(clknet_1_0__leaf_net300),
    .A1(clknet_1_0__leaf_net506),
    .A2(net929),
    .A3(net978),
    .S0(net816),
    .S1(clknet_1_1__leaf_net833),
    .X(net511));
 sky130_fd_sc_hd__mux4_1 c623 (.A0(clknet_1_1__leaf_net506),
    .A1(clknet_1_1__leaf_net508),
    .A2(clknet_1_1__leaf_net934),
    .A3(net769),
    .S0(net976),
    .S1(clknet_1_0__leaf_net924),
    .X(net512));
 sky130_fd_sc_hd__mux4_1 c624 (.A0(net511),
    .A1(net481),
    .A2(net1036),
    .A3(clknet_1_0__leaf_net924),
    .S0(net827),
    .S1(net838),
    .X(net513));
 sky130_fd_sc_hd__mux4_1 c625 (.A0(net512),
    .A1(net1008),
    .A2(net213),
    .A3(net925),
    .S0(net820),
    .S1(net944),
    .X(net514));
 sky130_fd_sc_hd__mux4_1 c626 (.A0(net988),
    .A1(net1000),
    .A2(clknet_1_1__leaf_net483),
    .A3(net1008),
    .S0(clknet_1_1__leaf_net510),
    .S1(net827),
    .X(net515));
 sky130_fd_sc_hd__mux4_1 c627 (.A0(net481),
    .A1(net113),
    .A2(net928),
    .A3(net1030),
    .S0(net716),
    .S1(clknet_1_0__leaf_net924),
    .X(net516));
 sky130_fd_sc_hd__mux4_1 c628 (.A0(clknet_1_1__leaf_net508),
    .A1(net930),
    .A2(net1036),
    .A3(clknet_1_0__leaf_net762),
    .S0(net771),
    .S1(net1024),
    .X(net935));
 sky130_fd_sc_hd__mux4_1 c629 (.A0(net455),
    .A1(net507),
    .A2(clknet_1_1__leaf_net483),
    .A3(net928),
    .S0(clknet_1_0__leaf_net927),
    .S1(net836),
    .X(net517));
 sky130_fd_sc_hd__mux4_2 c63 (.A0(net0),
    .A1(net904),
    .A2(net900),
    .A3(net899),
    .S0(net912),
    .S1(net906),
    .X(net1));
 sky130_fd_sc_hd__mux4_1 c630 (.A0(net516),
    .A1(clknet_1_1__leaf_net515),
    .A2(clknet_1_1__leaf_net517),
    .A3(net212),
    .S0(clknet_1_0__leaf_net762),
    .S1(clknet_1_1__leaf_net834),
    .X(net518));
 sky130_fd_sc_hd__mux4_1 c631 (.A0(net455),
    .A1(net1035),
    .A2(net1030),
    .A3(net923),
    .S0(clknet_1_1__leaf_net833),
    .S1(clknet_1_0__leaf_net834),
    .X(net973));
 sky130_fd_sc_hd__mux4_2 c632 (.A0(net896),
    .A1(clknet_1_1__leaf_net973),
    .A2(clknet_1_0__leaf_net510),
    .A3(net814),
    .S0(net817),
    .S1(net933),
    .X(net922));
 sky130_fd_sc_hd__mux4_1 c633 (.A0(net513),
    .A1(clknet_1_1__leaf_net517),
    .A2(clknet_1_0__leaf_net922),
    .A3(clknet_1_0__leaf_net300),
    .S0(clknet_1_0__leaf_net508),
    .S1(net722),
    .X(net519));
 sky130_fd_sc_hd__mux4_1 c634 (.A0(clknet_1_0__leaf_net517),
    .A1(clknet_1_1__leaf_net922),
    .A2(clknet_1_1__leaf_net510),
    .A3(net716),
    .S0(net722),
    .S1(clknet_1_1__leaf_net834),
    .X(net520));
 sky130_fd_sc_hd__mux4_1 c635 (.A0(net213),
    .A1(net1036),
    .A2(net717),
    .A3(net929),
    .S0(clknet_1_0__leaf_net798),
    .S1(clknet_1_0__leaf_net834),
    .X(net521));
 sky130_fd_sc_hd__mux4_2 c636 (.A0(net521),
    .A1(net931),
    .A2(clknet_1_0__leaf_net922),
    .A3(clknet_1_0__leaf_net762),
    .S0(net814),
    .S1(net836),
    .X(net522));
 sky130_fd_sc_hd__mux4_1 c637 (.A0(net514),
    .A1(net284),
    .A2(clknet_1_0__leaf_net515),
    .A3(clknet_1_1__leaf_net510),
    .S0(clknet_1_0__leaf_net517),
    .S1(net722),
    .X(net523));
 sky130_fd_sc_hd__mux4_1 c64 (.A0(net3),
    .A1(net910),
    .A2(net909),
    .A3(net906),
    .S0(net902),
    .S1(net900),
    .X(net2));
 sky130_fd_sc_hd__mux4_2 c65 (.A0(net865),
    .A1(net882),
    .A2(net878),
    .A3(net879),
    .S0(net889),
    .S1(net1044),
    .X(net3));
 sky130_fd_sc_hd__a21bo_2 c66 (.A1(net899),
    .A2(net915),
    .B1_N(net1051),
    .X(net4));
 sky130_fd_sc_hd__buf_1 c660 (.A(net696),
    .X(net524));
 sky130_fd_sc_hd__clkbuf_1 c661 (.A(net696),
    .X(net525));
 sky130_fd_sc_hd__a21bo_1 c662 (.A1(net431),
    .A2(net1014),
    .B1_N(net982),
    .X(net526));
 sky130_fd_sc_hd__mux4_1 c663 (.A0(net1068),
    .A1(net1016),
    .A2(net1002),
    .A3(net981),
    .S0(net1014),
    .S1(net418),
    .X(net527));
 sky130_fd_sc_hd__clkbuf_1 c664 (.A(net719),
    .X(net528));
 sky130_fd_sc_hd__a21bo_1 c665 (.A1(net994),
    .A2(net424),
    .B1_N(net1011),
    .X(net529));
 sky130_fd_sc_hd__a21bo_1 c666 (.A1(net1011),
    .A2(net1014),
    .B1_N(net529),
    .X(net530));
 sky130_fd_sc_hd__a21bo_1 c667 (.A1(net982),
    .A2(net994),
    .B1_N(net823),
    .X(net531));
 sky130_fd_sc_hd__mux4_2 c668 (.A0(net529),
    .A1(net214),
    .A2(net1014),
    .A3(net982),
    .S0(net1011),
    .S1(net723),
    .X(net532));
 sky130_fd_sc_hd__clkbuf_2 c669 (.A(net719),
    .X(net533));
 sky130_fd_sc_hd__a31o_1 c67 (.A1(net902),
    .A2(net907),
    .A3(net885),
    .B1(net908),
    .X(net5));
 sky130_fd_sc_hd__mux4_1 c670 (.A0(net532),
    .A1(net994),
    .A2(net533),
    .A3(clknet_1_0__leaf_net425),
    .S0(net1016),
    .S1(net1014),
    .X(net534));
 sky130_fd_sc_hd__a21bo_1 c671 (.A1(net533),
    .A2(net994),
    .B1_N(net730),
    .X(net535));
 sky130_fd_sc_hd__mux4_1 c672 (.A0(net530),
    .A1(net531),
    .A2(net533),
    .A3(net1014),
    .S0(net1012),
    .S1(net1021),
    .X(net536));
 sky130_fd_sc_hd__a41o_1 c673 (.A1(net532),
    .A2(net1011),
    .A3(net535),
    .A4(net533),
    .B1(net1014),
    .X(net537));
 sky130_fd_sc_hd__a31o_1 c674 (.A1(net217),
    .A2(net533),
    .A3(net1011),
    .B1(net728),
    .X(net538));
 sky130_fd_sc_hd__mux4_1 c675 (.A0(net430),
    .A1(net530),
    .A2(net1047),
    .A3(net533),
    .S0(net431),
    .S1(net532),
    .X(net539));
 sky130_fd_sc_hd__mux4_1 c676 (.A0(net419),
    .A1(net533),
    .A2(net1014),
    .A3(net728),
    .S0(clknet_1_0__leaf_net742),
    .S1(net1021),
    .X(net540));
 sky130_fd_sc_hd__dlymetal6s2s_1 c677 (.A(net719),
    .X(net541));
 sky130_fd_sc_hd__a41o_1 c678 (.A1(net1011),
    .A2(net696),
    .A3(net728),
    .A4(clknet_1_1__leaf_net742),
    .B1(net1021),
    .X(net542));
 sky130_fd_sc_hd__a21bo_1 c679 (.A1(net529),
    .A2(net535),
    .B1_N(clknet_1_0__leaf_net542),
    .X(net543));
 sky130_fd_sc_hd__a21bo_1 c68 (.A1(net908),
    .A2(net2),
    .B1_N(net1032),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 c680 (.A(net719),
    .X(net544));
 sky130_fd_sc_hd__mux4_1 c681 (.A0(net544),
    .A1(net531),
    .A2(net524),
    .A3(net1014),
    .S0(net1011),
    .S1(clknet_1_0__leaf_net742),
    .X(net545));
 sky130_fd_sc_hd__a41o_1 c682 (.A1(net979),
    .A2(net1015),
    .A3(net1047),
    .A4(net696),
    .B1(clknet_1_0__leaf_net778),
    .X(net546));
 sky130_fd_sc_hd__a31o_2 c683 (.A1(net1015),
    .A2(net1016),
    .A3(net700),
    .B1(net1021),
    .X(net547));
 sky130_fd_sc_hd__a31o_1 c684 (.A1(net524),
    .A2(net896),
    .A3(net547),
    .B1(net1012),
    .X(net548));
 sky130_fd_sc_hd__mux4_1 c685 (.A0(net421),
    .A1(clknet_1_0__leaf_net542),
    .A2(net443),
    .A3(net328),
    .S0(net1045),
    .S1(net842),
    .X(net549));
 sky130_fd_sc_hd__a41o_1 c686 (.A1(net983),
    .A2(net441),
    .A3(net1016),
    .A4(clknet_1_0__leaf_net542),
    .B1(net823),
    .X(net550));
 sky130_fd_sc_hd__mux4_2 c687 (.A0(net530),
    .A1(net1014),
    .A2(net1011),
    .A3(net443),
    .S0(net228),
    .S1(net748),
    .X(net551));
 sky130_fd_sc_hd__a41o_1 c688 (.A1(net1046),
    .A2(net1012),
    .A3(clknet_1_0__leaf_net542),
    .A4(net748),
    .B1(net825),
    .X(net552));
 sky130_fd_sc_hd__a41o_1 c689 (.A1(net543),
    .A2(net443),
    .A3(net983),
    .A4(net979),
    .B1(clknet_1_1__leaf_net742),
    .X(net553));
 sky130_fd_sc_hd__a41o_2 c69 (.A1(net912),
    .A2(net1051),
    .A3(net1037),
    .A4(net900),
    .B1(net1039),
    .X(net7));
 sky130_fd_sc_hd__a41o_2 c690 (.A1(net551),
    .A2(net1016),
    .A3(net1047),
    .A4(net547),
    .B1(net748),
    .X(net554));
 sky130_fd_sc_hd__sdfbbn_2 c691 (.CLK_N(clknet_4_0_0_clk),
    .D(net526),
    .RESET_B(net554),
    .SCD(net876),
    .SCE(net823),
    .SET_B(net825),
    .Q(net556),
    .Q_N(net555));
 sky130_fd_sc_hd__mux4_1 c692 (.A0(net548),
    .A1(net555),
    .A2(net1015),
    .A3(net1016),
    .S0(net983),
    .S1(net653),
    .X(net557));
 sky130_fd_sc_hd__a31o_1 c693 (.A1(net1015),
    .A2(net551),
    .A3(net78),
    .B1(net1012),
    .X(net558));
 sky130_fd_sc_hd__mux4_1 c694 (.A0(clknet_1_0__leaf_net552),
    .A1(net983),
    .A2(net441),
    .A3(net214),
    .S0(net554),
    .S1(net547),
    .X(net559));
 sky130_fd_sc_hd__a41o_1 c695 (.A1(net548),
    .A2(net1012),
    .A3(net983),
    .A4(net653),
    .B1(clknet_1_0__leaf_net742),
    .X(net560));
 sky130_fd_sc_hd__mux4_1 c696 (.A0(net535),
    .A1(net1011),
    .A2(net1015),
    .A3(net983),
    .S0(net551),
    .S1(net753),
    .X(net561));
 sky130_fd_sc_hd__a41o_1 c697 (.A1(clknet_1_0__leaf_net552),
    .A2(net1016),
    .A3(clknet_1_1__leaf_net560),
    .A4(clknet_1_1__leaf_net742),
    .B1(net1021),
    .X(net562));
 sky130_fd_sc_hd__mux4_1 c698 (.A0(net556),
    .A1(net561),
    .A2(net1067),
    .A3(net979),
    .S0(net889),
    .S1(net741),
    .X(net563));
 sky130_fd_sc_hd__a41o_1 c699 (.A1(net443),
    .A2(net441),
    .A3(net555),
    .A4(net228),
    .B1(net1077),
    .X(net564));
 sky130_fd_sc_hd__a21bo_1 c70 (.A1(net888),
    .A2(net3),
    .B1_N(net7),
    .X(net8));
 sky130_fd_sc_hd__a41o_1 c700 (.A1(clknet_1_0__leaf_net562),
    .A2(net979),
    .A3(clknet_1_0__leaf_net560),
    .A4(net653),
    .B1(net1077),
    .X(net565));
 sky130_fd_sc_hd__mux4_1 c701 (.A0(net558),
    .A1(clknet_1_1__leaf_net562),
    .A2(clknet_1_1__leaf_net552),
    .A3(net729),
    .S0(net842),
    .S1(net843),
    .X(net566));
 sky130_fd_sc_hd__mux4_1 c702 (.A0(net228),
    .A1(net979),
    .A2(clknet_1_0__leaf_net562),
    .A3(net524),
    .S0(net729),
    .S1(net844),
    .X(net567));
 sky130_fd_sc_hd__mux4_1 c703 (.A0(clknet_1_0__leaf_net560),
    .A1(net1043),
    .A2(net729),
    .A3(net754),
    .S0(net844),
    .S1(net845),
    .X(net568));
 sky130_fd_sc_hd__mux4_1 c704 (.A0(net554),
    .A1(net557),
    .A2(net981),
    .A3(net556),
    .S0(net983),
    .S1(net824),
    .X(net569));
 sky130_fd_sc_hd__mux4_1 c705 (.A0(net558),
    .A1(net991),
    .A2(net1000),
    .A3(net1043),
    .S0(net983),
    .S1(net754),
    .X(net570));
 sky130_fd_sc_hd__mux4_2 c706 (.A0(net424),
    .A1(net990),
    .A2(net1035),
    .A3(net824),
    .S0(net1021),
    .S1(net846),
    .X(net571));
 sky130_fd_sc_hd__mux4_2 c707 (.A0(net547),
    .A1(net983),
    .A2(clknet_1_1__leaf_net474),
    .A3(net557),
    .S0(net720),
    .S1(net1021),
    .X(net572));
 sky130_fd_sc_hd__mux4_1 c708 (.A0(net561),
    .A1(net1033),
    .A2(net1012),
    .A3(net1016),
    .S0(net832),
    .S1(net847),
    .X(net573));
 sky130_fd_sc_hd__mux4_1 c709 (.A0(clknet_1_0__leaf_net474),
    .A1(net376),
    .A2(net1047),
    .A3(net1021),
    .S0(net848),
    .S1(net849),
    .X(net574));
 sky130_fd_sc_hd__a21bo_1 c71 (.A1(net8),
    .A2(net915),
    .B1_N(net1037),
    .X(net9));
 sky130_fd_sc_hd__mux4_1 c710 (.A0(net557),
    .A1(clknet_1_0__leaf_net568),
    .A2(clknet_1_0__leaf_net474),
    .A3(net1033),
    .S0(net555),
    .S1(net849),
    .X(net575));
 sky130_fd_sc_hd__mux4_1 c711 (.A0(net424),
    .A1(net1002),
    .A2(net981),
    .A3(net653),
    .S0(net832),
    .S1(net849),
    .X(net576));
 sky130_fd_sc_hd__mux4_1 c712 (.A0(net376),
    .A1(net1029),
    .A2(net832),
    .A3(net1021),
    .S0(net842),
    .S1(net845),
    .X(net577));
 sky130_fd_sc_hd__mux4_1 c713 (.A0(net376),
    .A1(net558),
    .A2(net1046),
    .A3(net1041),
    .S0(net824),
    .S1(net851),
    .X(net578));
 sky130_fd_sc_hd__mux4_1 c714 (.A0(net571),
    .A1(net576),
    .A2(net983),
    .A3(net541),
    .S0(net845),
    .S1(net849),
    .X(net579));
 sky130_fd_sc_hd__mux4_1 c715 (.A0(net577),
    .A1(net981),
    .A2(net576),
    .A3(clknet_1_0__leaf_net474),
    .S0(net824),
    .S1(clknet_1_0__leaf_net852),
    .X(net580));
 sky130_fd_sc_hd__mux4_1 c716 (.A0(net561),
    .A1(net988),
    .A2(net1013),
    .A3(net571),
    .S0(net1087),
    .S1(net1072),
    .X(net581));
 sky130_fd_sc_hd__mux4_1 c717 (.A0(net576),
    .A1(net1041),
    .A2(net751),
    .A3(net824),
    .S0(net842),
    .S1(clknet_1_0__leaf_net852),
    .X(net582));
 sky130_fd_sc_hd__mux4_1 c718 (.A0(net554),
    .A1(net571),
    .A2(clknet_1_1__leaf_net568),
    .A3(net842),
    .S0(net847),
    .S1(clknet_1_0__leaf_net852),
    .X(net583));
 sky130_fd_sc_hd__mux4_1 c719 (.A0(clknet_1_1__leaf_net474),
    .A1(net1013),
    .A2(net846),
    .A3(net848),
    .S0(net850),
    .S1(clknet_1_1__leaf_net854),
    .X(net584));
 sky130_fd_sc_hd__a21bo_2 c72 (.A1(net915),
    .A2(net9),
    .B1_N(net8),
    .X(net10));
 sky130_fd_sc_hd__mux4_1 c720 (.A0(net1016),
    .A1(net992),
    .A2(clknet_1_1__leaf_net706),
    .A3(net1029),
    .S0(net849),
    .S1(net851),
    .X(net585));
 sky130_fd_sc_hd__mux4_1 c721 (.A0(net547),
    .A1(net1047),
    .A2(clknet_1_0__leaf_net585),
    .A3(net751),
    .S0(net845),
    .S1(clknet_1_0__leaf_net854),
    .X(net586));
 sky130_fd_sc_hd__mux4_1 c722 (.A0(net1016),
    .A1(clknet_1_1__leaf_net585),
    .A2(net1000),
    .A3(net554),
    .S0(net113),
    .S1(net841),
    .X(net587));
 sky130_fd_sc_hd__mux4_1 c723 (.A0(clknet_1_0__leaf_net568),
    .A1(net586),
    .A2(net547),
    .A3(net751),
    .S0(net842),
    .S1(net851),
    .X(net588));
 sky130_fd_sc_hd__mux4_1 c724 (.A0(clknet_1_0__leaf_net474),
    .A1(net576),
    .A2(net541),
    .A3(net699),
    .S0(net720),
    .S1(clknet_1_1__leaf_net854),
    .X(net589));
 sky130_fd_sc_hd__mux4_1 c725 (.A0(net571),
    .A1(clknet_1_1__leaf_net474),
    .A2(net720),
    .A3(net751),
    .S0(net842),
    .S1(clknet_1_0__leaf_net854),
    .X(net590));
 sky130_fd_sc_hd__mux4_1 c726 (.A0(net237),
    .A1(net1035),
    .A2(net981),
    .A3(net813),
    .S0(net841),
    .S1(clknet_1_1__leaf_net853),
    .X(net591));
 sky130_fd_sc_hd__mux4_1 c727 (.A0(net541),
    .A1(net984),
    .A2(clknet_1_1__leaf_net542),
    .A3(net988),
    .S0(net838),
    .S1(net842),
    .X(net592));
 sky130_fd_sc_hd__mux4_1 c728 (.A0(net237),
    .A1(net1030),
    .A2(net753),
    .A3(net1024),
    .S0(net850),
    .S1(net856),
    .X(net593));
 sky130_fd_sc_hd__mux4_1 c729 (.A0(clknet_1_0__leaf_net592),
    .A1(clknet_1_0__leaf_net386),
    .A2(net328),
    .A3(clknet_1_0__leaf_net483),
    .S0(net753),
    .S1(net856),
    .X(net594));
 sky130_fd_sc_hd__a41o_1 c73 (.A1(net917),
    .A2(net10),
    .A3(net1037),
    .A4(net1032),
    .B1(net133),
    .X(net11));
 sky130_fd_sc_hd__mux4_1 c730 (.A0(clknet_1_1__leaf_net592),
    .A1(net1030),
    .A2(net844),
    .A3(clknet_1_1__leaf_net852),
    .S0(net855),
    .S1(net857),
    .X(net595));
 sky130_fd_sc_hd__mux4_1 c731 (.A0(clknet_1_0__leaf_net483),
    .A1(net984),
    .A2(clknet_1_1__leaf_net386),
    .A3(net394),
    .S0(net556),
    .S1(net1030),
    .X(net596));
 sky130_fd_sc_hd__mux4_1 c732 (.A0(clknet_1_0__leaf_net592),
    .A1(clknet_1_1__leaf_net542),
    .A2(net741),
    .A3(net754),
    .S0(net844),
    .S1(net859),
    .X(net597));
 sky130_fd_sc_hd__mux4_1 c733 (.A0(net597),
    .A1(net556),
    .A2(net455),
    .A3(net997),
    .S0(net832),
    .S1(net856),
    .X(net598));
 sky130_fd_sc_hd__mux4_1 c734 (.A0(clknet_1_0__leaf_net483),
    .A1(net1035),
    .A2(clknet_1_0__leaf_net595),
    .A3(clknet_1_1__leaf_net592),
    .S0(net1024),
    .S1(net1021),
    .X(net599));
 sky130_fd_sc_hd__mux4_1 c735 (.A0(net984),
    .A1(clknet_1_0__leaf_net592),
    .A2(clknet_1_1__leaf_net591),
    .A3(net1046),
    .S0(net715),
    .S1(net859),
    .X(net600));
 sky130_fd_sc_hd__mux4_1 c736 (.A0(net455),
    .A1(net284),
    .A2(net725),
    .A3(net741),
    .S0(net857),
    .S1(net860),
    .X(net601));
 sky130_fd_sc_hd__mux4_1 c737 (.A0(clknet_1_1__leaf_net592),
    .A1(clknet_1_1__leaf_net595),
    .A2(net601),
    .A3(net1013),
    .S0(clknet_1_1__leaf_net542),
    .S1(net697),
    .X(net602));
 sky130_fd_sc_hd__mux4_1 c738 (.A0(clknet_1_0__leaf_net386),
    .A1(clknet_1_0__leaf_net591),
    .A2(net1002),
    .A3(net716),
    .S0(net736),
    .S1(net858),
    .X(net603));
 sky130_fd_sc_hd__mux4_1 c739 (.A0(net541),
    .A1(net725),
    .A2(net736),
    .A3(net842),
    .S0(net844),
    .S1(clknet_1_0__leaf_net853),
    .X(net604));
 sky130_fd_sc_hd__a41o_4 c74 (.A1(net11),
    .A2(net1044),
    .A3(net10),
    .A4(net1037),
    .B1(net1032),
    .X(net12));
 sky130_fd_sc_hd__mux4_1 c740 (.A0(clknet_1_0__leaf_net591),
    .A1(net984),
    .A2(net1045),
    .A3(net751),
    .S0(net832),
    .S1(net858),
    .X(net605));
 sky130_fd_sc_hd__mux4_1 c741 (.A0(net113),
    .A1(clknet_1_0__leaf_net483),
    .A2(clknet_1_1__leaf_net604),
    .A3(clknet_1_1__leaf_net542),
    .S0(net751),
    .S1(clknet_1_1__leaf_net853),
    .X(net606));
 sky130_fd_sc_hd__mux4_1 c742 (.A0(net1033),
    .A1(net284),
    .A2(net981),
    .A3(net715),
    .S0(net751),
    .S1(net837),
    .X(net607));
 sky130_fd_sc_hd__mux4_1 c743 (.A0(clknet_1_1__leaf_net606),
    .A1(net997),
    .A2(net454),
    .A3(net1030),
    .S0(net736),
    .S1(net751),
    .X(net608));
 sky130_fd_sc_hd__mux4_1 c744 (.A0(net1013),
    .A1(clknet_1_0__leaf_net595),
    .A2(net984),
    .A3(clknet_1_0__leaf_net604),
    .S0(net725),
    .S1(net855),
    .X(net609));
 sky130_fd_sc_hd__mux4_1 c745 (.A0(net394),
    .A1(clknet_1_1__leaf_net604),
    .A2(net607),
    .A3(net984),
    .S0(net697),
    .S1(clknet_1_1__leaf_net852),
    .X(net610));
 sky130_fd_sc_hd__mux4_1 c746 (.A0(net593),
    .A1(clknet_1_0__leaf_net604),
    .A2(clknet_1_0__leaf_net386),
    .A3(net724),
    .S0(clknet_1_0__leaf_net853),
    .S1(net855),
    .X(net611));
 sky130_fd_sc_hd__mux4_1 c747 (.A0(net601),
    .A1(clknet_1_0__leaf_net606),
    .A2(clknet_1_1__leaf_net386),
    .A3(net1030),
    .S0(net699),
    .S1(net838),
    .X(net612));
 sky130_fd_sc_hd__mux4_1 c748 (.A0(net601),
    .A1(net1005),
    .A2(net1003),
    .A3(net1033),
    .S0(net716),
    .S1(net741),
    .X(net613));
 sky130_fd_sc_hd__mux4_1 c749 (.A0(net991),
    .A1(net1000),
    .A2(net1046),
    .A3(clknet_1_0__leaf_net798),
    .S0(net840),
    .S1(net850),
    .X(net614));
 sky130_fd_sc_hd__a41o_1 c75 (.A1(net9),
    .A2(net917),
    .A3(net11),
    .A4(net10),
    .B1(net878),
    .X(net13));
 sky130_fd_sc_hd__mux4_1 c750 (.A0(clknet_1_1__leaf_net542),
    .A1(net1000),
    .A2(clknet_1_0__leaf_net510),
    .A3(net993),
    .S0(clknet_1_0__leaf_net798),
    .S1(net840),
    .X(net615));
 sky130_fd_sc_hd__mux4_1 c751 (.A0(net997),
    .A1(clknet_1_0__leaf_net522),
    .A2(net724),
    .A3(net747),
    .S0(net821),
    .S1(net860),
    .X(net616));
 sky130_fd_sc_hd__mux4_2 c752 (.A0(net1048),
    .A1(net614),
    .A2(clknet_1_1__leaf_net522),
    .A3(net747),
    .S0(net846),
    .S1(net860),
    .X(net617));
 sky130_fd_sc_hd__mux4_1 c753 (.A0(clknet_1_1__leaf_net617),
    .A1(net997),
    .A2(clknet_1_0__leaf_net778),
    .A3(net813),
    .S0(net817),
    .S1(net832),
    .X(net618));
 sky130_fd_sc_hd__mux4_2 c754 (.A0(clknet_1_0__leaf_net522),
    .A1(clknet_1_0__leaf_net617),
    .A2(net736),
    .A3(net752),
    .S0(net1024),
    .S1(net850),
    .X(net619));
 sky130_fd_sc_hd__mux4_1 c755 (.A0(net1045),
    .A1(clknet_1_1__leaf_net510),
    .A2(net1048),
    .A3(net716),
    .S0(net752),
    .S1(net844),
    .X(net620));
 sky130_fd_sc_hd__mux4_1 c756 (.A0(clknet_1_0__leaf_net510),
    .A1(clknet_1_1__leaf_net542),
    .A2(clknet_1_1__leaf_net522),
    .A3(net455),
    .S0(net724),
    .S1(clknet_1_0__leaf_net798),
    .X(net621));
 sky130_fd_sc_hd__mux4_1 c757 (.A0(net607),
    .A1(net621),
    .A2(net752),
    .A3(clknet_1_0__leaf_net798),
    .S0(net832),
    .S1(net844),
    .X(net622));
 sky130_fd_sc_hd__mux4_1 c758 (.A0(net1005),
    .A1(net284),
    .A2(clknet_1_1__leaf_net706),
    .A3(clknet_1_0__leaf_net778),
    .S0(net813),
    .S1(net846),
    .X(net623));
 sky130_fd_sc_hd__mux4_1 c759 (.A0(net284),
    .A1(net616),
    .A2(net1033),
    .A3(clknet_1_0__leaf_net483),
    .S0(net741),
    .S1(net842),
    .X(net624));
 sky130_fd_sc_hd__a41o_2 c76 (.A1(net1032),
    .A2(net908),
    .A3(net13),
    .A4(net899),
    .B1(net2),
    .X(net14));
 sky130_fd_sc_hd__mux4_1 c760 (.A0(net993),
    .A1(net697),
    .A2(net736),
    .A3(net747),
    .S0(net813),
    .S1(net840),
    .X(net625));
 sky130_fd_sc_hd__mux4_1 c761 (.A0(net613),
    .A1(net997),
    .A2(net620),
    .A3(net625),
    .S0(net752),
    .S1(net840),
    .X(net626));
 sky130_fd_sc_hd__mux4_1 c762 (.A0(clknet_1_0__leaf_net623),
    .A1(clknet_1_0__leaf_net510),
    .A2(net697),
    .A3(net716),
    .S0(clknet_1_0__leaf_net778),
    .S1(clknet_1_0__leaf_net815),
    .X(net627));
 sky130_fd_sc_hd__mux4_1 c763 (.A0(net626),
    .A1(net627),
    .A2(net736),
    .A3(net741),
    .S0(net832),
    .S1(net837),
    .X(net628));
 sky130_fd_sc_hd__mux4_1 c764 (.A0(clknet_1_1__leaf_net623),
    .A1(net615),
    .A2(net625),
    .A3(net628),
    .S0(net1003),
    .S1(net896),
    .X(net629));
 sky130_fd_sc_hd__a41o_1 c77 (.A1(net9),
    .A2(net11),
    .A3(net878),
    .A4(net873),
    .B1(net8),
    .X(net15));
 sky130_fd_sc_hd__mux4_2 c78 (.A0(net2),
    .A1(net9),
    .A2(net915),
    .A3(net7),
    .S0(net12),
    .S1(net11),
    .X(net16));
 sky130_fd_sc_hd__a21bo_2 c79 (.A1(net904),
    .A2(net13),
    .B1_N(net10),
    .X(net17));
 sky130_fd_sc_hd__a21bo_1 c80 (.A1(net12),
    .A2(net6),
    .B1_N(net10),
    .X(net18));
 sky130_fd_sc_hd__a41o_2 c81 (.A1(net881),
    .A2(net998),
    .A3(net1032),
    .A4(net14),
    .B1(net1039),
    .X(net19));
 sky130_fd_sc_hd__a21bo_1 c82 (.A1(net16),
    .A2(net14),
    .B1_N(net910),
    .X(net20));
 sky130_fd_sc_hd__a21bo_2 c83 (.A1(net15),
    .A2(net8),
    .B1_N(net20),
    .X(net21));
 sky130_fd_sc_hd__a41o_1 c84 (.A1(net21),
    .A2(net16),
    .A3(net14),
    .A4(net998),
    .B1(net8),
    .X(net22));
 sky130_fd_sc_hd__mux4_2 c85 (.A0(net22),
    .A1(net21),
    .A2(net10),
    .A3(net998),
    .S0(net1032),
    .S1(net20),
    .X(net23));
 sky130_fd_sc_hd__mux4_1 c86 (.A0(net18),
    .A1(net22),
    .A2(net23),
    .A3(net21),
    .S0(net1043),
    .S1(net19),
    .X(net24));
 sky130_fd_sc_hd__mux4_1 c87 (.A0(net24),
    .A1(net997),
    .A2(net998),
    .A3(net882),
    .S0(net23),
    .S1(net22),
    .X(net25));
 sky130_fd_sc_hd__a21bo_4 c88 (.A1(net13),
    .A2(net919),
    .B1_N(net133),
    .X(net943));
 sky130_fd_sc_hd__a21bo_1 c89 (.A1(net914),
    .A2(net1032),
    .B1_N(net890),
    .X(net26));
 sky130_fd_sc_hd__a21bo_1 c90 (.A1(net8),
    .A2(net900),
    .B1_N(net872),
    .X(net27));
 sky130_fd_sc_hd__a21bo_1 c91 (.A1(net26),
    .A2(net885),
    .B1_N(net18),
    .X(net28));
 sky130_fd_sc_hd__a21bo_1 c92 (.A1(net25),
    .A2(net22),
    .B1_N(net27),
    .X(net29));
 sky130_fd_sc_hd__a21bo_1 c93 (.A1(net919),
    .A2(net25),
    .B1_N(net28),
    .X(net30));
 sky130_fd_sc_hd__a21bo_2 c94 (.A1(net28),
    .A2(net891),
    .B1_N(net30),
    .X(net31));
 sky130_fd_sc_hd__a21bo_1 c95 (.A1(net873),
    .A2(net29),
    .B1_N(net907),
    .X(net32));
 sky130_fd_sc_hd__buf_1 c96 (.A(net665),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_1 c97 (.A(net665),
    .X(net34));
 sky130_fd_sc_hd__sdfrbp_1 c98 (.CLK(clknet_4_14_0_clk),
    .D(net27),
    .RESET_B(net31),
    .SCD(net30),
    .SCE(net1010),
    .Q(net36),
    .Q_N(net35));
 sky130_fd_sc_hd__a31o_1 c99 (.A1(net910),
    .A2(net1037),
    .A3(net1039),
    .B1(net1009),
    .X(net37));
 sky130_fd_sc_hd__a41o_1 merge765 (.A1(net83),
    .A2(net418),
    .A3(net419),
    .A4(net88),
    .B1(net802),
    .X(net630));
 sky130_fd_sc_hd__mux4_1 merge766 (.A0(net31),
    .A1(net44),
    .A2(net872),
    .A3(net907),
    .S0(clknet_1_0__leaf_net48),
    .S1(net32),
    .X(net631));
 sky130_fd_sc_hd__mux4_1 merge767 (.A0(net419),
    .A1(clknet_1_0__leaf_net425),
    .A2(net982),
    .A3(net1057),
    .S0(net424),
    .S1(net217),
    .X(net632));
 sky130_fd_sc_hd__a41o_1 merge768 (.A1(net29),
    .A2(net31),
    .A3(net28),
    .A4(net16),
    .B1(net25),
    .X(net633));
 sky130_fd_sc_hd__a41o_1 merge769 (.A1(net240),
    .A2(net980),
    .A3(net131),
    .A4(net644),
    .B1(net657),
    .X(net634));
 sky130_fd_sc_hd__a41o_1 merge770 (.A1(net1053),
    .A2(net208),
    .A3(net980),
    .A4(net82),
    .B1(net214),
    .X(net635));
 sky130_fd_sc_hd__a41o_1 merge771 (.A1(net420),
    .A2(net419),
    .A3(net421),
    .A4(net76),
    .B1(net424),
    .X(net636));
 sky130_fd_sc_hd__mux4_1 merge772 (.A0(net211),
    .A1(net320),
    .A2(net990),
    .A3(net74),
    .S0(net420),
    .S1(clknet_1_1__leaf_net425),
    .X(net637));
 sky130_fd_sc_hd__mux4_1 merge773 (.A0(net231),
    .A1(net975),
    .A2(clknet_1_1__leaf_net246),
    .A3(net243),
    .S0(clknet_1_0__leaf_net245),
    .S1(net131),
    .X(net638));
 sky130_fd_sc_hd__mux4_1 merge774 (.A0(clknet_1_0__leaf_net425),
    .A1(net524),
    .A2(net419),
    .A3(net533),
    .S0(net418),
    .S1(net700),
    .X(net639));
 sky130_fd_sc_hd__mux4_1 merge775 (.A0(net418),
    .A1(net982),
    .A2(net1068),
    .A3(net531),
    .S0(net532),
    .S1(net1011),
    .X(net640));
 sky130_fd_sc_hd__xnor2_1 merge776 (.A(net53),
    .B(net59),
    .Y(net641));
 sky130_fd_sc_hd__xnor2_1 merge777 (.A(net176),
    .B(net186),
    .Y(net642));
 sky130_fd_sc_hd__dfrbp_2 merge778 (.CLK(clknet_4_10_0_clk),
    .D(net125),
    .RESET_B(net126),
    .Q(net644),
    .Q_N(net643));
 sky130_fd_sc_hd__xnor2_1 merge779 (.A(net287),
    .B(net304),
    .Y(net645));
 sky130_fd_sc_hd__xnor2_1 merge780 (.A(net509),
    .B(net519),
    .Y(net646));
 sky130_fd_sc_hd__xnor2_1 merge781 (.A(net152),
    .B(net139),
    .Y(net647));
 sky130_fd_sc_hd__dfrbp_1 merge782 (.CLK(clknet_4_2_0_clk),
    .D(net319),
    .RESET_B(net323),
    .Q(net649),
    .Q_N(net648));
 sky130_fd_sc_hd__dfrtn_1 merge783 (.CLK_N(clknet_4_2_0_clk),
    .D(net337),
    .RESET_B(net338),
    .Q(net650));
 sky130_fd_sc_hd__xnor2_1 merge784 (.A(net362),
    .B(net361),
    .Y(net651));
 sky130_fd_sc_hd__xnor2_1 merge785 (.A(net444),
    .B(net456),
    .Y(net652));
 sky130_fd_sc_hd__dfrtp_1 merge786 (.CLK(clknet_4_1_0_clk),
    .D(net553),
    .RESET_B(net559),
    .Q(net653));
 sky130_fd_sc_hd__xnor2_1 merge787 (.A(net109),
    .B(net110),
    .Y(net654));
 sky130_fd_sc_hd__xnor2_1 merge788 (.A(net472),
    .B(net480),
    .Y(net655));
 sky130_fd_sc_hd__xnor2_1 merge789 (.A(net410),
    .B(net411),
    .Y(net656));
 sky130_fd_sc_hd__dfrtp_1 merge790 (.CLK(clknet_4_10_0_clk),
    .D(net227),
    .Q(net233));
 sky130_fd_sc_hd__xnor2_1 merge791 (.A(net527),
    .B(net536),
    .Y(net658));
 sky130_fd_sc_hd__dfrtp_1 merge792 (.CLK(clknet_4_15_0_clk),
    .RESET_B(net305),
    .Q(net306));
 sky130_fd_sc_hd__xnor2_1 merge793 (.A(net437),
    .B(net630),
    .Y(net659));
 sky130_fd_sc_hd__xnor2_1 merge794 (.A(net382),
    .B(net398),
    .Y(net660));
 sky130_fd_sc_hd__dfsbp_1 merge795 (.CLK(clknet_4_9_0_clk),
    .D(net283),
    .SET_B(net271),
    .Q(net662),
    .Q_N(net661));
 sky130_fd_sc_hd__xnor2_2 merge796 (.A(net629),
    .B(net619),
    .Y(net663));
 sky130_fd_sc_hd__xnor2_1 merge797 (.A(net491),
    .B(net494),
    .Y(net664));
 sky130_fd_sc_hd__dfsbp_1 merge798 (.CLK(clknet_4_14_0_clk),
    .D(net47),
    .SET_B(net633),
    .Q(net666),
    .Q_N(net665));
 sky130_fd_sc_hd__dfstp_1 merge799 (.CLK(clknet_4_14_0_clk),
    .D(net163),
    .SET_B(net164),
    .Q(net960));
 sky130_fd_sc_hd__xnor2_1 merge800 (.A(net594),
    .B(net605),
    .Y(net667));
 sky130_fd_sc_hd__dfstp_4 merge801 (.CLK(clknet_4_2_0_clk),
    .D(net218),
    .SET_B(net210),
    .Q(net668));
 sky130_fd_sc_hd__xnor2_4 merge802 (.A(net578),
    .B(net572),
    .Y(net669));
 sky130_fd_sc_hd__xnor2_1 merge803 (.A(net252),
    .B(net256),
    .Y(net670));
 sky130_fd_sc_hd__xnor2_1 merge804 (.A(net460),
    .B(net457),
    .Y(net671));
 sky130_fd_sc_hd__dfstp_1 merge805 (.CLK(clknet_4_3_0_clk),
    .D(net374),
    .SET_B(net638),
    .Q(net672));
 sky130_fd_sc_hd__dlrbn_2 merge806 (.D(net216),
    .GATE_N(clknet_4_8_0_clk),
    .RESET_B(net236),
    .Q(net674),
    .Q_N(net673));
 sky130_fd_sc_hd__dlrbn_1 merge807 (.D(net354),
    .GATE_N(clknet_4_2_0_clk),
    .RESET_B(net635),
    .Q(net676),
    .Q_N(net675));
 sky130_fd_sc_hd__xnor2_2 merge808 (.A(net413),
    .B(net417),
    .Y(net677));
 sky130_fd_sc_hd__xnor2_1 merge809 (.A(net482),
    .B(net520),
    .Y(net678));
 sky130_fd_sc_hd__xnor2_1 merge810 (.A(net142),
    .B(net143),
    .Y(net679));
 sky130_fd_sc_hd__dlrbp_1 merge811 (.D(net151),
    .GATE(clknet_4_14_0_clk),
    .RESET_B(net154),
    .Q(net681),
    .Q_N(net680));
 sky130_fd_sc_hd__dlrbp_1 merge812 (.D(net664),
    .GATE(clknet_4_7_0_clk),
    .RESET_B(net502),
    .Q(net683),
    .Q_N(net682));
 sky130_fd_sc_hd__dlrtn_1 merge813 (.D(net352),
    .GATE_N(clknet_4_3_0_clk),
    .RESET_B(net655),
    .Q(net684));
 sky130_fd_sc_hd__dlrtn_1 merge814 (.D(net652),
    .GATE_N(clknet_4_3_0_clk),
    .RESET_B(net449),
    .Q(net685));
 sky130_fd_sc_hd__xnor2_1 merge815 (.A(net584),
    .B(net622),
    .Y(net686));
 sky130_fd_sc_hd__xnor2_1 merge816 (.A(net663),
    .B(net646),
    .Y(net687));
 sky130_fd_sc_hd__xnor2_1 merge817 (.A(net588),
    .B(net611),
    .Y(net688));
 sky130_fd_sc_hd__xnor2_1 merge818 (.A(net416),
    .B(net290),
    .Y(net689));
 sky130_fd_sc_hd__xnor2_1 merge819 (.A(net642),
    .B(net63),
    .Y(net690));
 sky130_fd_sc_hd__xnor2_1 merge820 (.A(net387),
    .B(net293),
    .Y(net691));
 sky130_fd_sc_hd__xnor2_1 merge821 (.A(net609),
    .B(net598),
    .Y(net692));
 sky130_fd_sc_hd__xnor2_1 merge822 (.A(net193),
    .B(net631),
    .Y(net693));
 sky130_fd_sc_hd__xnor2_1 merge823 (.A(net589),
    .B(net570),
    .Y(net694));
 sky130_fd_sc_hd__xnor2_1 merge824 (.A(net167),
    .B(net150),
    .Y(net695));
 sky130_fd_sc_hd__dlrtn_1 merge825 (.D(net632),
    .GATE_N(clknet_4_0_0_clk),
    .RESET_B(net658),
    .Q(net696));
 sky130_fd_sc_hd__dlrtp_1 merge826 (.D(net600),
    .GATE(clknet_4_5_0_clk),
    .RESET_B(net624),
    .Q(net697));
 sky130_fd_sc_hd__dlrtp_1 merge827 (.D(net654),
    .GATE(clknet_4_10_0_clk),
    .RESET_B(net111),
    .Q(net698));
 sky130_fd_sc_hd__dlrtp_2 merge828 (.D(net370),
    .GATE(clknet_4_12_0_clk),
    .RESET_B(net677),
    .Q(net953));
 sky130_fd_sc_hd__edfxbp_1 merge829 (.CLK(clknet_4_0_0_clk),
    .D(net538),
    .DE(net688),
    .Q(net700),
    .Q_N(net699));
 sky130_fd_sc_hd__xnor2_1 merge830 (.A(net660),
    .B(net656),
    .Y(net701));
 sky130_fd_sc_hd__edfxtp_1 merge831 (.CLK(clknet_4_15_0_clk),
    .D(net41),
    .DE(net195),
    .Q(net702));
 sky130_fd_sc_hd__xnor2_1 merge832 (.A(net258),
    .B(net299),
    .Y(net703));
 sky130_fd_sc_hd__xnor2_1 merge833 (.A(net634),
    .B(net388),
    .Y(net704));
 sky130_fd_sc_hd__sdlclkp_1 merge834 (.CLK(clknet_4_13_0_clk),
    .GATE(net406),
    .SCE(net402),
    .GCLK(net945));
 sky130_fd_sc_hd__sdlclkp_2 merge835 (.CLK(clknet_4_14_0_clk),
    .GATE(net645),
    .SCE(net647),
    .GCLK(net705));
 sky130_fd_sc_hd__sdlclkp_4 merge836 (.CLK(clknet_4_0_0_clk),
    .GATE(net636),
    .SCE(net686),
    .GCLK(net706));
 sky130_fd_sc_hd__xnor2_1 merge837 (.A(net670),
    .B(net260),
    .Y(net707));
 sky130_fd_sc_hd__dfrbp_1 merge838 (.CLK(clknet_4_11_0_clk),
    .D(net132),
    .Q(net709),
    .Q_N(net708));
 sky130_fd_sc_hd__xnor2_1 merge839 (.A(net379),
    .B(net385),
    .Y(net710));
 sky130_fd_sc_hd__xnor2_1 merge840 (.A(net651),
    .B(net669),
    .Y(net711));
 sky130_fd_sc_hd__xnor2_1 merge841 (.A(net383),
    .B(net384),
    .Y(net712));
 sky130_fd_sc_hd__dfrbp_1 merge842 (.CLK(clknet_4_3_0_clk),
    .D(net313),
    .RESET_B(net367),
    .Q(net714),
    .Q_N(net713));
 sky130_fd_sc_hd__dfrtn_1 merge843 (.CLK_N(clknet_4_4_0_clk),
    .D(net667),
    .RESET_B(net468),
    .Q(net715));
 sky130_fd_sc_hd__dfrtp_4 merge844 (.CLK(clknet_4_5_0_clk),
    .D(net687),
    .RESET_B(net596),
    .Q(net716));
 sky130_fd_sc_hd__dfrtp_2 merge845 (.CLK(clknet_4_4_0_clk),
    .D(net678),
    .RESET_B(net476),
    .Q(net717));
 sky130_fd_sc_hd__xnor2_1 merge846 (.A(net637),
    .B(net477),
    .Y(net718));
 sky130_fd_sc_hd__dfrtp_1 merge847 (.CLK(clknet_4_0_0_clk),
    .D(net640),
    .RESET_B(net639),
    .Q(net719));
 sky130_fd_sc_hd__dfsbp_1 merge848 (.CLK(clknet_4_4_0_clk),
    .D(net488),
    .SET_B(net694),
    .Q(net721),
    .Q_N(net720));
 sky130_fd_sc_hd__dfsbp_2 merge849 (.CLK(clknet_4_0_0_clk),
    .D(net432),
    .SET_B(net518),
    .Q(net723),
    .Q_N(net722));
 sky130_fd_sc_hd__dfstp_2 merge850 (.CLK(clknet_4_5_0_clk),
    .D(net692),
    .SET_B(net479),
    .Q(net724));
 sky130_fd_sc_hd__dfstp_2 merge851 (.CLK(clknet_4_5_0_clk),
    .D(net689),
    .SET_B(net599),
    .Q(net725));
 sky130_fd_sc_hd__dfstp_2 merge852 (.CLK(clknet_4_2_0_clk),
    .D(net427),
    .SET_B(net671),
    .Q(net726));
 sky130_fd_sc_hd__dlrbn_2 merge853 (.D(net537),
    .GATE_N(clknet_4_0_0_clk),
    .RESET_B(net279),
    .Q(net728),
    .Q_N(net727));
 sky130_fd_sc_hd__dlrbn_1 merge854 (.D(net436),
    .GATE_N(clknet_4_0_0_clk),
    .RESET_B(net565),
    .Q(net730),
    .Q_N(net729));
 sky130_fd_sc_hd__dlrbp_1 merge855 (.D(net178),
    .GATE(clknet_4_7_0_clk),
    .RESET_B(net489),
    .Q(net732),
    .Q_N(net731));
 sky130_fd_sc_hd__dlrbp_1 merge856 (.D(net703),
    .GATE(clknet_4_12_0_clk),
    .RESET_B(net278),
    .Q(net734),
    .Q_N(net733));
 sky130_fd_sc_hd__dlrtn_1 merge857 (.D(net414),
    .GATE_N(clknet_4_13_0_clk),
    .RESET_B(net405),
    .Q(net735));
 sky130_fd_sc_hd__dlrtn_2 merge858 (.D(net612),
    .GATE_N(clknet_4_5_0_clk),
    .RESET_B(net602),
    .Q(net736));
 sky130_fd_sc_hd__dlrtn_2 merge859 (.D(net695),
    .GATE_N(clknet_4_12_0_clk),
    .RESET_B(net294),
    .Q(net961));
 sky130_fd_sc_hd__dlrtp_1 merge860 (.D(net189),
    .GATE(clknet_4_15_0_clk),
    .RESET_B(net641),
    .Q(net949));
 sky130_fd_sc_hd__dlrtp_2 merge861 (.D(net659),
    .GATE(clknet_4_2_0_clk),
    .RESET_B(net718),
    .Q(net737));
 sky130_fd_sc_hd__dlrtp_2 merge862 (.D(net704),
    .GATE(clknet_4_9_0_clk),
    .RESET_B(net710),
    .Q(net738));
 sky130_fd_sc_hd__edfxbp_1 merge863 (.CLK(clknet_4_11_0_clk),
    .DE(net263),
    .Q(net740),
    .Q_N(net266));
 sky130_fd_sc_hd__edfxtp_1 merge864 (.CLK(clknet_4_4_0_clk),
    .D(net546),
    .DE(net610),
    .Q(net741));
 sky130_fd_sc_hd__sdlclkp_1 merge865 (.CLK(clknet_4_0_0_clk),
    .GATE(net539),
    .SCE(net550),
    .GCLK(net742));
 sky130_fd_sc_hd__sdlclkp_2 merge866 (.CLK(clknet_4_14_0_clk),
    .GATE(net148),
    .SCE(net693),
    .GCLK(net743));
 sky130_fd_sc_hd__sdlclkp_4 merge867 (.CLK(clknet_4_14_0_clk),
    .GATE(net679),
    .SCE(net690),
    .GCLK(net744));
 sky130_fd_sc_hd__dfrbp_2 merge868 (.CLK(clknet_4_9_0_clk),
    .D(net269),
    .RESET_B(net291),
    .Q(net746),
    .Q_N(net745));
 sky130_fd_sc_hd__dfrbp_1 merge869 (.CLK(clknet_4_1_0_clk),
    .D(net549),
    .RESET_B(net608),
    .Q(net748),
    .Q_N(net747));
 sky130_fd_sc_hd__dfrtn_1 merge870 (.CLK_N(clknet_4_14_0_clk),
    .D(net711),
    .RESET_B(net180),
    .Q(net749));
 sky130_fd_sc_hd__dfrtp_1 merge871 (.CLK(clknet_4_10_0_clk),
    .D(net114),
    .RESET_B(net707),
    .Q(net750));
 sky130_fd_sc_hd__dfrtp_4 merge872 (.CLK(clknet_4_12_0_clk),
    .D(net691),
    .RESET_B(net701),
    .Q(net962));
 sky130_fd_sc_hd__dfrtp_4 merge873 (.CLK(clknet_4_4_0_clk),
    .D(net603),
    .RESET_B(net581),
    .Q(net751));
 sky130_fd_sc_hd__dfsbp_2 merge874 (.CLK(clknet_4_5_0_clk),
    .D(net712),
    .SET_B(net618),
    .Q(net955),
    .Q_N(net752));
 sky130_fd_sc_hd__dfsbp_1 merge875 (.CLK(clknet_4_0_0_clk),
    .D(net564),
    .SET_B(net540),
    .Q(net754),
    .Q_N(net753));
 sky130_fd_sc_hd__dfxbp_1 s876 (.CLK(clknet_4_14_0_clk),
    .D(net43),
    .Q(net756),
    .Q_N(net755));
 sky130_fd_sc_hd__dfxbp_2 s877 (.CLK(clknet_4_10_0_clk),
    .D(net108),
    .Q(net758),
    .Q_N(net757));
 sky130_fd_sc_hd__dfxtp_2 s878 (.CLK(clknet_4_11_0_clk),
    .D(net120),
    .Q(net963));
 sky130_fd_sc_hd__dfxtp_2 s879 (.CLK(clknet_4_14_0_clk),
    .D(net144),
    .Q(net759));
 sky130_fd_sc_hd__dfxtp_4 s880 (.CLK(clknet_4_11_0_clk),
    .D(net155),
    .Q(net966));
 sky130_fd_sc_hd__dlclkp_1 s881 (.CLK(clknet_4_11_0_clk),
    .GATE(net156),
    .GCLK(net760));
 sky130_fd_sc_hd__dlclkp_2 s882 (.CLK(clknet_4_14_0_clk),
    .GATE(net157),
    .GCLK(net761));
 sky130_fd_sc_hd__dlclkp_4 s883 (.CLK(clknet_4_14_0_clk),
    .GATE(net158),
    .GCLK(net762));
 sky130_fd_sc_hd__dlxbn_1 s884 (.D(net159),
    .GATE_N(clknet_4_15_0_clk),
    .Q(net764),
    .Q_N(net763));
 sky130_fd_sc_hd__dlxbn_2 s885 (.D(net160),
    .GATE_N(clknet_4_15_0_clk),
    .Q(net929),
    .Q_N(net765));
 sky130_fd_sc_hd__dlxbp_1 s886 (.D(net161),
    .GATE(clknet_4_15_0_clk),
    .Q(net767),
    .Q_N(net766));
 sky130_fd_sc_hd__dlxtn_2 s887 (.D(net162),
    .GATE_N(clknet_4_15_0_clk),
    .Q(net768));
 sky130_fd_sc_hd__dlxtn_2 s888 (.D(net165),
    .GATE_N(clknet_4_13_0_clk),
    .Q(net769));
 sky130_fd_sc_hd__dlxtn_2 s889 (.D(net166),
    .GATE_N(clknet_4_13_0_clk),
    .Q(net770));
 sky130_fd_sc_hd__dlxtp_1 s890 (.D(net170),
    .GATE(clknet_4_13_0_clk),
    .Q(net771));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s891 (.D(net173),
    .SLEEP_B(clknet_4_13_0_clk),
    .Q(net772));
 sky130_fd_sc_hd__dfxbp_1 s892 (.CLK(clknet_4_15_0_clk),
    .D(net183),
    .Q(net956),
    .Q_N(net773));
 sky130_fd_sc_hd__dfxbp_1 s893 (.CLK(clknet_4_15_0_clk),
    .D(net187),
    .Q(net775),
    .Q_N(net774));
 sky130_fd_sc_hd__dfxtp_1 s894 (.CLK(clknet_4_15_0_clk),
    .D(net190),
    .Q(net776));
 sky130_fd_sc_hd__dfxtp_2 s895 (.CLK(clknet_4_8_0_clk),
    .D(net219),
    .Q(net777));
 sky130_fd_sc_hd__dfxtp_2 s896 (.CLK(clknet_4_8_0_clk),
    .D(net226),
    .Q(net923));
 sky130_fd_sc_hd__dlclkp_1 s897 (.CLK(clknet_4_8_0_clk),
    .GATE(net235),
    .GCLK(net778));
 sky130_fd_sc_hd__dlclkp_2 s898 (.CLK(clknet_4_8_0_clk),
    .GATE(net239),
    .GCLK(net779));
 sky130_fd_sc_hd__dlclkp_4 s899 (.CLK(clknet_4_10_0_clk),
    .GATE(net244),
    .GCLK(net780));
 sky130_fd_sc_hd__dlxbn_2 s900 (.D(net248),
    .GATE_N(clknet_4_9_0_clk),
    .Q(net782),
    .Q_N(net781));
 sky130_fd_sc_hd__dlxbn_2 s901 (.D(net259),
    .GATE_N(clknet_4_8_0_clk),
    .Q(net976),
    .Q_N(net783));
 sky130_fd_sc_hd__dlxbp_1 s902 (.D(net262),
    .GATE(clknet_4_8_0_clk),
    .Q(net785),
    .Q_N(net784));
 sky130_fd_sc_hd__dlxtn_2 s903 (.D(net264),
    .GATE_N(clknet_4_9_0_clk),
    .Q(net786));
 sky130_fd_sc_hd__dlxtn_2 s904 (.D(net265),
    .GATE_N(clknet_4_9_0_clk),
    .Q(net787));
 sky130_fd_sc_hd__dlxtn_1 s905 (.D(net267),
    .GATE_N(clknet_4_11_0_clk),
    .Q(net788));
 sky130_fd_sc_hd__dlxtp_1 s906 (.D(net268),
    .GATE(clknet_4_9_0_clk),
    .Q(net789));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s907 (.D(net270),
    .SLEEP_B(clknet_4_9_0_clk),
    .Q(net790));
 sky130_fd_sc_hd__dfxbp_1 s908 (.CLK(clknet_4_9_0_clk),
    .D(net274),
    .Q(net970),
    .Q_N(net791));
 sky130_fd_sc_hd__dfxbp_1 s909 (.CLK(clknet_4_6_0_clk),
    .D(net276),
    .Q(net793),
    .Q_N(net792));
 sky130_fd_sc_hd__dfxtp_1 s910 (.CLK(clknet_4_12_0_clk),
    .D(net277),
    .Q(net794));
 sky130_fd_sc_hd__dfxtp_2 s911 (.CLK(clknet_4_9_0_clk),
    .D(net280),
    .Q(net795));
 sky130_fd_sc_hd__dfxtp_2 s912 (.CLK(clknet_4_13_0_clk),
    .D(net286),
    .Q(net796));
 sky130_fd_sc_hd__dlclkp_1 s913 (.CLK(clknet_4_13_0_clk),
    .GATE(net298),
    .GCLK(net797));
 sky130_fd_sc_hd__dlclkp_2 s914 (.CLK(clknet_4_12_0_clk),
    .GATE(net301),
    .GCLK(net798));
 sky130_fd_sc_hd__dlclkp_4 s915 (.CLK(clknet_4_2_0_clk),
    .GATE(net325),
    .GCLK(net799));
 sky130_fd_sc_hd__dlxbn_2 s916 (.D(net326),
    .GATE_N(clknet_4_2_0_clk),
    .Q(net801),
    .Q_N(net800));
 sky130_fd_sc_hd__dlxbn_1 s917 (.D(net327),
    .GATE_N(clknet_4_2_0_clk),
    .Q(net803),
    .Q_N(net802));
 sky130_fd_sc_hd__dlxbp_1 s918 (.D(net336),
    .GATE(clknet_4_3_0_clk),
    .Q(net805),
    .Q_N(net804));
 sky130_fd_sc_hd__dlxtn_2 s919 (.D(net349),
    .GATE_N(clknet_4_2_0_clk),
    .Q(net806));
 sky130_fd_sc_hd__dlxtn_2 s920 (.D(net350),
    .GATE_N(clknet_4_3_0_clk),
    .Q(net939));
 sky130_fd_sc_hd__dlxtn_2 s921 (.D(net353),
    .GATE_N(clknet_4_3_0_clk),
    .Q(net807));
 sky130_fd_sc_hd__dlxtp_1 s922 (.D(net355),
    .GATE(clknet_4_6_0_clk),
    .Q(net808));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s923 (.D(net380),
    .SLEEP_B(clknet_4_6_0_clk),
    .Q(net951));
 sky130_fd_sc_hd__dfxbp_1 s924 (.CLK(clknet_4_6_0_clk),
    .D(net381),
    .Q(net810),
    .Q_N(net809));
 sky130_fd_sc_hd__dfxbp_1 s925 (.CLK(clknet_4_9_0_clk),
    .D(net389),
    .Q(net812),
    .Q_N(net811));
 sky130_fd_sc_hd__dfxtp_4 s926 (.CLK(clknet_4_12_0_clk),
    .D(net392),
    .Q(net978));
 sky130_fd_sc_hd__dfxtp_2 s927 (.CLK(clknet_4_6_0_clk),
    .D(net395),
    .Q(net813));
 sky130_fd_sc_hd__dfxtp_2 s928 (.CLK(clknet_4_12_0_clk),
    .D(net399),
    .Q(net814));
 sky130_fd_sc_hd__dlclkp_1 s929 (.CLK(clknet_4_12_0_clk),
    .GATE(net404),
    .GCLK(net927));
 sky130_fd_sc_hd__dlclkp_2 s930 (.CLK(clknet_4_7_0_clk),
    .GATE(net407),
    .GCLK(net815));
 sky130_fd_sc_hd__dlclkp_4 s931 (.CLK(clknet_4_13_0_clk),
    .GATE(net408),
    .GCLK(net924));
 sky130_fd_sc_hd__dlxbn_1 s932 (.D(net409),
    .GATE_N(clknet_4_7_0_clk),
    .Q(net817),
    .Q_N(net816));
 sky130_fd_sc_hd__dlxbn_1 s933 (.D(net412),
    .GATE_N(clknet_4_13_0_clk),
    .Q(net819),
    .Q_N(net818));
 sky130_fd_sc_hd__dlxbp_1 s934 (.D(net415),
    .GATE(clknet_4_13_0_clk),
    .Q(net821),
    .Q_N(net820));
 sky130_fd_sc_hd__dlxtn_2 s935 (.D(net434),
    .GATE_N(clknet_4_0_0_clk),
    .Q(net822));
 sky130_fd_sc_hd__dlxtn_1 s936 (.D(net435),
    .GATE_N(clknet_4_0_0_clk),
    .Q(net823));
 sky130_fd_sc_hd__dlxtn_2 s937 (.D(net438),
    .GATE_N(clknet_4_1_0_clk),
    .Q(net824));
 sky130_fd_sc_hd__dlxtp_1 s938 (.D(net458),
    .GATE(clknet_4_0_0_clk),
    .Q(net825));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s939 (.D(net459),
    .SLEEP_B(clknet_4_1_0_clk),
    .Q(net936));
 sky130_fd_sc_hd__dfxbp_2 s940 (.CLK(clknet_4_6_0_clk),
    .D(net463),
    .Q(net827),
    .Q_N(net826));
 sky130_fd_sc_hd__dfxbp_1 s941 (.CLK(clknet_4_1_0_clk),
    .D(net466),
    .Q(net829),
    .Q_N(net828));
 sky130_fd_sc_hd__dfxtp_1 s942 (.CLK(clknet_4_1_0_clk),
    .D(net470),
    .Q(net830));
 sky130_fd_sc_hd__dfxtp_2 s943 (.CLK(clknet_4_6_0_clk),
    .D(net473),
    .Q(net831));
 sky130_fd_sc_hd__dfxtp_4 s944 (.CLK(clknet_4_4_0_clk),
    .D(net478),
    .Q(net832));
 sky130_fd_sc_hd__dlclkp_1 s945 (.CLK(clknet_4_7_0_clk),
    .GATE(net495),
    .GCLK(net833));
 sky130_fd_sc_hd__dlclkp_2 s946 (.CLK(clknet_4_7_0_clk),
    .GATE(net496),
    .GCLK(net834));
 sky130_fd_sc_hd__dlclkp_4 s947 (.CLK(clknet_4_7_0_clk),
    .GATE(net497),
    .GCLK(net835));
 sky130_fd_sc_hd__dlxbn_2 s948 (.D(net501),
    .GATE_N(clknet_4_5_0_clk),
    .Q(net933),
    .Q_N(net836));
 sky130_fd_sc_hd__dlxbn_2 s949 (.D(net503),
    .GATE_N(clknet_4_5_0_clk),
    .Q(net838),
    .Q_N(net837));
 sky130_fd_sc_hd__dlxbp_1 s950 (.D(net504),
    .GATE(clknet_4_7_0_clk),
    .Q(net944),
    .Q_N(net839));
 sky130_fd_sc_hd__dlxtn_1 s951 (.D(net523),
    .GATE_N(clknet_4_5_0_clk),
    .Q(net840));
 sky130_fd_sc_hd__dlxtn_1 s952 (.D(net534),
    .GATE_N(clknet_4_0_0_clk),
    .Q(net841));
 sky130_fd_sc_hd__dlxtn_4 s953 (.D(net545),
    .GATE_N(clknet_4_0_0_clk),
    .Q(net842));
 sky130_fd_sc_hd__dlxtp_1 s954 (.D(net563),
    .GATE(clknet_4_1_0_clk),
    .Q(net843));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s955 (.D(net566),
    .SLEEP_B(clknet_4_1_0_clk),
    .Q(net844));
 sky130_fd_sc_hd__dfxbp_1 s956 (.CLK(clknet_4_1_0_clk),
    .D(net567),
    .Q(net846),
    .Q_N(net845));
 sky130_fd_sc_hd__dfxbp_1 s957 (.CLK(clknet_4_1_0_clk),
    .D(net569),
    .Q(net848),
    .Q_N(net847));
 sky130_fd_sc_hd__dfxtp_2 s958 (.CLK(clknet_4_1_0_clk),
    .D(net573),
    .Q(net849));
 sky130_fd_sc_hd__dfxtp_1 s959 (.CLK(clknet_4_4_0_clk),
    .D(net574),
    .Q(net850));
 sky130_fd_sc_hd__dfxtp_1 s960 (.CLK(clknet_4_1_0_clk),
    .D(net575),
    .Q(net851));
 sky130_fd_sc_hd__dlclkp_1 s961 (.CLK(clknet_4_4_0_clk),
    .GATE(net579),
    .GCLK(net852));
 sky130_fd_sc_hd__dlclkp_2 s962 (.CLK(clknet_4_4_0_clk),
    .GATE(net580),
    .GCLK(net853));
 sky130_fd_sc_hd__dlclkp_4 s963 (.CLK(clknet_4_4_0_clk),
    .GATE(net582),
    .GCLK(net854));
 sky130_fd_sc_hd__dlxbn_1 s964 (.D(net583),
    .GATE_N(clknet_4_4_0_clk),
    .Q(net856),
    .Q_N(net855));
 sky130_fd_sc_hd__dlxbn_1 s965 (.D(net587),
    .GATE_N(clknet_4_4_0_clk),
    .Q(net858),
    .Q_N(net857));
 sky130_fd_sc_hd__dlxbp_1 s966 (.D(net590),
    .GATE(clknet_4_4_0_clk),
    .Q(net860),
    .Q_N(net859));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Right_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Right_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Right_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Right_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Right_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Right_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Right_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Right_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Right_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Right_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Right_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Right_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Right_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Right_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Right_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Right_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Right_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Right_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Right_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Right_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Right_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_161 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_162 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_163 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_164 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_165 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_166 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_167 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_168 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_169 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_170 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_171 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_172 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_173 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_174 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_175 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_176 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_177 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_178 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_179 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_180 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_181 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_182 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Left_183 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Left_184 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Left_185 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Left_186 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Left_187 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Left_188 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Left_189 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Left_190 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Left_191 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Left_192 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Left_193 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Left_194 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Left_195 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Left_196 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Left_197 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Left_198 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Left_199 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Left_200 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Left_201 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Left_202 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Left_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1347 ();
 sky130_fd_sc_hd__buf_12 input1 (.A(in0),
    .X(net133));
 sky130_fd_sc_hd__clkbuf_2 input2 (.A(in1),
    .X(net861));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(in10),
    .X(net862));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(in11),
    .X(net863));
 sky130_fd_sc_hd__buf_1 input5 (.A(in12),
    .X(net864));
 sky130_fd_sc_hd__clkbuf_4 input6 (.A(in13),
    .X(net865));
 sky130_fd_sc_hd__clkbuf_4 input7 (.A(in14),
    .X(net866));
 sky130_fd_sc_hd__buf_1 input8 (.A(in15),
    .X(net867));
 sky130_fd_sc_hd__dlymetal6s2s_1 input9 (.A(in16),
    .X(net868));
 sky130_fd_sc_hd__buf_1 input10 (.A(in17),
    .X(net869));
 sky130_fd_sc_hd__buf_1 input11 (.A(in18),
    .X(net870));
 sky130_fd_sc_hd__buf_1 input12 (.A(in19),
    .X(net871));
 sky130_fd_sc_hd__clkbuf_4 input13 (.A(in2),
    .X(net872));
 sky130_fd_sc_hd__buf_1 input14 (.A(in20),
    .X(net873));
 sky130_fd_sc_hd__buf_1 input15 (.A(in21),
    .X(net874));
 sky130_fd_sc_hd__buf_1 input16 (.A(in22),
    .X(net875));
 sky130_fd_sc_hd__buf_2 input17 (.A(in23),
    .X(net876));
 sky130_fd_sc_hd__dlymetal6s2s_1 input18 (.A(in24),
    .X(net877));
 sky130_fd_sc_hd__clkbuf_4 input19 (.A(in25),
    .X(net878));
 sky130_fd_sc_hd__buf_2 input20 (.A(in26),
    .X(net879));
 sky130_fd_sc_hd__buf_2 input21 (.A(in27),
    .X(net880));
 sky130_fd_sc_hd__clkbuf_1 input22 (.A(in28),
    .X(net881));
 sky130_fd_sc_hd__buf_4 input23 (.A(in29),
    .X(net882));
 sky130_fd_sc_hd__buf_1 input24 (.A(in3),
    .X(net883));
 sky130_fd_sc_hd__buf_1 input25 (.A(in30),
    .X(net884));
 sky130_fd_sc_hd__clkbuf_4 input26 (.A(in31),
    .X(net885));
 sky130_fd_sc_hd__buf_1 input27 (.A(in32),
    .X(net886));
 sky130_fd_sc_hd__buf_1 input28 (.A(in33),
    .X(net887));
 sky130_fd_sc_hd__clkbuf_1 input29 (.A(in34),
    .X(net888));
 sky130_fd_sc_hd__buf_4 input30 (.A(in35),
    .X(net889));
 sky130_fd_sc_hd__buf_1 input31 (.A(in36),
    .X(net890));
 sky130_fd_sc_hd__buf_2 input32 (.A(in37),
    .X(net891));
 sky130_fd_sc_hd__buf_1 input33 (.A(in38),
    .X(net892));
 sky130_fd_sc_hd__dlymetal6s2s_1 input34 (.A(in39),
    .X(net893));
 sky130_fd_sc_hd__clkbuf_2 input35 (.A(in4),
    .X(net894));
 sky130_fd_sc_hd__buf_1 input36 (.A(in40),
    .X(net895));
 sky130_fd_sc_hd__buf_4 input37 (.A(in41),
    .X(net896));
 sky130_fd_sc_hd__dlymetal6s2s_1 input38 (.A(in42),
    .X(net897));
 sky130_fd_sc_hd__clkbuf_1 input39 (.A(in43),
    .X(net898));
 sky130_fd_sc_hd__buf_1 input40 (.A(in44),
    .X(net899));
 sky130_fd_sc_hd__clkbuf_2 input41 (.A(in45),
    .X(net900));
 sky130_fd_sc_hd__clkbuf_1 input42 (.A(in46),
    .X(net901));
 sky130_fd_sc_hd__buf_1 input43 (.A(in47),
    .X(net902));
 sky130_fd_sc_hd__buf_1 input44 (.A(in48),
    .X(net903));
 sky130_fd_sc_hd__clkbuf_1 input45 (.A(in49),
    .X(net904));
 sky130_fd_sc_hd__buf_1 input46 (.A(in5),
    .X(net905));
 sky130_fd_sc_hd__clkbuf_2 input47 (.A(in50),
    .X(net906));
 sky130_fd_sc_hd__buf_1 input48 (.A(in51),
    .X(net907));
 sky130_fd_sc_hd__buf_4 input49 (.A(in52),
    .X(net908));
 sky130_fd_sc_hd__clkbuf_2 input50 (.A(in53),
    .X(net909));
 sky130_fd_sc_hd__buf_1 input51 (.A(in54),
    .X(net910));
 sky130_fd_sc_hd__buf_1 input52 (.A(in55),
    .X(net911));
 sky130_fd_sc_hd__buf_1 input53 (.A(in56),
    .X(net912));
 sky130_fd_sc_hd__clkbuf_4 input54 (.A(in57),
    .X(net913));
 sky130_fd_sc_hd__buf_1 input55 (.A(in58),
    .X(net914));
 sky130_fd_sc_hd__dlymetal6s2s_1 input56 (.A(in59),
    .X(net915));
 sky130_fd_sc_hd__buf_1 input57 (.A(in6),
    .X(net916));
 sky130_fd_sc_hd__buf_1 input58 (.A(in60),
    .X(net917));
 sky130_fd_sc_hd__buf_1 input59 (.A(in61),
    .X(net918));
 sky130_fd_sc_hd__buf_1 input60 (.A(in7),
    .X(net919));
 sky130_fd_sc_hd__clkbuf_2 input61 (.A(in8),
    .X(net920));
 sky130_fd_sc_hd__buf_1 input62 (.A(in9),
    .X(net921));
 sky130_fd_sc_hd__clkbuf_1 output63 (.A(clknet_1_1__leaf_net922),
    .X(out0));
 sky130_fd_sc_hd__buf_2 output64 (.A(net1026),
    .X(out1));
 sky130_fd_sc_hd__clkbuf_1 output65 (.A(clknet_1_1__leaf_net924),
    .X(out10));
 sky130_fd_sc_hd__buf_2 output66 (.A(net925),
    .X(out11));
 sky130_fd_sc_hd__buf_2 output67 (.A(net926),
    .X(out12));
 sky130_fd_sc_hd__clkbuf_1 output68 (.A(clknet_1_1__leaf_net927),
    .X(out13));
 sky130_fd_sc_hd__buf_2 output69 (.A(net928),
    .X(out14));
 sky130_fd_sc_hd__buf_2 output70 (.A(net929),
    .X(out15));
 sky130_fd_sc_hd__buf_2 output71 (.A(net930),
    .X(out16));
 sky130_fd_sc_hd__buf_2 output72 (.A(net931),
    .X(out17));
 sky130_fd_sc_hd__buf_2 output73 (.A(net932),
    .X(out18));
 sky130_fd_sc_hd__buf_2 output74 (.A(net933),
    .X(out19));
 sky130_fd_sc_hd__clkbuf_1 output75 (.A(clknet_1_0__leaf_net934),
    .X(out2));
 sky130_fd_sc_hd__clkbuf_1 output76 (.A(net935),
    .X(out20));
 sky130_fd_sc_hd__buf_2 output77 (.A(net936),
    .X(out21));
 sky130_fd_sc_hd__clkbuf_1 output78 (.A(clknet_1_1__leaf_net937),
    .X(out22));
 sky130_fd_sc_hd__clkbuf_1 output79 (.A(clknet_1_1__leaf_net938),
    .X(out23));
 sky130_fd_sc_hd__buf_2 output80 (.A(net1023),
    .X(out24));
 sky130_fd_sc_hd__buf_2 output81 (.A(net940),
    .X(out25));
 sky130_fd_sc_hd__clkbuf_1 output82 (.A(net941),
    .X(out27));
 sky130_fd_sc_hd__clkbuf_4 output83 (.A(net942),
    .X(out28));
 sky130_fd_sc_hd__clkbuf_4 output84 (.A(net943),
    .X(out29));
 sky130_fd_sc_hd__buf_2 output85 (.A(net944),
    .X(out3));
 sky130_fd_sc_hd__clkbuf_1 output86 (.A(clknet_1_1__leaf_net945),
    .X(out30));
 sky130_fd_sc_hd__clkbuf_1 output87 (.A(clknet_1_1__leaf_net946),
    .X(out31));
 sky130_fd_sc_hd__clkbuf_1 output88 (.A(clknet_1_1__leaf_net947),
    .X(out32));
 sky130_fd_sc_hd__buf_2 output89 (.A(net948),
    .X(out34));
 sky130_fd_sc_hd__clkbuf_4 output90 (.A(net949),
    .X(out36));
 sky130_fd_sc_hd__buf_2 output91 (.A(net950),
    .X(out38));
 sky130_fd_sc_hd__buf_2 output92 (.A(net951),
    .X(out39));
 sky130_fd_sc_hd__clkbuf_1 output93 (.A(clknet_1_0__leaf_net952),
    .X(out4));
 sky130_fd_sc_hd__buf_2 output94 (.A(net953),
    .X(out40));
 sky130_fd_sc_hd__clkbuf_1 output95 (.A(clknet_1_1__leaf_net954),
    .X(out41));
 sky130_fd_sc_hd__buf_2 output96 (.A(net955),
    .X(out42));
 sky130_fd_sc_hd__buf_2 output97 (.A(net956),
    .X(out43));
 sky130_fd_sc_hd__clkbuf_1 output98 (.A(clknet_1_1__leaf_net957),
    .X(out44));
 sky130_fd_sc_hd__clkbuf_1 output99 (.A(net958),
    .X(out45));
 sky130_fd_sc_hd__clkbuf_1 output100 (.A(clknet_1_1__leaf_net959),
    .X(out46));
 sky130_fd_sc_hd__buf_2 output101 (.A(net960),
    .X(out47));
 sky130_fd_sc_hd__buf_2 output102 (.A(net961),
    .X(out48));
 sky130_fd_sc_hd__buf_2 output103 (.A(net962),
    .X(out49));
 sky130_fd_sc_hd__buf_2 output104 (.A(net963),
    .X(out5));
 sky130_fd_sc_hd__clkbuf_1 output105 (.A(net964),
    .X(out50));
 sky130_fd_sc_hd__clkbuf_1 output106 (.A(clknet_1_1__leaf_net965),
    .X(out51));
 sky130_fd_sc_hd__clkbuf_4 output107 (.A(net966),
    .X(out52));
 sky130_fd_sc_hd__clkbuf_4 output108 (.A(net967),
    .X(out53));
 sky130_fd_sc_hd__buf_2 output109 (.A(net968),
    .X(out54));
 sky130_fd_sc_hd__clkbuf_4 output110 (.A(net969),
    .X(out55));
 sky130_fd_sc_hd__clkbuf_4 output111 (.A(net970),
    .X(out56));
 sky130_fd_sc_hd__clkbuf_1 output112 (.A(clknet_1_1__leaf_net971),
    .X(out57));
 sky130_fd_sc_hd__clkbuf_1 output113 (.A(clknet_1_1__leaf_net972),
    .X(out58));
 sky130_fd_sc_hd__clkbuf_1 output114 (.A(clknet_1_0__leaf_net973),
    .X(out6));
 sky130_fd_sc_hd__clkbuf_1 output115 (.A(clknet_1_1__leaf_net974),
    .X(out60));
 sky130_fd_sc_hd__buf_2 output116 (.A(net975),
    .X(out61));
 sky130_fd_sc_hd__buf_2 output117 (.A(net976),
    .X(out7));
 sky130_fd_sc_hd__clkbuf_1 output118 (.A(clknet_1_1__leaf_net977),
    .X(out8));
 sky130_fd_sc_hd__buf_2 output119 (.A(net978),
    .X(out9));
 sky130_fd_sc_hd__buf_2 fanout120 (.A(net447),
    .X(net979));
 sky130_fd_sc_hd__clkbuf_4 fanout121 (.A(net209),
    .X(net980));
 sky130_fd_sc_hd__clkbuf_4 fanout122 (.A(net328),
    .X(net981));
 sky130_fd_sc_hd__buf_2 fanout123 (.A(net320),
    .X(net982));
 sky130_fd_sc_hd__clkbuf_4 fanout124 (.A(net985),
    .X(net983));
 sky130_fd_sc_hd__buf_1 fanout125 (.A(net985),
    .X(net984));
 sky130_fd_sc_hd__buf_4 fanout126 (.A(net344),
    .X(net985));
 sky130_fd_sc_hd__clkbuf_4 fanout127 (.A(net318),
    .X(net986));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout128 (.A(net318),
    .X(net987));
 sky130_fd_sc_hd__buf_4 fanout129 (.A(net104),
    .X(net988));
 sky130_fd_sc_hd__clkbuf_4 fanout130 (.A(net204),
    .X(net989));
 sky130_fd_sc_hd__clkbuf_4 fanout131 (.A(net203),
    .X(net990));
 sky130_fd_sc_hd__clkbuf_2 fanout132 (.A(net203),
    .X(net991));
 sky130_fd_sc_hd__buf_2 fanout133 (.A(net993),
    .X(net992));
 sky130_fd_sc_hd__buf_2 fanout134 (.A(net372),
    .X(net993));
 sky130_fd_sc_hd__buf_4 fanout135 (.A(net312),
    .X(net994));
 sky130_fd_sc_hd__buf_4 fanout136 (.A(net310),
    .X(net995));
 sky130_fd_sc_hd__clkbuf_4 fanout137 (.A(net90),
    .X(net996));
 sky130_fd_sc_hd__buf_4 fanout138 (.A(net18),
    .X(net997));
 sky130_fd_sc_hd__clkbuf_4 fanout139 (.A(net17),
    .X(net998));
 sky130_fd_sc_hd__buf_6 fanout140 (.A(net196),
    .X(net999));
 sky130_fd_sc_hd__buf_4 fanout141 (.A(net122),
    .X(net1000));
 sky130_fd_sc_hd__buf_12 fanout142 (.A(net81),
    .X(net1001));
 sky130_fd_sc_hd__buf_8 fanout143 (.A(net77),
    .X(net1002));
 sky130_fd_sc_hd__clkbuf_8 fanout144 (.A(net115),
    .X(net1003));
 sky130_fd_sc_hd__buf_8 fanout145 (.A(net78),
    .X(net1004));
 sky130_fd_sc_hd__buf_4 fanout146 (.A(net97),
    .X(net1005));
 sky130_fd_sc_hd__buf_12 fanout147 (.A(net1007),
    .X(net1006));
 sky130_fd_sc_hd__buf_8 fanout148 (.A(net72),
    .X(net1007));
 sky130_fd_sc_hd__buf_2 fanout149 (.A(net1010),
    .X(net1008));
 sky130_fd_sc_hd__clkbuf_4 fanout150 (.A(net1010),
    .X(net1009));
 sky130_fd_sc_hd__buf_2 fanout151 (.A(net34),
    .X(net1010));
 sky130_fd_sc_hd__buf_2 fanout152 (.A(net1012),
    .X(net1011));
 sky130_fd_sc_hd__buf_2 fanout153 (.A(net1013),
    .X(net1012));
 sky130_fd_sc_hd__clkbuf_2 fanout154 (.A(net528),
    .X(net1013));
 sky130_fd_sc_hd__buf_2 fanout155 (.A(net525),
    .X(net1014));
 sky130_fd_sc_hd__buf_1 fanout156 (.A(net525),
    .X(net1015));
 sky130_fd_sc_hd__buf_2 fanout157 (.A(net422),
    .X(net1016));
 sky130_fd_sc_hd__clkbuf_2 fanout158 (.A(net422),
    .X(net1017));
 sky130_fd_sc_hd__clkbuf_4 fanout159 (.A(net249),
    .X(net1018));
 sky130_fd_sc_hd__clkbuf_4 fanout160 (.A(net70),
    .X(net1019));
 sky130_fd_sc_hd__buf_12 fanout161 (.A(net70),
    .X(net1020));
 sky130_fd_sc_hd__clkbuf_4 fanout162 (.A(net841),
    .X(net1021));
 sky130_fd_sc_hd__buf_4 fanout163 (.A(net951),
    .X(net1022));
 sky130_fd_sc_hd__clkbuf_4 fanout164 (.A(net939),
    .X(net1023));
 sky130_fd_sc_hd__buf_4 fanout165 (.A(net788),
    .X(net1024));
 sky130_fd_sc_hd__buf_2 fanout166 (.A(net788),
    .X(net1025));
 sky130_fd_sc_hd__buf_4 fanout167 (.A(net923),
    .X(net1026));
 sky130_fd_sc_hd__buf_4 fanout168 (.A(net963),
    .X(net1027));
 sky130_fd_sc_hd__clkbuf_4 fanout169 (.A(net750),
    .X(net1028));
 sky130_fd_sc_hd__buf_2 max_cap170 (.A(net749),
    .X(net1029));
 sky130_fd_sc_hd__buf_4 fanout171 (.A(net698),
    .X(net1030));
 sky130_fd_sc_hd__buf_2 fanout172 (.A(net698),
    .X(net1031));
 sky130_fd_sc_hd__clkbuf_4 fanout173 (.A(net5),
    .X(net1032));
 sky130_fd_sc_hd__buf_4 max_cap174 (.A(net215),
    .X(net1033));
 sky130_fd_sc_hd__buf_8 fanout175 (.A(net68),
    .X(net1034));
 sky130_fd_sc_hd__clkbuf_8 fanout176 (.A(net865),
    .X(net1035));
 sky130_fd_sc_hd__buf_4 fanout177 (.A(net918),
    .X(net1036));
 sky130_fd_sc_hd__clkbuf_2 fanout178 (.A(net918),
    .X(net1037));
 sky130_fd_sc_hd__buf_4 fanout179 (.A(net903),
    .X(net1038));
 sky130_fd_sc_hd__buf_2 fanout180 (.A(net903),
    .X(net1039));
 sky130_fd_sc_hd__clkbuf_4 fanout181 (.A(net1041),
    .X(net1040));
 sky130_fd_sc_hd__buf_2 fanout182 (.A(net901),
    .X(net1041));
 sky130_fd_sc_hd__buf_4 fanout183 (.A(net894),
    .X(net1042));
 sky130_fd_sc_hd__buf_4 fanout184 (.A(net891),
    .X(net1043));
 sky130_fd_sc_hd__buf_4 fanout185 (.A(net890),
    .X(net1044));
 sky130_fd_sc_hd__clkbuf_8 fanout186 (.A(net885),
    .X(net1045));
 sky130_fd_sc_hd__buf_4 fanout187 (.A(net872),
    .X(net1046));
 sky130_fd_sc_hd__clkbuf_4 fanout188 (.A(net1048),
    .X(net1047));
 sky130_fd_sc_hd__clkbuf_4 fanout189 (.A(net133),
    .X(net1048));
 sky130_fd_sc_hd__buf_8 fanout190 (.A(net1050),
    .X(net1049));
 sky130_fd_sc_hd__buf_12 fanout191 (.A(net1051),
    .X(net1050));
 sky130_fd_sc_hd__buf_12 fanout192 (.A(net133),
    .X(net1051));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net854 (.A(net854),
    .X(clknet_0_net854));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net854 (.A(clknet_0_net854),
    .X(clknet_1_0__leaf_net854));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net854 (.A(clknet_0_net854),
    .X(clknet_1_1__leaf_net854));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net706 (.A(net706),
    .X(clknet_0_net706));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net706 (.A(clknet_0_net706),
    .X(clknet_1_0__leaf_net706));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net706 (.A(clknet_0_net706),
    .X(clknet_1_1__leaf_net706));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net623 (.A(net623),
    .X(clknet_0_net623));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net623 (.A(clknet_0_net623),
    .X(clknet_1_0__leaf_net623));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net623 (.A(clknet_0_net623),
    .X(clknet_1_1__leaf_net623));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net585 (.A(net585),
    .X(clknet_0_net585));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net585 (.A(clknet_0_net585),
    .X(clknet_1_0__leaf_net585));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net585 (.A(clknet_0_net585),
    .X(clknet_1_1__leaf_net585));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net425 (.A(net425),
    .X(clknet_0_net425));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net425 (.A(clknet_0_net425),
    .X(clknet_1_0__leaf_net425));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net425 (.A(clknet_0_net425),
    .X(clknet_1_1__leaf_net425));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net433 (.A(net433),
    .X(clknet_0_net433));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net433 (.A(clknet_0_net433),
    .X(clknet_1_0__leaf_net433));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net433 (.A(clknet_0_net433),
    .X(clknet_1_1__leaf_net433));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net423 (.A(net423),
    .X(clknet_0_net423));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net423 (.A(clknet_0_net423),
    .X(clknet_1_0__leaf_net423));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net423 (.A(clknet_0_net423),
    .X(clknet_1_1__leaf_net423));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net934 (.A(net934),
    .X(clknet_0_net934));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net934 (.A(clknet_0_net934),
    .X(clknet_1_0__leaf_net934));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net934 (.A(clknet_0_net934),
    .X(clknet_1_1__leaf_net934));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net517 (.A(net517),
    .X(clknet_0_net517));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net517 (.A(clknet_0_net517),
    .X(clknet_1_0__leaf_net517));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net517 (.A(clknet_0_net517),
    .X(clknet_1_1__leaf_net517));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net490 (.A(net490),
    .X(clknet_0_net490));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net490 (.A(clknet_0_net490),
    .X(clknet_1_0__leaf_net490));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net490 (.A(clknet_0_net490),
    .X(clknet_1_1__leaf_net490));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net493 (.A(net493),
    .X(clknet_0_net493));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net493 (.A(clknet_0_net493),
    .X(clknet_1_0__leaf_net493));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net493 (.A(clknet_0_net493),
    .X(clknet_1_1__leaf_net493));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net835 (.A(net835),
    .X(clknet_0_net835));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net835 (.A(clknet_0_net835),
    .X(clknet_1_0__leaf_net835));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net835 (.A(clknet_0_net835),
    .X(clknet_1_1__leaf_net835));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net499 (.A(net499),
    .X(clknet_0_net499));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net499 (.A(clknet_0_net499),
    .X(clknet_1_0__leaf_net499));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net499 (.A(clknet_0_net499),
    .X(clknet_1_1__leaf_net499));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net498 (.A(net498),
    .X(clknet_0_net498));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net498 (.A(clknet_0_net498),
    .X(clknet_1_0__leaf_net498));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net498 (.A(clknet_0_net498),
    .X(clknet_1_1__leaf_net498));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net833 (.A(net833),
    .X(clknet_0_net833));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net833 (.A(clknet_0_net833),
    .X(clknet_1_0__leaf_net833));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net833 (.A(clknet_0_net833),
    .X(clknet_1_1__leaf_net833));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net973 (.A(net973),
    .X(clknet_0_net973));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net973 (.A(clknet_0_net973),
    .X(clknet_1_0__leaf_net973));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net973 (.A(clknet_0_net973),
    .X(clknet_1_1__leaf_net973));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net922 (.A(net922),
    .X(clknet_0_net922));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net922 (.A(clknet_0_net922),
    .X(clknet_1_0__leaf_net922));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net922 (.A(clknet_0_net922),
    .X(clknet_1_1__leaf_net922));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net522 (.A(net522),
    .X(clknet_0_net522));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net522 (.A(clknet_0_net522),
    .X(clknet_1_0__leaf_net522));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net522 (.A(clknet_0_net522),
    .X(clknet_1_1__leaf_net522));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net617 (.A(net617),
    .X(clknet_0_net617));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net617 (.A(clknet_0_net617),
    .X(clknet_1_0__leaf_net617));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net617 (.A(clknet_0_net617),
    .X(clknet_1_1__leaf_net617));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net834 (.A(net834),
    .X(clknet_0_net834));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net834 (.A(clknet_0_net834),
    .X(clknet_1_0__leaf_net834));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net834 (.A(clknet_0_net834),
    .X(clknet_1_1__leaf_net834));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net508 (.A(net508),
    .X(clknet_0_net508));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net508 (.A(clknet_0_net508),
    .X(clknet_1_0__leaf_net508));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net508 (.A(clknet_0_net508),
    .X(clknet_1_1__leaf_net508));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net510 (.A(net510),
    .X(clknet_0_net510));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net510 (.A(clknet_0_net510),
    .X(clknet_1_0__leaf_net510));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net510 (.A(clknet_0_net510),
    .X(clknet_1_1__leaf_net510));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net515 (.A(net515),
    .X(clknet_0_net515));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net515 (.A(clknet_0_net515),
    .X(clknet_1_0__leaf_net515));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net515 (.A(clknet_0_net515),
    .X(clknet_1_1__leaf_net515));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net483 (.A(net483),
    .X(clknet_0_net483));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net483 (.A(clknet_0_net483),
    .X(clknet_1_0__leaf_net483));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net483 (.A(clknet_0_net483),
    .X(clknet_1_1__leaf_net483));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net606 (.A(net606),
    .X(clknet_0_net606));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net606 (.A(clknet_0_net606),
    .X(clknet_1_0__leaf_net606));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net606 (.A(clknet_0_net606),
    .X(clknet_1_1__leaf_net606));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net465 (.A(net465),
    .X(clknet_0_net465));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net465 (.A(clknet_0_net465),
    .X(clknet_1_0__leaf_net465));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net465 (.A(clknet_0_net465),
    .X(clknet_1_1__leaf_net465));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net471 (.A(net471),
    .X(clknet_0_net471));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net471 (.A(clknet_0_net471),
    .X(clknet_1_0__leaf_net471));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net471 (.A(clknet_0_net471),
    .X(clknet_1_1__leaf_net471));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net461 (.A(net461),
    .X(clknet_0_net461));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net461 (.A(clknet_0_net461),
    .X(clknet_1_0__leaf_net461));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net461 (.A(clknet_0_net461),
    .X(clknet_1_1__leaf_net461));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net474 (.A(net474),
    .X(clknet_0_net474));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net474 (.A(clknet_0_net474),
    .X(clknet_1_0__leaf_net474));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net474 (.A(clknet_0_net474),
    .X(clknet_1_1__leaf_net474));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net853 (.A(net853),
    .X(clknet_0_net853));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net853 (.A(clknet_0_net853),
    .X(clknet_1_0__leaf_net853));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net853 (.A(clknet_0_net853),
    .X(clknet_1_1__leaf_net853));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net604 (.A(net604),
    .X(clknet_0_net604));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net604 (.A(clknet_0_net604),
    .X(clknet_1_0__leaf_net604));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net604 (.A(clknet_0_net604),
    .X(clknet_1_1__leaf_net604));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net591 (.A(net591),
    .X(clknet_0_net591));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net591 (.A(clknet_0_net591),
    .X(clknet_1_0__leaf_net591));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net591 (.A(clknet_0_net591),
    .X(clknet_1_1__leaf_net591));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net469 (.A(net469),
    .X(clknet_0_net469));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net469 (.A(clknet_0_net469),
    .X(clknet_1_0__leaf_net469));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net469 (.A(clknet_0_net469),
    .X(clknet_1_1__leaf_net469));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net852 (.A(net852),
    .X(clknet_0_net852));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net852 (.A(clknet_0_net852),
    .X(clknet_1_0__leaf_net852));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net852 (.A(clknet_0_net852),
    .X(clknet_1_1__leaf_net852));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net595 (.A(net595),
    .X(clknet_0_net595));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net595 (.A(clknet_0_net595),
    .X(clknet_1_0__leaf_net595));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net595 (.A(clknet_0_net595),
    .X(clknet_1_1__leaf_net595));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net924 (.A(net924),
    .X(clknet_0_net924));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net924 (.A(clknet_0_net924),
    .X(clknet_1_0__leaf_net924));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net924 (.A(clknet_0_net924),
    .X(clknet_1_1__leaf_net924));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net815 (.A(net815),
    .X(clknet_0_net815));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net815 (.A(clknet_0_net815),
    .X(clknet_1_0__leaf_net815));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net815 (.A(clknet_0_net815),
    .X(clknet_1_1__leaf_net815));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net927 (.A(net927),
    .X(clknet_0_net927));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net927 (.A(clknet_0_net927),
    .X(clknet_1_0__leaf_net927));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net927 (.A(clknet_0_net927),
    .X(clknet_1_1__leaf_net927));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net506 (.A(net506),
    .X(clknet_0_net506));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net506 (.A(clknet_0_net506),
    .X(clknet_1_0__leaf_net506));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net506 (.A(clknet_0_net506),
    .X(clknet_1_1__leaf_net506));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net954 (.A(net954),
    .X(clknet_0_net954));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net954 (.A(clknet_0_net954),
    .X(clknet_1_0__leaf_net954));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net954 (.A(clknet_0_net954),
    .X(clknet_1_1__leaf_net954));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net938 (.A(net938),
    .X(clknet_0_net938));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net938 (.A(clknet_0_net938),
    .X(clknet_1_0__leaf_net938));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net938 (.A(clknet_0_net938),
    .X(clknet_1_1__leaf_net938));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net977 (.A(net977),
    .X(clknet_0_net977));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net977 (.A(clknet_0_net977),
    .X(clknet_1_0__leaf_net977));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net977 (.A(clknet_0_net977),
    .X(clknet_1_1__leaf_net977));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net799 (.A(net799),
    .X(clknet_0_net799));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net799 (.A(clknet_0_net799),
    .X(clknet_1_0__leaf_net799));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net799 (.A(clknet_0_net799),
    .X(clknet_1_1__leaf_net799));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net330 (.A(net330),
    .X(clknet_0_net330));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net330 (.A(clknet_0_net330),
    .X(clknet_1_0__leaf_net330));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net330 (.A(clknet_0_net330),
    .X(clknet_1_1__leaf_net330));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net798 (.A(net798),
    .X(clknet_0_net798));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net798 (.A(clknet_0_net798),
    .X(clknet_1_0__leaf_net798));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net798 (.A(clknet_0_net798),
    .X(clknet_1_1__leaf_net798));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net303 (.A(net303),
    .X(clknet_0_net303));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net303 (.A(clknet_0_net303),
    .X(clknet_1_0__leaf_net303));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net303 (.A(clknet_0_net303),
    .X(clknet_1_1__leaf_net303));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net705 (.A(net705),
    .X(clknet_0_net705));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net705 (.A(clknet_0_net705),
    .X(clknet_1_0__leaf_net705));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net705 (.A(clknet_0_net705),
    .X(clknet_1_1__leaf_net705));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net302 (.A(net302),
    .X(clknet_0_net302));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net302 (.A(clknet_0_net302),
    .X(clknet_1_0__leaf_net302));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net302 (.A(clknet_0_net302),
    .X(clknet_1_1__leaf_net302));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net946 (.A(net946),
    .X(clknet_0_net946));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net946 (.A(clknet_0_net946),
    .X(clknet_1_0__leaf_net946));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net946 (.A(clknet_0_net946),
    .X(clknet_1_1__leaf_net946));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net397 (.A(net397),
    .X(clknet_0_net397));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net397 (.A(clknet_0_net397),
    .X(clknet_1_0__leaf_net397));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net397 (.A(clknet_0_net397),
    .X(clknet_1_1__leaf_net397));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net386 (.A(net386),
    .X(clknet_0_net386));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net386 (.A(clknet_0_net386),
    .X(clknet_1_0__leaf_net386));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net386 (.A(clknet_0_net386),
    .X(clknet_1_1__leaf_net386));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net952 (.A(net952),
    .X(clknet_0_net952));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net952 (.A(clknet_0_net952),
    .X(clknet_1_0__leaf_net952));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net952 (.A(clknet_0_net952),
    .X(clknet_1_1__leaf_net952));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net282 (.A(net282),
    .X(clknet_0_net282));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net282 (.A(clknet_0_net282),
    .X(clknet_1_0__leaf_net282));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net282 (.A(clknet_0_net282),
    .X(clknet_1_1__leaf_net282));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net761 (.A(net761),
    .X(clknet_0_net761));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net761 (.A(clknet_0_net761),
    .X(clknet_1_0__leaf_net761));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net761 (.A(clknet_0_net761),
    .X(clknet_1_1__leaf_net761));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net191 (.A(net191),
    .X(clknet_0_net191));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net191 (.A(clknet_0_net191),
    .X(clknet_1_0__leaf_net191));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net191 (.A(clknet_0_net191),
    .X(clknet_1_1__leaf_net191));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net743 (.A(net743),
    .X(clknet_0_net743));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net743 (.A(clknet_0_net743),
    .X(clknet_1_0__leaf_net743));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net743 (.A(clknet_0_net743),
    .X(clknet_1_1__leaf_net743));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net49 (.A(net49),
    .X(clknet_0_net49));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net49 (.A(clknet_0_net49),
    .X(clknet_1_0__leaf_net49));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net49 (.A(clknet_0_net49),
    .X(clknet_1_1__leaf_net49));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net971 (.A(net971),
    .X(clknet_0_net971));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net971 (.A(clknet_0_net971),
    .X(clknet_1_0__leaf_net971));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net971 (.A(clknet_0_net971),
    .X(clknet_1_1__leaf_net971));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net52 (.A(net52),
    .X(clknet_0_net52));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net52 (.A(clknet_0_net52),
    .X(clknet_1_0__leaf_net52));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net52 (.A(clknet_0_net52),
    .X(clknet_1_1__leaf_net52));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net57 (.A(net57),
    .X(clknet_0_net57));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net57 (.A(clknet_0_net57),
    .X(clknet_1_0__leaf_net57));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net57 (.A(clknet_0_net57),
    .X(clknet_1_1__leaf_net57));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net744 (.A(net744),
    .X(clknet_0_net744));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net744 (.A(clknet_0_net744),
    .X(clknet_1_0__leaf_net744));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net744 (.A(clknet_0_net744),
    .X(clknet_1_1__leaf_net744));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net179 (.A(net179),
    .X(clknet_0_net179));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net179 (.A(clknet_0_net179),
    .X(clknet_1_0__leaf_net179));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net179 (.A(clknet_0_net179),
    .X(clknet_1_1__leaf_net179));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net181 (.A(net181),
    .X(clknet_0_net181));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net181 (.A(clknet_0_net181),
    .X(clknet_1_0__leaf_net181));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net181 (.A(clknet_0_net181),
    .X(clknet_1_1__leaf_net181));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net937 (.A(net937),
    .X(clknet_0_net937));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net937 (.A(clknet_0_net937),
    .X(clknet_1_0__leaf_net937));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net937 (.A(clknet_0_net937),
    .X(clknet_1_1__leaf_net937));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net972 (.A(net972),
    .X(clknet_0_net972));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net972 (.A(clknet_0_net972),
    .X(clknet_1_0__leaf_net972));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net972 (.A(clknet_0_net972),
    .X(clknet_1_1__leaf_net972));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net153 (.A(net153),
    .X(clknet_0_net153));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net153 (.A(clknet_0_net153),
    .X(clknet_1_0__leaf_net153));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net153 (.A(clknet_0_net153),
    .X(clknet_1_1__leaf_net153));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net797 (.A(net797),
    .X(clknet_0_net797));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net797 (.A(clknet_0_net797),
    .X(clknet_1_0__leaf_net797));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net797 (.A(clknet_0_net797),
    .X(clknet_1_1__leaf_net797));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net947 (.A(net947),
    .X(clknet_0_net947));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net947 (.A(clknet_0_net947),
    .X(clknet_1_0__leaf_net947));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net947 (.A(net1060),
    .X(clknet_1_1__leaf_net947));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net401 (.A(net401),
    .X(clknet_0_net401));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net401 (.A(clknet_0_net401),
    .X(clknet_1_0__leaf_net401));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net401 (.A(clknet_0_net401),
    .X(clknet_1_1__leaf_net401));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net945 (.A(net945),
    .X(clknet_0_net945));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net945 (.A(clknet_0_net945),
    .X(clknet_1_0__leaf_net945));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net945 (.A(clknet_0_net945),
    .X(clknet_1_1__leaf_net945));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net403 (.A(net403),
    .X(clknet_0_net403));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net403 (.A(clknet_0_net403),
    .X(clknet_1_0__leaf_net403));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net403 (.A(clknet_0_net403),
    .X(clknet_1_1__leaf_net403));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net300 (.A(net300),
    .X(clknet_0_net300));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net300 (.A(clknet_0_net300),
    .X(clknet_1_0__leaf_net300));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net300 (.A(clknet_0_net300),
    .X(clknet_1_1__leaf_net300));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net145 (.A(net145),
    .X(clknet_0_net145));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net145 (.A(clknet_0_net145),
    .X(clknet_1_0__leaf_net145));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net145 (.A(clknet_0_net145),
    .X(clknet_1_1__leaf_net145));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net62 (.A(net62),
    .X(clknet_0_net62));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net62 (.A(clknet_0_net62),
    .X(clknet_1_0__leaf_net62));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net62 (.A(clknet_0_net62),
    .X(clknet_1_1__leaf_net62));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net182 (.A(net182),
    .X(clknet_0_net182));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net182 (.A(clknet_0_net182),
    .X(clknet_1_0__leaf_net182));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net182 (.A(clknet_0_net182),
    .X(clknet_1_1__leaf_net182));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net188 (.A(net188),
    .X(clknet_0_net188));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net188 (.A(clknet_0_net188),
    .X(clknet_1_0__leaf_net188));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net188 (.A(clknet_0_net188),
    .X(clknet_1_1__leaf_net188));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net185 (.A(net185),
    .X(clknet_0_net185));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net185 (.A(clknet_0_net185),
    .X(clknet_1_0__leaf_net185));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net185 (.A(clknet_0_net185),
    .X(clknet_1_1__leaf_net185));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net184 (.A(net184),
    .X(clknet_0_net184));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net184 (.A(clknet_0_net184),
    .X(clknet_1_0__leaf_net184));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net184 (.A(clknet_0_net184),
    .X(clknet_1_1__leaf_net184));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net67 (.A(net67),
    .X(clknet_0_net67));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net67 (.A(clknet_0_net67),
    .X(clknet_1_0__leaf_net67));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net67 (.A(clknet_0_net67),
    .X(clknet_1_1__leaf_net67));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net959 (.A(net959),
    .X(clknet_0_net959));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net959 (.A(clknet_0_net959),
    .X(clknet_1_0__leaf_net959));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net959 (.A(clknet_0_net959),
    .X(clknet_1_1__leaf_net959));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net974 (.A(net974),
    .X(clknet_0_net974));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net974 (.A(clknet_0_net974),
    .X(clknet_1_0__leaf_net974));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net974 (.A(clknet_0_net974),
    .X(clknet_1_1__leaf_net974));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net177 (.A(net177),
    .X(clknet_0_net177));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net177 (.A(clknet_0_net177),
    .X(clknet_1_0__leaf_net177));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net177 (.A(clknet_0_net177),
    .X(clknet_1_1__leaf_net177));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net60 (.A(net60),
    .X(clknet_0_net60));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net60 (.A(clknet_0_net60),
    .X(clknet_1_0__leaf_net60));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net60 (.A(clknet_0_net60),
    .X(clknet_1_1__leaf_net60));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net56 (.A(net56),
    .X(clknet_0_net56));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net56 (.A(clknet_0_net56),
    .X(clknet_1_0__leaf_net56));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net56 (.A(clknet_0_net56),
    .X(clknet_1_1__leaf_net56));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net965 (.A(net965),
    .X(clknet_0_net965));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net965 (.A(clknet_0_net965),
    .X(clknet_1_0__leaf_net965));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net965 (.A(clknet_0_net965),
    .X(clknet_1_1__leaf_net965));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net54 (.A(net54),
    .X(clknet_0_net54));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net54 (.A(clknet_0_net54),
    .X(clknet_1_0__leaf_net54));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net54 (.A(clknet_0_net54),
    .X(clknet_1_1__leaf_net54));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net48 (.A(net48),
    .X(clknet_0_net48));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net48 (.A(clknet_0_net48),
    .X(clknet_1_0__leaf_net48));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net48 (.A(clknet_0_net48),
    .X(clknet_1_1__leaf_net48));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net50 (.A(net50),
    .X(clknet_0_net50));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net50 (.A(clknet_0_net50),
    .X(clknet_1_0__leaf_net50));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net50 (.A(clknet_0_net50),
    .X(clknet_1_1__leaf_net50));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net171 (.A(net171),
    .X(clknet_0_net171));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net171 (.A(clknet_0_net171),
    .X(clknet_1_0__leaf_net171));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net171 (.A(clknet_0_net171),
    .X(clknet_1_1__leaf_net171));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net957 (.A(net957),
    .X(clknet_0_net957));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net957 (.A(clknet_0_net957),
    .X(clknet_1_0__leaf_net957));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net957 (.A(clknet_0_net957),
    .X(clknet_1_1__leaf_net957));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net762 (.A(net762),
    .X(clknet_0_net762));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net762 (.A(clknet_0_net762),
    .X(clknet_1_0__leaf_net762));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net762 (.A(clknet_0_net762),
    .X(clknet_1_1__leaf_net762));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net780 (.A(net780),
    .X(clknet_0_net780));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net780 (.A(clknet_0_net780),
    .X(clknet_1_0__leaf_net780));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net780 (.A(clknet_0_net780),
    .X(clknet_1_1__leaf_net780));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net273 (.A(net273),
    .X(clknet_0_net273));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net273 (.A(clknet_0_net273),
    .X(clknet_1_0__leaf_net273));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net273 (.A(clknet_0_net273),
    .X(clknet_1_1__leaf_net273));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net275 (.A(net275),
    .X(clknet_0_net275));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net275 (.A(clknet_0_net275),
    .X(clknet_1_0__leaf_net275));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net275 (.A(clknet_0_net275),
    .X(clknet_1_1__leaf_net275));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net251 (.A(net251),
    .X(clknet_0_net251));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net251 (.A(clknet_0_net251),
    .X(clknet_1_0__leaf_net251));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net251 (.A(clknet_0_net251),
    .X(clknet_1_1__leaf_net251));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net257 (.A(net257),
    .X(clknet_0_net257));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net257 (.A(clknet_0_net257),
    .X(clknet_1_0__leaf_net257));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net257 (.A(clknet_0_net257),
    .X(clknet_1_1__leaf_net257));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net253 (.A(net253),
    .X(clknet_0_net253));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net253 (.A(clknet_0_net253),
    .X(clknet_1_0__leaf_net253));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net253 (.A(clknet_0_net253),
    .X(clknet_1_1__leaf_net253));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net246 (.A(net246),
    .X(clknet_0_net246));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net246 (.A(clknet_0_net246),
    .X(clknet_1_0__leaf_net246));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net246 (.A(clknet_0_net246),
    .X(clknet_1_1__leaf_net246));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net475 (.A(net475),
    .X(clknet_0_net475));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net475 (.A(clknet_0_net475),
    .X(clknet_1_0__leaf_net475));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net475 (.A(clknet_0_net475),
    .X(clknet_1_1__leaf_net475));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net462 (.A(net462),
    .X(clknet_0_net462));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net462 (.A(clknet_0_net462),
    .X(clknet_1_0__leaf_net462));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net462 (.A(clknet_0_net462),
    .X(clknet_1_1__leaf_net462));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net369 (.A(net369),
    .X(clknet_0_net369));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net369 (.A(clknet_0_net369),
    .X(clknet_1_0__leaf_net369));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net369 (.A(clknet_0_net369),
    .X(clknet_1_1__leaf_net369));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net245 (.A(net245),
    .X(clknet_0_net245));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net245 (.A(clknet_0_net245),
    .X(clknet_1_0__leaf_net245));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net245 (.A(clknet_0_net245),
    .X(clknet_1_1__leaf_net245));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net396 (.A(net396),
    .X(clknet_0_net396));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net396 (.A(clknet_0_net396),
    .X(clknet_1_0__leaf_net396));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net396 (.A(clknet_0_net396),
    .X(clknet_1_1__leaf_net396));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net779 (.A(net779),
    .X(clknet_0_net779));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net779 (.A(clknet_0_net779),
    .X(clknet_1_0__leaf_net779));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net779 (.A(clknet_0_net779),
    .X(clknet_1_1__leaf_net779));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net250 (.A(net250),
    .X(clknet_0_net250));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net250 (.A(clknet_0_net250),
    .X(clknet_1_0__leaf_net250));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net250 (.A(clknet_0_net250),
    .X(clknet_1_1__leaf_net250));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net778 (.A(net778),
    .X(clknet_0_net778));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net778 (.A(clknet_0_net778),
    .X(clknet_1_0__leaf_net778));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net778 (.A(clknet_0_net778),
    .X(clknet_1_1__leaf_net778));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net238 (.A(net238),
    .X(clknet_0_net238));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net238 (.A(clknet_0_net238),
    .X(clknet_1_0__leaf_net238));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net238 (.A(clknet_0_net238),
    .X(clknet_1_1__leaf_net238));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net332 (.A(net332),
    .X(clknet_0_net332));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net332 (.A(clknet_0_net332),
    .X(clknet_1_0__leaf_net332));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net332 (.A(clknet_0_net332),
    .X(clknet_1_1__leaf_net332));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net331 (.A(net331),
    .X(clknet_0_net331));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net331 (.A(clknet_0_net331),
    .X(clknet_1_0__leaf_net331));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net331 (.A(clknet_0_net331),
    .X(clknet_1_1__leaf_net331));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net760 (.A(net760),
    .X(clknet_0_net760));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net760 (.A(clknet_0_net760),
    .X(clknet_1_0__leaf_net760));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net760 (.A(clknet_0_net760),
    .X(clknet_1_1__leaf_net760));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net742 (.A(net742),
    .X(clknet_0_net742));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net742 (.A(clknet_0_net742),
    .X(clknet_1_0__leaf_net742));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net742 (.A(clknet_0_net742),
    .X(clknet_1_1__leaf_net742));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net562 (.A(net562),
    .X(clknet_0_net562));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net562 (.A(clknet_0_net562),
    .X(clknet_1_0__leaf_net562));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net562 (.A(clknet_0_net562),
    .X(clknet_1_1__leaf_net562));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net560 (.A(net560),
    .X(clknet_0_net560));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net560 (.A(clknet_0_net560),
    .X(clknet_1_0__leaf_net560));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net560 (.A(clknet_0_net560),
    .X(clknet_1_1__leaf_net560));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net568 (.A(net568),
    .X(clknet_0_net568));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net568 (.A(clknet_0_net568),
    .X(clknet_1_0__leaf_net568));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net568 (.A(clknet_0_net568),
    .X(clknet_1_1__leaf_net568));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net542 (.A(net542),
    .X(clknet_0_net542));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net542 (.A(clknet_0_net542),
    .X(clknet_1_0__leaf_net542));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net542 (.A(clknet_0_net542),
    .X(clknet_1_1__leaf_net542));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net592 (.A(net592),
    .X(clknet_0_net592));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net592 (.A(clknet_0_net592),
    .X(clknet_1_0__leaf_net592));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net592 (.A(clknet_0_net592),
    .X(clknet_1_1__leaf_net592));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net552 (.A(net552),
    .X(clknet_0_net552));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net552 (.A(clknet_0_net552),
    .X(clknet_1_0__leaf_net552));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net552 (.A(clknet_0_net552),
    .X(clknet_1_1__leaf_net552));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer1 (.A(net77),
    .X(net1052));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer2 (.A(net1052),
    .X(net1053));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer3 (.A(net1052),
    .X(net1054));
 sky130_fd_sc_hd__clkbuf_1 clone4 (.A(net133),
    .X(net1055));
 sky130_fd_sc_hd__dlygate4sd3_1 rebuffer5 (.A(net68),
    .X(net1056));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer6 (.A(net78),
    .X(net1057));
 sky130_fd_sc_hd__clkbuf_1 clone7 (.A(net1050),
    .X(net1058));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer8 (.A(net70),
    .X(net1059));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer9 (.A(clknet_0_net947),
    .X(net1060));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer10 (.A(net1050),
    .X(net1061));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer11 (.A(net1065),
    .X(net1062));
 sky130_fd_sc_hd__clkbuf_1 clone12 (.A(net78),
    .X(net1063));
 sky130_fd_sc_hd__clkbuf_1 clone13 (.A(net68),
    .X(net1064));
 sky130_fd_sc_hd__clkbuf_1 clone14 (.A(net72),
    .X(net1065));
 sky130_fd_sc_hd__clkbuf_1 clone15 (.A(net70),
    .X(net1066));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer16 (.A(net1102),
    .X(net1067));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer17 (.A(net1067),
    .X(net1068));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer18 (.A(net1001),
    .X(net1069));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer19 (.A(net1001),
    .X(net1070));
 sky130_fd_sc_hd__clkbuf_1 clone20 (.A(net1007),
    .X(net1071));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(net851),
    .X(net1072));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(net785),
    .X(net1073));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(net648),
    .X(net1074));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(net805),
    .X(net1075));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(net790),
    .X(net1076));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(net843),
    .X(net1077));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(net786),
    .X(net1078));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(net308),
    .X(net1079));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(net451),
    .X(net1080));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(net757),
    .X(net1081));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(net806),
    .X(net1082));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(net801),
    .X(net1083));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(net334),
    .X(net1084));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(net969),
    .X(net1085));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(net765),
    .X(net1086));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(net849),
    .X(net1087));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(net746),
    .X(net1088));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_A (.DIODE(clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(in0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(in1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(in10));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(in11));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(in12));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(in13));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(in14));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(in15));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(in16));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(in17));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(in18));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(in19));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(in2));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(in20));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(in21));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(in22));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(in23));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(in24));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(in25));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(in26));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(in27));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_A (.DIODE(in28));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_A (.DIODE(in29));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_A (.DIODE(in3));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_A (.DIODE(in30));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_A (.DIODE(in31));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_A (.DIODE(in32));
 sky130_fd_sc_hd__diode_2 ANTENNA_input28_A (.DIODE(in33));
 sky130_fd_sc_hd__diode_2 ANTENNA_input29_A (.DIODE(in34));
 sky130_fd_sc_hd__diode_2 ANTENNA_input30_A (.DIODE(in35));
 sky130_fd_sc_hd__diode_2 ANTENNA_input31_A (.DIODE(in36));
 sky130_fd_sc_hd__diode_2 ANTENNA_input32_A (.DIODE(in37));
 sky130_fd_sc_hd__diode_2 ANTENNA_input33_A (.DIODE(in38));
 sky130_fd_sc_hd__diode_2 ANTENNA_input34_A (.DIODE(in39));
 sky130_fd_sc_hd__diode_2 ANTENNA_input35_A (.DIODE(in4));
 sky130_fd_sc_hd__diode_2 ANTENNA_input36_A (.DIODE(in40));
 sky130_fd_sc_hd__diode_2 ANTENNA_input37_A (.DIODE(in41));
 sky130_fd_sc_hd__diode_2 ANTENNA_input38_A (.DIODE(in42));
 sky130_fd_sc_hd__diode_2 ANTENNA_input39_A (.DIODE(in43));
 sky130_fd_sc_hd__diode_2 ANTENNA_input40_A (.DIODE(in44));
 sky130_fd_sc_hd__diode_2 ANTENNA_input41_A (.DIODE(in45));
 sky130_fd_sc_hd__diode_2 ANTENNA_input42_A (.DIODE(in46));
 sky130_fd_sc_hd__diode_2 ANTENNA_input43_A (.DIODE(in47));
 sky130_fd_sc_hd__diode_2 ANTENNA_input44_A (.DIODE(in48));
 sky130_fd_sc_hd__diode_2 ANTENNA_input45_A (.DIODE(in49));
 sky130_fd_sc_hd__diode_2 ANTENNA_input46_A (.DIODE(in5));
 sky130_fd_sc_hd__diode_2 ANTENNA_input47_A (.DIODE(in50));
 sky130_fd_sc_hd__diode_2 ANTENNA_input48_A (.DIODE(in51));
 sky130_fd_sc_hd__diode_2 ANTENNA_input49_A (.DIODE(in52));
 sky130_fd_sc_hd__diode_2 ANTENNA_input50_A (.DIODE(in53));
 sky130_fd_sc_hd__diode_2 ANTENNA_input51_A (.DIODE(in54));
 sky130_fd_sc_hd__diode_2 ANTENNA_input52_A (.DIODE(in55));
 sky130_fd_sc_hd__diode_2 ANTENNA_input53_A (.DIODE(in56));
 sky130_fd_sc_hd__diode_2 ANTENNA_input54_A (.DIODE(in57));
 sky130_fd_sc_hd__diode_2 ANTENNA_input55_A (.DIODE(in58));
 sky130_fd_sc_hd__diode_2 ANTENNA_input56_A (.DIODE(in59));
 sky130_fd_sc_hd__diode_2 ANTENNA_input57_A (.DIODE(in6));
 sky130_fd_sc_hd__diode_2 ANTENNA_input58_A (.DIODE(in60));
 sky130_fd_sc_hd__diode_2 ANTENNA_input59_A (.DIODE(in61));
 sky130_fd_sc_hd__diode_2 ANTENNA_input60_A (.DIODE(in7));
 sky130_fd_sc_hd__diode_2 ANTENNA_input61_A (.DIODE(in8));
 sky130_fd_sc_hd__diode_2 ANTENNA_input62_A (.DIODE(in9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c63_A0 (.DIODE(net0));
 sky130_fd_sc_hd__diode_2 ANTENNA_c62_X (.DIODE(net0));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_A0 (.DIODE(net0));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_A2 (.DIODE(net0));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_A1 (.DIODE(net0));
 sky130_fd_sc_hd__diode_2 ANTENNA_c198_A3 (.DIODE(net0));
 sky130_fd_sc_hd__diode_2 ANTENNA_c63_X (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_A2 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_A1 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout129_A (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_A0 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_X (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c228_A0 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c222_A3 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_A3 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c206_A4 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_A3 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_A3 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_A0 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_S1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_A3 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_A2 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_X (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c232_A3 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c221_S0 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c220_A0 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_A2 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_A4 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_A2 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_A1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c183_A3 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_X (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_A0 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_S0 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_A1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c611_A0 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_A2 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_A2 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_S0 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c191_A2 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_A1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_A3 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_X (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout144_A (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c183_A1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_A0 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_X (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_A0 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_A2 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c346_A1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_A1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_A1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_S0 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_A3 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_A2 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_S1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c184_A0 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c183_X (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c80_A1 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_c78_S0 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_c74_X (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_A2 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_A0 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_A3 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_c350_A1 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_A0 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_c212_A2 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_A0 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_SCD (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_A3 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_A1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_S1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_A1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c191_A1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c190_A2 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_X (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_A0 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_A1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_A3 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_A2 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_A0 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_X (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_A1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_A1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_A1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_c212_A1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_c203_B1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_SCE (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_c198_A4 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_A0 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_c194_X (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_c235_A1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_c229_A0 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_c221_A3 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_c220_A2 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_A2 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_c212_A3 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_A0 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_SET_B (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_A0 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_c205_A2 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_c203_X (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_c234_A0 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_A0 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_A0 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_c221_A2 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_Q (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_A1 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_A3 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_A1 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_A0 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_A2 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_A2 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA_c215_A4 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_A1 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_X (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout139_A (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_c126_B1 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_c123_B1_N (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_c395_A1 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_c79_X (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge855_D (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA_c244_X (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout138_A (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_c86_A0 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_A1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_c91_B1_N (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_c80_X (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_c86_S1 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c81_X (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c610_A2 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_A1 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_A2 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_A1 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_A0 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_A0 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_A1 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout132_A (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout131_A (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA_c271_X (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout130_A (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_A3 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_A3 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_c272_X (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_c543_S0 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_c528_A1 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_D (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_c279_A3 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_c277_A1 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_c275_X (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge770_A2 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA_c539_A1 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_A3 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_A4 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA_c278_A0 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA_c276_X (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout121_A (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_A2 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_c496_A1 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_c277_X (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_c86_A3 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_c85_A1 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_c84_A1 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_c83_X (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_A2 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_A2 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_A0 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_c208_A2 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_A3 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_A3 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_S0 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_S0 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_S0 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA_c368_A3 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_A3 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_Q_N (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_A0 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_A2 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_A1 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_A1 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_A1 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA_c283_A0 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_Q (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge770_B1 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_A3 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA_c668_A1 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_SCE (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_A3 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA_c405_B1_N (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_A4 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_Q_N (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap174_A (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_c393_A1 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_c323_S1 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_Q (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge767_S1 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA_c674_A1 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA_c546_A0 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA_c540_SCE (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_A2 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_A1 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA_c283_X (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_A2 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_A2 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_A0 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA_c313_A1 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_A2 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_A0 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_A2 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_X (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA_c566_A1 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_c558_A3 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_A0 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_A3 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_A1 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_A2 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_B1_N (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_X (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_c702_A0 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_A4 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA_c687_S0 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA_c565_SET_B (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA_c561_A2 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA_c560_A1 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_A3 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_A1 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_A2 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_A2 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_X (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge773_A0 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_c571_A1 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_A0 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_c297_X (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_A3 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_A1 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c431_A1 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_B1_N (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_A1 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_A3 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_S0 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_A1 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_A1 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_A2 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_X (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_A0 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A0 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_A2 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA_c559_SCD (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA_c555_A1 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_RESET_B (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_A3 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_X (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_A0 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_A2 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c321_A1 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_X (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge853_RESET_B (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA_c346_X (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA_c759_A0 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_A1 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_c742_A1 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_A1 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_A1 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_A2 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_S0 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_A2 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_A4 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_X (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_c70_A2 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_X (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c64_A0 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_A0 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_A1 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_A2 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout136_A (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_A2 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA_c399_X (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_A0 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_A3 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_c430_A1 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_A1 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_c413_A1 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_c412_A3 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_c409_A2 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_c404_X (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_c558_A1 (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA_c547_S0 (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA_c545_A2 (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA_c544_A3 (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA_c532_A4 (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_S0 (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_A1 (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA_c413_A2 (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA_c411_A3 (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA_c410_X (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout122_A (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA_c685_A3 (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_A2 (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_X (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_A0 (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_A1 (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_A0 (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_A1 (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_A2 (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA_c427_D (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA_c424_S1 (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_X (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_A1 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_A1 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_A3 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_c427_Q_N (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_A0 (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_A1 (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA_c434_A2 (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_D (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA_c427_Q (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_A2 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA_c458_A2 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_A1 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_Q_N (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA_c98_Q (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c393_A0 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c248_A0 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c222_A1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_A0 (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_A0 (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_A1 (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_S1 (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA_c577_A2 (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_A0 (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_A3 (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_S0 (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_X (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_A0 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_A1 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_A0 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_A1 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_A2 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_X (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA_c613_A0 (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_S0 (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_A3 (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_A1 (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_S0 (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_A0 (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_A3 (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_A3 (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_X (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA_c237_A1 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_c106_SCE (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_c104_A3 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_c103_A4 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_c102_SCD (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_c101_A1 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_c100_X (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_c745_A0 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_A3 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA_c613_A2 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_A0 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_A1 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_A1 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_X (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA_c66_X (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_c368_A2 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_A0 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_A1 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_c235_A0 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_c221_A1 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_c105_A1 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_A4 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_A0 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_A3 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_c236_A0 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_c112_B1_N (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_c109_S0 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_c105_A3 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_c102_Q_N (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge774_A2 (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge771_A2 (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge767_A0 (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge765_A3 (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA_c676_A0 (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA_c548_A2 (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA_c545_A3 (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA_c540_D (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA_c538_SCE (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA_c529_X (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge771_A3 (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA_c685_A0 (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA_c565_RESET_B (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA_c532_X (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge771_B1 (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge767_S0 (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_A0 (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_A0 (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA_c665_A2 (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA_c547_A2 (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA_c546_A1 (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA_c545_S1 (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA_c536_A1 (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA_c535_X (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_A0 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_A0 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_A1 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_S0 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA_c564_B1 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA_c560_X (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA_c743_A2 (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_A3 (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_A1 (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_A2 (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA_c566_A2 (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA_c565_Q_N (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_A3 (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_A0 (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_A2 (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_A0 (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_A0 (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_A2 (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA_c565_Q (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_A0 (.DIODE(net481));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_A1 (.DIODE(net481));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_A0 (.DIODE(net481));
 sky130_fd_sc_hd__diode_2 ANTENNA_c611_A3 (.DIODE(net481));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_A1 (.DIODE(net481));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_A3 (.DIODE(net481));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_A2 (.DIODE(net481));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_X (.DIODE(net481));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge849_SET_B (.DIODE(net518));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_X (.DIODE(net518));
 sky130_fd_sc_hd__diode_2 ANTENNA_c739_A0 (.DIODE(net541));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A0 (.DIODE(net541));
 sky130_fd_sc_hd__diode_2 ANTENNA_c724_A2 (.DIODE(net541));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_A3 (.DIODE(net541));
 sky130_fd_sc_hd__diode_2 ANTENNA_c677_X (.DIODE(net541));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_A1 (.DIODE(net556));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_S0 (.DIODE(net556));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_A3 (.DIODE(net556));
 sky130_fd_sc_hd__diode_2 ANTENNA_c698_A0 (.DIODE(net556));
 sky130_fd_sc_hd__diode_2 ANTENNA_c691_Q (.DIODE(net556));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge769_B1 (.DIODE(net657));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_SCD (.DIODE(net657));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_B1_N (.DIODE(net657));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_A3 (.DIODE(net657));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_A4 (.DIODE(net657));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_A2 (.DIODE(net657));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_S1 (.DIODE(net657));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_A2 (.DIODE(net657));
 sky130_fd_sc_hd__diode_2 ANTENNA_c295_A1 (.DIODE(net657));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge801_Q (.DIODE(net668));
 sky130_fd_sc_hd__diode_2 ANTENNA_c365_A3 (.DIODE(net668));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_A3 (.DIODE(net668));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_B1_N (.DIODE(net668));
 sky130_fd_sc_hd__diode_2 ANTENNA_c297_B1_N (.DIODE(net668));
 sky130_fd_sc_hd__diode_2 ANTENNA_c295_A2 (.DIODE(net668));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_S0 (.DIODE(net668));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_B1 (.DIODE(net668));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_SCE (.DIODE(net668));
 sky130_fd_sc_hd__diode_2 ANTENNA_c279_B1 (.DIODE(net668));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge840_B (.DIODE(net669));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge802_Y (.DIODE(net669));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone13_A (.DIODE(net1096));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer5_A (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout175_A (.DIODE(net1096));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_A4 (.DIODE(net1096));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_X (.DIODE(net1096));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge836_SCE (.DIODE(net686));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge815_Y (.DIODE(net686));
 sky130_fd_sc_hd__diode_2 ANTENNA_c253_A1 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_c243_A0 (.DIODE(net1091));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_B1 (.DIODE(net1091));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_S0 (.DIODE(net1091));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_S1 (.DIODE(net1091));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_A0 (.DIODE(net1091));
 sky130_fd_sc_hd__diode_2 ANTENNA_c143_A4 (.DIODE(net1091));
 sky130_fd_sc_hd__diode_2 ANTENNA_c140_A2 (.DIODE(net1091));
 sky130_fd_sc_hd__diode_2 ANTENNA_c138_A2 (.DIODE(net1091));
 sky130_fd_sc_hd__diode_2 ANTENNA_c136_A2 (.DIODE(net1091));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_X (.DIODE(net1091));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge829_Q_N (.DIODE(net699));
 sky130_fd_sc_hd__diode_2 ANTENNA_c747_S0 (.DIODE(net699));
 sky130_fd_sc_hd__diode_2 ANTENNA_c724_A3 (.DIODE(net699));
 sky130_fd_sc_hd__diode_2 ANTENNA_c78_A3 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_c70_B1_N (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_c69_X (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_A0 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_A2 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_A0 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_A1 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_c216_A3 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_c203_A4 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone15_A (.DIODE(net1097));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer8_A (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout161_A (.DIODE(net1097));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout160_A (.DIODE(net1097));
 sky130_fd_sc_hd__diode_2 ANTENNA_c134_X (.DIODE(net1097));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge831_Q (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA_c395_A4 (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA_c394_S0 (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA_c393_S0 (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA_c109_S1 (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA_c108_S1 (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA_c107_A4 (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge870_D (.DIODE(net711));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge840_Y (.DIODE(net711));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge844_Q (.DIODE(net716));
 sky130_fd_sc_hd__diode_2 ANTENNA_c762_A3 (.DIODE(net716));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A3 (.DIODE(net716));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_S0 (.DIODE(net716));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_A3 (.DIODE(net716));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_A3 (.DIODE(net716));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_S0 (.DIODE(net716));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge845_Q (.DIODE(net717));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_A2 (.DIODE(net717));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_A3 (.DIODE(net717));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_S0 (.DIODE(net717));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_A2 (.DIODE(net717));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge849_Q_N (.DIODE(net722));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_S1 (.DIODE(net722));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_S0 (.DIODE(net722));
 sky130_fd_sc_hd__diode_2 ANTENNA_c633_S1 (.DIODE(net722));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge850_Q (.DIODE(net724));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_S0 (.DIODE(net724));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_A2 (.DIODE(net724));
 sky130_fd_sc_hd__diode_2 ANTENNA_c746_A3 (.DIODE(net724));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_S1 (.DIODE(net724));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_A3 (.DIODE(net724));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_A3 (.DIODE(net724));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge851_Q (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA_c744_S0 (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA_c739_A1 (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_A2 (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_S1 (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA_c373_A3 (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_A2 (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge853_Q_N (.DIODE(net727));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_A3 (.DIODE(net727));
 sky130_fd_sc_hd__diode_2 ANTENNA_c350_A3 (.DIODE(net727));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_A0 (.DIODE(net727));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge855_Q (.DIODE(net732));
 sky130_fd_sc_hd__diode_2 ANTENNA_c252_S1 (.DIODE(net732));
 sky130_fd_sc_hd__diode_2 ANTENNA_c249_A3 (.DIODE(net732));
 sky130_fd_sc_hd__diode_2 ANTENNA_c248_A3 (.DIODE(net732));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge856_Q (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA_c446_A2 (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA_c371_A2 (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_S0 (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_A3 (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge861_Q (.DIODE(net737));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_S0 (.DIODE(net737));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_S1 (.DIODE(net737));
 sky130_fd_sc_hd__diode_2 ANTENNA_c549_S1 (.DIODE(net737));
 sky130_fd_sc_hd__diode_2 ANTENNA_c541_A (.DIODE(net737));
 sky130_fd_sc_hd__diode_2 ANTENNA_c535_A (.DIODE(net737));
 sky130_fd_sc_hd__diode_2 ANTENNA_c533_A (.DIODE(net737));
 sky130_fd_sc_hd__diode_2 ANTENNA_c531_A (.DIODE(net737));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge772_A3 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_S1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_A4 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_B1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_c143_A2 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_A2 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_S0 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_A1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_c138_X (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge863_Q (.DIODE(net740));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_A3 (.DIODE(net740));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_RESET_B (.DIODE(net740));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_A2 (.DIODE(net740));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_A3 (.DIODE(net740));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge864_Q (.DIODE(net741));
 sky130_fd_sc_hd__diode_2 ANTENNA_c763_A3 (.DIODE(net741));
 sky130_fd_sc_hd__diode_2 ANTENNA_c759_S0 (.DIODE(net741));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_S1 (.DIODE(net741));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_A3 (.DIODE(net741));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_A2 (.DIODE(net741));
 sky130_fd_sc_hd__diode_2 ANTENNA_c698_S1 (.DIODE(net741));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge869_Q_N (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA_c760_A3 (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_A3 (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_A3 (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge873_Q (.DIODE(net751));
 sky130_fd_sc_hd__diode_2 ANTENNA_c743_S1 (.DIODE(net751));
 sky130_fd_sc_hd__diode_2 ANTENNA_c742_S0 (.DIODE(net751));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_S0 (.DIODE(net751));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_A3 (.DIODE(net751));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_A3 (.DIODE(net751));
 sky130_fd_sc_hd__diode_2 ANTENNA_c723_A3 (.DIODE(net751));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_A3 (.DIODE(net751));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_A2 (.DIODE(net751));
 sky130_fd_sc_hd__diode_2 ANTENNA_s876_Q (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA_c257_A3 (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA_c226_S0 (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA_c118_B1 (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold30_A (.DIODE(net757));
 sky130_fd_sc_hd__diode_2 ANTENNA_s877_Q_N (.DIODE(net757));
 sky130_fd_sc_hd__diode_2 ANTENNA_c566_A3 (.DIODE(net757));
 sky130_fd_sc_hd__diode_2 ANTENNA_c556_B1 (.DIODE(net757));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_A3 (.DIODE(net757));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_S1 (.DIODE(net757));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_B1 (.DIODE(net757));
 sky130_fd_sc_hd__diode_2 ANTENNA_s877_Q (.DIODE(net758));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_S0 (.DIODE(net758));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_S0 (.DIODE(net758));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_S0 (.DIODE(net758));
 sky130_fd_sc_hd__diode_2 ANTENNA_c446_B1 (.DIODE(net758));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_S0 (.DIODE(net758));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_S1 (.DIODE(net758));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge771_A4 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_A1 (.DIODE(net1093));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_A0 (.DIODE(net1093));
 sky130_fd_sc_hd__diode_2 ANTENNA_c562_A4 (.DIODE(net1094));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_B1 (.DIODE(net1094));
 sky130_fd_sc_hd__diode_2 ANTENNA_c313_A3 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_c159_S0 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_A1 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_A3 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_c140_X (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold35_A (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_s885_Q_N (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_S1 (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_A3 (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_S0 (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_c259_A2 (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_c242_S1 (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_c239_A1 (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_c229_S0 (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_S1 (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_S1 (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_s887_Q (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_A2 (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_S0 (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_A3 (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_S0 (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA_c371_A3 (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_S0 (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_S0 (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA_c230_S1 (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA_s888_Q (.DIODE(net769));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_A3 (.DIODE(net769));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_A2 (.DIODE(net769));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_S0 (.DIODE(net769));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_S1 (.DIODE(net769));
 sky130_fd_sc_hd__diode_2 ANTENNA_c241_S1 (.DIODE(net769));
 sky130_fd_sc_hd__diode_2 ANTENNA_c239_A3 (.DIODE(net769));
 sky130_fd_sc_hd__diode_2 ANTENNA_c236_S0 (.DIODE(net769));
 sky130_fd_sc_hd__diode_2 ANTENNA_c235_S0 (.DIODE(net769));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_S1 (.DIODE(net769));
 sky130_fd_sc_hd__diode_2 ANTENNA_s889_Q (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c502_A3 (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_A3 (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_S1 (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_S0 (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c236_S1 (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c235_S1 (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c234_S1 (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c231_S1 (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_s890_Q (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_S0 (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_A2 (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_A3 (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_A2 (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_A3 (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_c239_S0 (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_c238_S1 (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_c237_S1 (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_s895_Q (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_A3 (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_S1 (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_S1 (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_B1 (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_S1 (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_S1 (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_c286_B1 (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net779_A (.DIODE(net779));
 sky130_fd_sc_hd__diode_2 ANTENNA_s898_GCLK (.DIODE(net779));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone12_A (.DIODE(net1095));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer6_A (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout145_A (.DIODE(net1095));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_S0 (.DIODE(net1095));
 sky130_fd_sc_hd__diode_2 ANTENNA_c693_A3 (.DIODE(net1095));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_X (.DIODE(net1095));
 sky130_fd_sc_hd__diode_2 ANTENNA_s900_Q_N (.DIODE(net781));
 sky130_fd_sc_hd__diode_2 ANTENNA_c371_S0 (.DIODE(net781));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_S0 (.DIODE(net781));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_S0 (.DIODE(net781));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_S1 (.DIODE(net781));
 sky130_fd_sc_hd__diode_2 ANTENNA_s900_Q (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_S0 (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_A3 (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_S1 (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_S1 (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_S1 (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_s901_Q_N (.DIODE(net783));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_A3 (.DIODE(net783));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_S0 (.DIODE(net783));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_S1 (.DIODE(net783));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_B1 (.DIODE(net783));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_S1 (.DIODE(net783));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold27_A (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_s903_Q (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_S1 (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_S1 (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_A3 (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_S0 (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_S0 (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_S1 (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_s904_Q (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_A2 (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_S0 (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_S1 (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_S0 (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_S1 (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c364_S1 (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c350_S0 (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_s906_Q (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_S0 (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_S1 (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_A2 (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_S0 (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_B1 (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_s912_Q (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_S0 (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_A3 (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA_c373_S0 (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA_c369_S1 (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_S1 (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA_c218_A0 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_S1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_A3 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_A3 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_A2 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_B1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_c148_A3 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_B1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_A3 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_X (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_s916_Q_N (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_S1 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_S0 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_S0 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold32_A (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_s916_Q (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_A3 (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_A2 (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_s921_Q (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_S0 (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_A3 (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_S0 (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_S1 (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_B1 (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_S1 (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_S1 (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_s922_Q (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_S0 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_S0 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_S1 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_S1 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_SET_B (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_s927_Q (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c760_S0 (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_S0 (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_A3 (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A3 (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_S1 (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c482_S1 (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_s928_Q (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_S0 (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_A3 (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_S1 (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_S1 (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_c502_S0 (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_c494_A3 (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_s934_Q (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_S0 (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_A2 (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_S1 (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_s935_Q (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_S1 (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_c582_A3 (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_S1 (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_c558_B1 (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_c547_S1 (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_c546_S1 (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_s937_Q (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_A3 (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_S0 (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_S0 (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_A3 (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_S1 (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_S0 (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_s940_Q_N (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_S0 (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_S1 (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_c582_S0 (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_S1 (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge765_A1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_c270_B1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_A2 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_A0 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_X (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_s943_Q (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_S1 (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c614_S0 (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_S0 (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_S1 (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_S1 (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_S1 (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_S1 (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c586_S1 (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_s944_Q (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c763_S0 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c757_S0 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_S1 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_S0 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_S0 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_A2 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_S0 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_S0 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_s949_Q (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_c747_S1 (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_S0 (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_S1 (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_S1 (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout162_A (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_S1 (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_S0 (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_s952_Q (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_s953_Q (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_c759_S1 (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_c739_A3 (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_S1 (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_S0 (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_c723_S0 (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_A3 (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_S0 (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_S0 (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_c701_S0 (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_c685_S1 (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_s955_Q (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c757_S1 (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_S1 (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c739_S0 (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_S0 (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_A2 (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c703_S0 (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c702_S1 (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_s956_Q (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_S1 (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_S0 (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_A2 (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_S1 (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_c241_A1 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_c238_A0 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_c232_A2 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_S1 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_c182_A3 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_A3 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_A3 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_X (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge765_A4 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_c403_A1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_A0 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_X (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_A0 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_c267_A1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_A0 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_A2 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_X (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout137_A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_c234_A1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_X (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_c228_A1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_A0 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_c218_A2 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_A3 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_c183_S0 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_c180_A1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_A1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_A2 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_A3 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_X (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout146_A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_A1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_c242_A3 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_c245_A1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_X (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_A0 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_A3 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_A1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_B1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_A2 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_c182_A2 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_A1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_S0 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_A3 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_B1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_X (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone4_A (.DIODE(net1099));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout192_A (.DIODE(net1099));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout189_A (.DIODE(net1099));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_X (.DIODE(net1099));
 sky130_fd_sc_hd__diode_2 ANTENNA_c88_B1_N (.DIODE(net1099));
 sky130_fd_sc_hd__diode_2 ANTENNA_c73_B1 (.DIODE(net1099));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout176_A (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_X (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_A0 (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_A2 (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_S0 (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_X (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_c414_A0 (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_c411_B1 (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_c403_S1 (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_c401_A2 (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_SCE (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_c269_A2 (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_c265_A2 (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_c148_A4 (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_c140_A3 (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_A2 (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_X (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_c180_A0 (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_A2 (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout187_A (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_X (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge766_A2 (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_c90_B1_N (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_c369_A0 (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_X (.DIODE(net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_A0 (.DIODE(net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_c158_A1 (.DIODE(net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_B1 (.DIODE(net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_X (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA_c691_SCD (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_A3 (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA_c286_A1 (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_A2 (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_A2 (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_X (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c77_A3 (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c75_B1 (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_A2 (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c62_S1 (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_A1 (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_SET_B (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c190_A3 (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_A1 (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_B1 (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_X (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_A3 (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_A3 (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_A1 (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_A2 (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_A3 (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_A2 (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_A2 (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_X (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_A2 (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c424_A0 (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_S0 (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_A3 (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c158_S1 (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_X (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c87_A3 (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_A1 (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_A0 (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_A2 (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_A1 (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_SCD (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_A4 (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_A2 (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_A2 (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_B1 (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout186_A (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_X (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_c91_A2 (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_c67_A3 (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_c323_S0 (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_X (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_A1 (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_B1_N (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_A3 (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_input30_X (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c698_S0 (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_S0 (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c582_A2 (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c560_A2 (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_A1 (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c321_A0 (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_A2 (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c286_A3 (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_A2 (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_A2 (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout184_A (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_input32_X (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c94_A2 (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout183_A (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_input35_X (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_A3 (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_A3 (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_A2 (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_input37_X (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c764_S1 (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_A2 (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_A0 (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_A2 (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_A3 (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c430_A2 (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_A0 (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_A1 (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_A2 (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_input38_X (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_A0 (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_A2 (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_B1 (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_input41_X (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_c90_A2 (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_c69_A4 (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_c64_S1 (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_c63_A2 (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_c107_A1 (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout180_A (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout179_A (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_input44_X (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_input49_X (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c76_A2 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c68_A1 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c67_B1 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_A0 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_A2 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_A3 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_A1 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c313_A2 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c229_A1 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_input50_X (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_c64_A2 (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_c208_A1 (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_c205_A0 (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_A1 (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_B1 (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_input54_X (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA_c62_A1 (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_B1 (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_A1 (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_S0 (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA_c232_A0 (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA_c222_A2 (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_SCD (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_A2 (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout178_A (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout177_A (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_input59_X (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout167_A (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_s896_Q (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_A3 (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_output66_A (.DIODE(net925));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_A3 (.DIODE(net925));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_S0 (.DIODE(net925));
 sky130_fd_sc_hd__diode_2 ANTENNA_c563_D (.DIODE(net925));
 sky130_fd_sc_hd__diode_2 ANTENNA_c559_Q (.DIODE(net925));
 sky130_fd_sc_hd__diode_2 ANTENNA_output67_A (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_A3 (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_A3 (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_c250_S0 (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_c244_A1 (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_c229_A2 (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_A2 (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_c226_A0 (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_A1 (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_c222_X (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_output69_A (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_A3 (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_A2 (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_A2 (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_A3 (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_A1 (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_A2 (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c586_A0 (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c543_A3 (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c531_X (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_output70_A (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_s885_Q (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_A3 (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_A2 (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_A3 (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_A3 (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_A3 (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c256_A3 (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c249_S1 (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c240_S0 (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_A3 (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_output71_A (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_A1 (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_A3 (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_A2 (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_c365_A1 (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_A1 (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_X (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_output72_A (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_A1 (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_A3 (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_c566_X (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_output73_A (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_A0 (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_A0 (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_A1 (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_Q (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_output74_A (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_s948_Q (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_S1 (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_S0 (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net934_A (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c536_X (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_output77_A (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_s939_Q (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_S0 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_S1 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c586_A3 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_S0 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c571_S1 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout164_A (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_s920_Q (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_A2 (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_S1 (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_A3 (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_S1 (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_output81_A (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_A2 (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_A0 (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_A3 (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_A3 (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_X (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_output83_A (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c392_A0 (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c125_A2 (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c122_A3 (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c120_B1 (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c117_A2 (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c113_Q (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_output84_A (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c88_X (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_A3 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c496_A2 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_A1 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c243_S0 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c121_B1_N (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c113_SET_B (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c104_A4 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net946_A (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_X (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_output91_A (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_A2 (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_A0 (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_A0 (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_RESET_B (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_A1 (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_A2 (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_X (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout163_A (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_output92_A (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_s923_Q (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_S1 (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_S1 (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_output94_A (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge828_Q (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_S0 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_A3 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_S1 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_output96_A (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge874_Q (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_A3 (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_A1 (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_A2 (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_output101_A (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge799_Q (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c392_S0 (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c247_A3 (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c240_A3 (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_output102_A (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge859_Q (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c370_A3 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c366_S1 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c364_A2 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c238_S0 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c235_A2 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_A2 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c220_S1 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_output103_A (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge872_Q (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_A3 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_S0 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_A2 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_A3 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_A1 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_A2 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_SCE (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout168_A (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_output104_A (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_s878_Q (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c393_S1 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_A2 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c251_S1 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_output107_A (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_s880_Q (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_S0 (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_S0 (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c258_A3 (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c247_S0 (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c246_S1 (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c245_S1 (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c234_A3 (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_A3 (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_S0 (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_output108_A (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_D (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c247_A2 (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c128_B1 (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c113_RESET_B (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c109_A2 (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c108_X (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_output111_A (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_s908_Q (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_S1 (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_c344_S1 (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_output116_A (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge773_A1 (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_SCD (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c344_A1 (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_A1 (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_S0 (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_A2 (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_X (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_output117_A (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_s901_Q (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_S0 (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_A3 (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_A3 (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_S1 (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_output119_A (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_s926_Q (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_A3 (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_S1 (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_S1 (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_S0 (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_c482_S0 (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_S1 (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_S1 (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout121_X (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_A1 (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_A3 (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_S0 (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge770_A3 (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge769_A2 (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c434_A3 (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_SCD (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c428_RESET_B (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_A3 (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c278_S0 (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout122_X (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_c742_A2 (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A2 (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_A2 (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_A1 (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_A2 (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_c663_A3 (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_c557_A1 (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_c538_SCD (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_c532_A2 (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_c530_A1 (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout123_X (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c528_B1_N (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c416_S0 (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c415_A3 (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c411_A4 (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c412_S1 (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge775_A1 (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge767_A2 (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c668_A3 (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c667_A1 (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c662_B1_N (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout124_X (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_S0 (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_A1 (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_S0 (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c696_A3 (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c695_A3 (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_A1 (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_S0 (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_A3 (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c686_A1 (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_A2 (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout126_X (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_A1 (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c431_S0 (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c434_S0 (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_A3 (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout124_A (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout125_A (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout127_X (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_c410_A2 (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_c409_A1 (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_c408_B1 (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_A2 (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_c564_A4 (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_c563_SCE (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_A1 (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_A2 (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_c549_A1 (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_c544_S0 (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout129_X (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_A3 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_S0 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_A3 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A3 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_A0 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_A1 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_A1 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_A2 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_A1 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_A1 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout130_X (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_A2 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c416_A3 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c412_A0 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_A0 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_A2 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_SET_B (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c278_A3 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c275_B1_N (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c274_B1_N (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c273_B (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout131_X (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_A1 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_A1 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge772_A2 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c532_A3 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_A2 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c402_B1 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_A3 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_SCD (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c273_A (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c427_RESET_B (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout132_X (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_A1 (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_A0 (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_A0 (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c587_A2 (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_A2 (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout133_X (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_S1 (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_A3 (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_A2 (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_A2 (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_A3 (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_A1 (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_A2 (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c720_A1 (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_A1 (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_A1 (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout134_X (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_S0 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_A3 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_A1 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_A0 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c760_A0 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_A3 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout133_A (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout135_X (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c402_A1 (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c404_A2 (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c412_S0 (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c413_A4 (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c528_A2 (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c671_A2 (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c670_A1 (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c667_A2 (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c665_A1 (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c538_RESET_B (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout136_X (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_A0 (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_A0 (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_A2 (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_S0 (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_S0 (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_A2 (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c540_SCD (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c414_A3 (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c413_A3 (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c400_A (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout137_X (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c232_A1 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c221_A0 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_S0 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c205_A3 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_A3 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_A2 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_A2 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c159_A2 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c158_A2 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_A3 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout138_X (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c87_A1 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c761_A1 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_A1 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_A0 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c743_A1 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_A3 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_A1 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_A0 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_A1 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_A2 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout139_X (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c240_A2 (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_B1 (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c220_A1 (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c203_A3 (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c84_A4 (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c85_A3 (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c81_A2 (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c102_SCE (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c87_A2 (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c226_A2 (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout140_X (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c431_A0 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_A2 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c278_A1 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c274_A2 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c276_A3 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c265_B1 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c283_S0 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c270_A3 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c400_B (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_SCD (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout141_X (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c194_A0 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c191_A3 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c368_A0 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_S0 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_A1 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_A1 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_A2 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_A2 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_A1 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c577_S1 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer19_A (.DIODE(net1103));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer18_A (.DIODE(net1103));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer16_A (.DIODE(net1102));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout142_X (.DIODE(net1103));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_A2 (.DIODE(net1103));
 sky130_fd_sc_hd__diode_2 ANTENNA_c267_B1_N (.DIODE(net1103));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_A4 (.DIODE(net1103));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_B1 (.DIODE(net1103));
 sky130_fd_sc_hd__diode_2 ANTENNA_c410_A3 (.DIODE(net1103));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout143_X (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_A4 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_A1 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c264_A (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_A1 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c663_A2 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_S0 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_A1 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_S0 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_S1 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_A2 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout144_X (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c184_A3 (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_S0 (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c180_S0 (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c372_A1 (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c344_A2 (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_S1 (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_A0 (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_A2 (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c764_S0 (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c502_A1 (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout146_X (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_A1 (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_A1 (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_A2 (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_A3 (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_A2 (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_c611_A1 (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_A0 (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_A1 (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_A3 (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_A3 (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone20_A (.DIODE(net1100));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout148_X (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_A1 (.DIODE(net1100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_A2 (.DIODE(net1100));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout147_A (.DIODE(net1100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_A1 (.DIODE(net1100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c399_B1_N (.DIODE(net1100));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout149_X (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_S0 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c370_A2 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_A3 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_A3 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c365_A0 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_A3 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_A1 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_A0 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_A0 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c502_A0 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout150_X (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c99_B1 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c108_S0 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c107_A3 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c103_B1 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c102_SET_B (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c101_B1_N (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c100_B1 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c222_S0 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c231_A3 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c230_A1 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout151_X (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_c98_SCE (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout150_A (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_c366_A2 (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_S0 (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout149_A (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout154_X (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_c744_A0 (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_A3 (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_A1 (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_A2 (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout153_A (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout157_X (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_A2 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_A0 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c720_A0 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_A3 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_A2 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_A3 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_A2 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c686_A3 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c670_S0 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c663_A1 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout158_X (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_A2 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c549_A2 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c544_A0 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c539_A4 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c536_A2 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout159_X (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_A3 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_A2 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_A2 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_SCE (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_A0 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_S0 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_A3 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_A2 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_A1 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_A1 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout160_X (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_A1 (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_A2 (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c228_A3 (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c222_A0 (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c220_S0 (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_A1 (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c205_S0 (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c198_B1 (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_A1 (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c184_S1 (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout162_X (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_S1 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_S1 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_S0 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_B1 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_B1 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c678_B1 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c676_S1 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c672_S1 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_A3 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_A3 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout163_X (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_S1 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_A3 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_A3 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_S0 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_S0 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_S0 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_S1 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_S0 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_S0 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_S0 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout164_X (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_A3 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_S1 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_output80_A (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_S1 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_A3 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c554_B1 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_A4 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_B1_N (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c437_S1 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_S1 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout165_X (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_S1 (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_S1 (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_S1 (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_A3 (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_S0 (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_S0 (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_A3 (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_S0 (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_A2 (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_S0 (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout167_X (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c611_S1 (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_A2 (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_A2 (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_A4 (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_S1 (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_output64_A (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c430_S0 (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_S1 (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c295_B1_N (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_B1_N (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout168_X (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c245_S0 (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c243_S1 (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_A2 (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c458_B1 (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_B1_N (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_S0 (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_S1 (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c191_S1 (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_S1 (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_B1 (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout169_X (.DIODE(net1028));
 sky130_fd_sc_hd__diode_2 ANTENNA_c180_S1 (.DIODE(net1028));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_S1 (.DIODE(net1028));
 sky130_fd_sc_hd__diode_2 ANTENNA_c183_S1 (.DIODE(net1028));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_B1 (.DIODE(net1028));
 sky130_fd_sc_hd__diode_2 ANTENNA_c446_A3 (.DIODE(net1028));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_S0 (.DIODE(net1028));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_S0 (.DIODE(net1028));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_B1 (.DIODE(net1028));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_A4 (.DIODE(net1028));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_SET_B (.DIODE(net1028));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap170_X (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_c720_A3 (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_A1 (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_A3 (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_A3 (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout171_X (.DIODE(net1030));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_S0 (.DIODE(net1030));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_S0 (.DIODE(net1030));
 sky130_fd_sc_hd__diode_2 ANTENNA_c747_A3 (.DIODE(net1030));
 sky130_fd_sc_hd__diode_2 ANTENNA_c743_A3 (.DIODE(net1030));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_S1 (.DIODE(net1030));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_A1 (.DIODE(net1030));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_A1 (.DIODE(net1030));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_A2 (.DIODE(net1030));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_A3 (.DIODE(net1030));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_A3 (.DIODE(net1030));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout172_X (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_S1 (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_S0 (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_S1 (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_B1_N (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_S0 (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_B1_N (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_A4 (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout173_X (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_c119_A3 (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_c118_A1 (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_c116_A2 (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_c89_A2 (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_c85_S0 (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_c81_A3 (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_c76_A1 (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_c74_B1 (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_c73_A4 (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_c68_B1_N (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap174_X (.DIODE(net1033));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_A3 (.DIODE(net1033));
 sky130_fd_sc_hd__diode_2 ANTENNA_c759_A2 (.DIODE(net1033));
 sky130_fd_sc_hd__diode_2 ANTENNA_c742_A0 (.DIODE(net1033));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_A3 (.DIODE(net1033));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_A1 (.DIODE(net1033));
 sky130_fd_sc_hd__diode_2 ANTENNA_c411_A2 (.DIODE(net1033));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout176_X (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA_c236_A1 (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_A4 (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA_c120_A3 (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA_c115_A1 (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_A1 (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A1 (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_A2 (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_A1 (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_A2 (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_B (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout177_X (.DIODE(net1036));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_A3 (.DIODE(net1036));
 sky130_fd_sc_hd__diode_2 ANTENNA_c203_A1 (.DIODE(net1036));
 sky130_fd_sc_hd__diode_2 ANTENNA_c183_A2 (.DIODE(net1036));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_A3 (.DIODE(net1036));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_A1 (.DIODE(net1036));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_A2 (.DIODE(net1036));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_A2 (.DIODE(net1036));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_A3 (.DIODE(net1036));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_A2 (.DIODE(net1036));
 sky130_fd_sc_hd__diode_2 ANTENNA_c372_A3 (.DIODE(net1036));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout179_X (.DIODE(net1038));
 sky130_fd_sc_hd__diode_2 ANTENNA_c180_A2 (.DIODE(net1038));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_A4 (.DIODE(net1038));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_A3 (.DIODE(net1038));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_A0 (.DIODE(net1038));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_A2 (.DIODE(net1038));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_A0 (.DIODE(net1038));
 sky130_fd_sc_hd__diode_2 ANTENNA_c366_A1 (.DIODE(net1038));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_S0 (.DIODE(net1038));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_A3 (.DIODE(net1038));
 sky130_fd_sc_hd__diode_2 ANTENNA_c234_A2 (.DIODE(net1038));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout180_X (.DIODE(net1039));
 sky130_fd_sc_hd__diode_2 ANTENNA_c99_A3 (.DIODE(net1039));
 sky130_fd_sc_hd__diode_2 ANTENNA_c81_B1 (.DIODE(net1039));
 sky130_fd_sc_hd__diode_2 ANTENNA_c69_B1 (.DIODE(net1039));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_A1 (.DIODE(net1039));
 sky130_fd_sc_hd__diode_2 ANTENNA_c215_A2 (.DIODE(net1039));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_S0 (.DIODE(net1039));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout181_X (.DIODE(net1040));
 sky130_fd_sc_hd__diode_2 ANTENNA_c249_A2 (.DIODE(net1040));
 sky130_fd_sc_hd__diode_2 ANTENNA_c243_A3 (.DIODE(net1040));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_A3 (.DIODE(net1040));
 sky130_fd_sc_hd__diode_2 ANTENNA_c131_A1 (.DIODE(net1040));
 sky130_fd_sc_hd__diode_2 ANTENNA_c127_S1 (.DIODE(net1040));
 sky130_fd_sc_hd__diode_2 ANTENNA_c119_A2 (.DIODE(net1040));
 sky130_fd_sc_hd__diode_2 ANTENNA_c482_A1 (.DIODE(net1040));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_A1 (.DIODE(net1040));
 sky130_fd_sc_hd__diode_2 ANTENNA_c368_A1 (.DIODE(net1040));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_A2 (.DIODE(net1040));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout182_X (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_c251_A1 (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout181_A (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_A1 (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_A3 (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_A1 (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_A4 (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout183_X (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_c183_A0 (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_A3 (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_A4 (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_A3 (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_c134_A4 (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_A2 (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_S0 (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_c545_S0 (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_A1 (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout184_X (.DIODE(net1043));
 sky130_fd_sc_hd__diode_2 ANTENNA_c86_S0 (.DIODE(net1043));
 sky130_fd_sc_hd__diode_2 ANTENNA_c231_A0 (.DIODE(net1043));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_A1 (.DIODE(net1043));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_A1 (.DIODE(net1043));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_SCD (.DIODE(net1043));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_B1_N (.DIODE(net1043));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_A3 (.DIODE(net1043));
 sky130_fd_sc_hd__diode_2 ANTENNA_c703_A1 (.DIODE(net1043));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_A2 (.DIODE(net1043));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_A3 (.DIODE(net1043));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout185_X (.DIODE(net1044));
 sky130_fd_sc_hd__diode_2 ANTENNA_c74_A2 (.DIODE(net1044));
 sky130_fd_sc_hd__diode_2 ANTENNA_c253_A0 (.DIODE(net1044));
 sky130_fd_sc_hd__diode_2 ANTENNA_c243_A1 (.DIODE(net1044));
 sky130_fd_sc_hd__diode_2 ANTENNA_c117_A1 (.DIODE(net1044));
 sky130_fd_sc_hd__diode_2 ANTENNA_c114_B1_N (.DIODE(net1044));
 sky130_fd_sc_hd__diode_2 ANTENNA_c105_S1 (.DIODE(net1044));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_S1 (.DIODE(net1044));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_A4 (.DIODE(net1044));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_A1 (.DIODE(net1044));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_A4 (.DIODE(net1044));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout186_X (.DIODE(net1045));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_A3 (.DIODE(net1045));
 sky130_fd_sc_hd__diode_2 ANTENNA_c256_A1 (.DIODE(net1045));
 sky130_fd_sc_hd__diode_2 ANTENNA_c252_A1 (.DIODE(net1045));
 sky130_fd_sc_hd__diode_2 ANTENNA_c246_A3 (.DIODE(net1045));
 sky130_fd_sc_hd__diode_2 ANTENNA_c194_A2 (.DIODE(net1045));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_B1 (.DIODE(net1045));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A0 (.DIODE(net1045));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_A2 (.DIODE(net1045));
 sky130_fd_sc_hd__diode_2 ANTENNA_c685_S0 (.DIODE(net1045));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_A1 (.DIODE(net1045));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout187_X (.DIODE(net1046));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_A3 (.DIODE(net1046));
 sky130_fd_sc_hd__diode_2 ANTENNA_c277_S1 (.DIODE(net1046));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_A2 (.DIODE(net1046));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_A3 (.DIODE(net1046));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_A2 (.DIODE(net1046));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_A1 (.DIODE(net1046));
 sky130_fd_sc_hd__diode_2 ANTENNA_c577_A3 (.DIODE(net1046));
 sky130_fd_sc_hd__diode_2 ANTENNA_c554_A3 (.DIODE(net1046));
 sky130_fd_sc_hd__diode_2 ANTENNA_c549_A0 (.DIODE(net1046));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_A1 (.DIODE(net1046));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout188_X (.DIODE(net1047));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_SET_B (.DIODE(net1047));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_A4 (.DIODE(net1047));
 sky130_fd_sc_hd__diode_2 ANTENNA_c407_B1_N (.DIODE(net1047));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_A1 (.DIODE(net1047));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_A2 (.DIODE(net1047));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_A3 (.DIODE(net1047));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_A3 (.DIODE(net1047));
 sky130_fd_sc_hd__diode_2 ANTENNA_c675_A2 (.DIODE(net1047));
 sky130_fd_sc_hd__diode_2 ANTENNA_c561_A3 (.DIODE(net1047));
 sky130_fd_sc_hd__diode_2 ANTENNA_c556_A2 (.DIODE(net1047));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout189_X (.DIODE(net1048));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A2 (.DIODE(net1048));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_A0 (.DIODE(net1048));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_A2 (.DIODE(net1048));
 sky130_fd_sc_hd__diode_2 ANTENNA_c529_B1_N (.DIODE(net1048));
 sky130_fd_sc_hd__diode_2 ANTENNA_c530_B1_N (.DIODE(net1048));
 sky130_fd_sc_hd__diode_2 ANTENNA_c539_B1 (.DIODE(net1048));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout188_A (.DIODE(net1048));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer10_A (.DIODE(net1050));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone7_A (.DIODE(net1101));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout191_X (.DIODE(net1101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c182_B1 (.DIODE(net1101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_A3 (.DIODE(net1101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_A4 (.DIODE(net1101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_S0 (.DIODE(net1101));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout190_A (.DIODE(net1101));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout192_X (.DIODE(net1051));
 sky130_fd_sc_hd__diode_2 ANTENNA_c69_A2 (.DIODE(net1098));
 sky130_fd_sc_hd__diode_2 ANTENNA_c66_B1_N (.DIODE(net1098));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_A3 (.DIODE(net1098));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout191_A (.DIODE(net1098));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_A3 (.DIODE(net1098));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_15_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_14_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_13_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_12_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_11_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_10_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_9_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_8_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_7_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_6_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_5_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_4_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_3_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_2_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_1_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_0_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_X (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c538_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c540_CLK_N (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c559_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c691_CLK_N (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge825_GATE_N (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge829_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge836_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge847_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge849_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge853_GATE_N (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge854_GATE_N (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge865_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge875_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s935_GATE_N (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s936_GATE_N (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s938_GATE (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s952_GATE_N (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s953_GATE_N (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_0_0_clk_X (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c563_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c565_CLK_N (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge786_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge869_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s937_GATE_N (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s939_SLEEP_B (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s941_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s942_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s954_GATE (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s955_SLEEP_B (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s956_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s957_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s958_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s960_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_1_0_clk_X (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_CLK_N (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_CLK_N (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c428_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge782_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge783_CLK_N (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge801_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge807_GATE_N (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge852_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge861_GATE (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s915_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s916_GATE_N (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s917_GATE_N (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s919_GATE_N (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_2_0_clk_X (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c427_CLK_N (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_CLK_N (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_CLK_N (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_CLK_N (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge805_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge813_GATE_N (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge814_GATE_N (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge842_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s918_GATE (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s920_GATE_N (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s921_GATE_N (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_3_0_clk_X (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge843_CLK_N (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge845_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge848_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge864_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge873_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s944_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s959_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s961_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s962_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s963_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s964_GATE_N (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s965_GATE_N (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s966_GATE (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_4_0_clk_X (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge826_GATE (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge844_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge850_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge851_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge858_GATE_N (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge874_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s948_GATE_N (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s949_GATE_N (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s951_GATE_N (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_5_0_clk_X (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s909_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s922_GATE (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s923_SLEEP_B (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s924_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s927_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s940_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s943_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_6_0_clk_X (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge812_GATE (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge855_GATE (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s930_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s932_GATE_N (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s945_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s946_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s947_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s950_GATE (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_7_0_clk_X (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge795_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge862_GATE (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge868_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s900_GATE_N (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s903_GATE_N (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s904_GATE_N (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s906_GATE (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s907_SLEEP_B (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s908_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s911_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s925_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_9_0_clk_X (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_CLK_N (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_CLK_N (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge838_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge863_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s878_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s880_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s881_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s905_GATE_N (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_11_0_clk_X (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge828_GATE (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge856_GATE (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge859_GATE_N (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge872_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s910_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s914_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s926_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s928_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s929_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_12_0_clk_X (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_CLK_N (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge834_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge857_GATE_N (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s888_GATE_N (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s889_GATE_N (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s890_GATE (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s891_SLEEP_B (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s912_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s913_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s931_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s933_GATE_N (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s934_GATE (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_13_0_clk_X (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c102_CLK_N (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c106_CLK_N (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c98_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge798_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge799_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge811_GATE (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge835_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge866_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge867_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge870_CLK_N (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s876_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s879_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s882_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s883_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_14_0_clk_X (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c113_CLK_N (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c129_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge792_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge831_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge860_GATE (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s884_GATE_N (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s885_GATE_N (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s886_GATE (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s887_GATE_N (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s892_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s893_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s894_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_15_0_clk_X (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net934_A (.DIODE(clknet_0_net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net934_A (.DIODE(clknet_0_net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net934_X (.DIODE(clknet_0_net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c544_A1 (.DIODE(clknet_1_0__leaf_net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_A1 (.DIODE(clknet_1_0__leaf_net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_A3 (.DIODE(clknet_1_0__leaf_net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_output75_A (.DIODE(clknet_1_0__leaf_net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net934_X (.DIODE(clknet_1_0__leaf_net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_A3 (.DIODE(clknet_1_1__leaf_net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_A1 (.DIODE(clknet_1_1__leaf_net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_A2 (.DIODE(clknet_1_1__leaf_net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_A1 (.DIODE(clknet_1_1__leaf_net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_A2 (.DIODE(clknet_1_1__leaf_net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net934_X (.DIODE(clknet_1_1__leaf_net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_S1 (.DIODE(clknet_1_1__leaf_net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_A3 (.DIODE(clknet_1_1__leaf_net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_output68_A (.DIODE(clknet_1_1__leaf_net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net927_X (.DIODE(clknet_1_1__leaf_net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_S0 (.DIODE(clknet_1_0__leaf_net705));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_A4 (.DIODE(clknet_1_0__leaf_net705));
 sky130_fd_sc_hd__diode_2 ANTENNA_c364_A1 (.DIODE(clknet_1_0__leaf_net705));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net705_X (.DIODE(clknet_1_0__leaf_net705));
 sky130_fd_sc_hd__diode_2 ANTENNA_c215_A3 (.DIODE(clknet_1_0__leaf_net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c216_A2 (.DIODE(clknet_1_0__leaf_net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_A2 (.DIODE(clknet_1_0__leaf_net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c220_A3 (.DIODE(clknet_1_0__leaf_net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c366_A3 (.DIODE(clknet_1_0__leaf_net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c372_S0 (.DIODE(clknet_1_0__leaf_net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net946_X (.DIODE(clknet_1_0__leaf_net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_A0 (.DIODE(clknet_1_1__leaf_net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_A2 (.DIODE(clknet_1_1__leaf_net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_A0 (.DIODE(clknet_1_1__leaf_net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_A3 (.DIODE(clknet_1_1__leaf_net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c482_A2 (.DIODE(clknet_1_1__leaf_net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_A3 (.DIODE(clknet_1_1__leaf_net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_A1 (.DIODE(clknet_1_1__leaf_net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_output87_A (.DIODE(clknet_1_1__leaf_net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net946_X (.DIODE(clknet_1_1__leaf_net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_A3 (.DIODE(clknet_1_1__leaf_net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_A2 (.DIODE(clknet_1_1__leaf_net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_c747_A2 (.DIODE(clknet_1_1__leaf_net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net386_X (.DIODE(clknet_1_1__leaf_net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_A0 (.DIODE(clknet_1_0__leaf_net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_A3 (.DIODE(clknet_1_0__leaf_net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_output93_A (.DIODE(clknet_1_0__leaf_net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net952_X (.DIODE(clknet_1_0__leaf_net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_A0 (.DIODE(clknet_1_0__leaf_net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_c218_A1 (.DIODE(clknet_1_0__leaf_net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_A2 (.DIODE(clknet_1_0__leaf_net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_A3 (.DIODE(clknet_1_0__leaf_net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_A2 (.DIODE(clknet_1_0__leaf_net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_A1 (.DIODE(clknet_1_0__leaf_net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net153_X (.DIODE(clknet_1_0__leaf_net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_A0 (.DIODE(clknet_1_1__leaf_net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_A2 (.DIODE(clknet_1_1__leaf_net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_c228_A2 (.DIODE(clknet_1_1__leaf_net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_c230_A2 (.DIODE(clknet_1_1__leaf_net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_c231_A2 (.DIODE(clknet_1_1__leaf_net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_D (.DIODE(clknet_1_1__leaf_net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_c365_A2 (.DIODE(clknet_1_1__leaf_net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_c369_A1 (.DIODE(clknet_1_1__leaf_net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net153_X (.DIODE(clknet_1_1__leaf_net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_S0 (.DIODE(clknet_1_1__leaf_net762));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_S0 (.DIODE(clknet_1_1__leaf_net762));
 sky130_fd_sc_hd__diode_2 ANTENNA_c229_A3 (.DIODE(clknet_1_1__leaf_net762));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_A2 (.DIODE(clknet_1_1__leaf_net762));
 sky130_fd_sc_hd__diode_2 ANTENNA_c365_S1 (.DIODE(clknet_1_1__leaf_net762));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net762_X (.DIODE(clknet_1_1__leaf_net762));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_SET_B (.DIODE(clknet_1_1__leaf_net779));
 sky130_fd_sc_hd__diode_2 ANTENNA_c392_S1 (.DIODE(clknet_1_1__leaf_net779));
 sky130_fd_sc_hd__diode_2 ANTENNA_c394_S1 (.DIODE(clknet_1_1__leaf_net779));
 sky130_fd_sc_hd__diode_2 ANTENNA_c395_B1 (.DIODE(clknet_1_1__leaf_net779));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net779_X (.DIODE(clknet_1_1__leaf_net779));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_A3 (.DIODE(clknet_1_0__leaf_net778));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_B1 (.DIODE(clknet_1_0__leaf_net778));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_A2 (.DIODE(clknet_1_0__leaf_net778));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_A3 (.DIODE(clknet_1_0__leaf_net778));
 sky130_fd_sc_hd__diode_2 ANTENNA_c762_S0 (.DIODE(clknet_1_0__leaf_net778));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net778_X (.DIODE(clknet_1_0__leaf_net778));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_S1 (.DIODE(clknet_1_1__leaf_net778));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_S1 (.DIODE(clknet_1_1__leaf_net778));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_A4 (.DIODE(clknet_1_1__leaf_net778));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_A2 (.DIODE(clknet_1_1__leaf_net778));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_A3 (.DIODE(clknet_1_1__leaf_net778));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net778_X (.DIODE(clknet_1_1__leaf_net778));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_A1 (.DIODE(net1052));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer3_A (.DIODE(net1052));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer2_A (.DIODE(net1052));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer1_X (.DIODE(net1052));
 sky130_fd_sc_hd__diode_2 ANTENNA_c231_A1 (.DIODE(net1055));
 sky130_fd_sc_hd__diode_2 ANTENNA_c242_S0 (.DIODE(net1055));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_S1 (.DIODE(net1055));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_A3 (.DIODE(net1055));
 sky130_fd_sc_hd__diode_2 ANTENNA_c126_A3 (.DIODE(net1055));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone4_X (.DIODE(net1055));
 sky130_fd_sc_hd__diode_2 ANTENNA_c230_A0 (.DIODE(net1056));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_A1 (.DIODE(net1056));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer5_X (.DIODE(net1056));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_A3 (.DIODE(net1063));
 sky130_fd_sc_hd__diode_2 ANTENNA_c403_A2 (.DIODE(net1063));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_A1 (.DIODE(net1063));
 sky130_fd_sc_hd__diode_2 ANTENNA_c286_A2 (.DIODE(net1063));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_A2 (.DIODE(net1063));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone12_X (.DIODE(net1063));
 sky130_fd_sc_hd__diode_2 ANTENNA_c529_A1 (.DIODE(net1065));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer11_A (.DIODE(net1065));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_A3 (.DIODE(net1065));
 sky130_fd_sc_hd__diode_2 ANTENNA_c402_A4 (.DIODE(net1065));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone14_X (.DIODE(net1065));
 sky130_fd_sc_hd__diode_2 ANTENNA_c266_A (.DIODE(net1066));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_A4 (.DIODE(net1066));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_B1_N (.DIODE(net1066));
 sky130_fd_sc_hd__diode_2 ANTENNA_c276_S0 (.DIODE(net1066));
 sky130_fd_sc_hd__diode_2 ANTENNA_c278_S1 (.DIODE(net1066));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone15_X (.DIODE(net1066));
 sky130_fd_sc_hd__diode_2 ANTENNA_c698_A2 (.DIODE(net1067));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer17_A (.DIODE(net1067));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer16_X (.DIODE(net1067));
 sky130_fd_sc_hd__diode_2 ANTENNA_c226_A3 (.DIODE(net1070));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer19_X (.DIODE(net1070));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(net1057));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer4 (.A(net373),
    .X(net1089));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer7 (.A(net1089),
    .X(net1090));
 sky130_fd_sc_hd__a21bo_1 clone8 (.A1(net916),
    .A2(net920),
    .B1_N(net1034),
    .X(net1091));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer12 (.A(net76),
    .X(net1092));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer13 (.A(net1092),
    .X(net1093));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer14 (.A(net1092),
    .X(net1094));
 sky130_fd_sc_hd__a41o_1 clone16 (.A1(net73),
    .A2(net74),
    .A3(net861),
    .A4(net1042),
    .B1(net1058),
    .X(net1095));
 sky130_fd_sc_hd__a21bo_1 clone17 (.A1(net916),
    .A2(net861),
    .B1_N(net1049),
    .X(net1096));
 sky130_fd_sc_hd__a41o_1 clone18 (.A1(net1034),
    .A2(net921),
    .A3(net871),
    .A4(net1042),
    .B1(net920),
    .X(net1097));
 sky130_fd_sc_hd__clkbuf_1 clone19 (.A(net133),
    .X(net1098));
 sky130_fd_sc_hd__clkbuf_1 clone21 (.A(in0),
    .X(net1099));
 sky130_fd_sc_hd__clkbuf_1 clone22 (.A(net72),
    .X(net1100));
 sky130_fd_sc_hd__clkbuf_1 clone23 (.A(net1051),
    .X(net1101));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer24 (.A(net1001),
    .X(net1102));
 sky130_fd_sc_hd__clkbuf_1 clone25 (.A(net81),
    .X(net1103));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_219 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_282 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_267 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_359 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_256 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_301 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_282 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_219 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_143 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_155 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_423 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_255 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_467 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_340 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_443 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_273 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_395 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_275 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_387 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_407 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_441 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_339 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_359 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_282 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_424 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_452 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_47 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_123 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_274 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_484 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_407 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_247 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_86 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_87 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_522 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_130 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_273 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_497 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_227 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_420 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_76 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_170 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_266 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_200 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_450 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_86 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_170 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_466 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_413 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_443 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_488 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_395 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_415 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_131 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_133 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_378 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_440 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_451 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_144 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_359 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_47 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_273 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_443 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_20 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_140 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_452 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_10 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_22 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_87 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_271 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_423 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_356 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_5 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_10 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_227 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_490 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_283 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_423 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_189 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_256 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_395 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_5 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_452 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_553 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_411 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_398 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_499 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_617 ();
endmodule
