module netlist_1 (clk,
    in0,
    in1,
    in10,
    in11,
    in12,
    in13,
    in14,
    in15,
    in16,
    in17,
    in18,
    in19,
    in2,
    in20,
    in21,
    in22,
    in23,
    in24,
    in25,
    in26,
    in27,
    in28,
    in29,
    in3,
    in30,
    in31,
    in32,
    in33,
    in34,
    in35,
    in36,
    in37,
    in38,
    in39,
    in4,
    in40,
    in41,
    in42,
    in43,
    in44,
    in45,
    in46,
    in47,
    in48,
    in49,
    in5,
    in50,
    in51,
    in52,
    in53,
    in54,
    in55,
    in56,
    in57,
    in58,
    in59,
    in6,
    in60,
    in61,
    in62,
    in63,
    in64,
    in65,
    in66,
    in67,
    in68,
    in69,
    in7,
    in70,
    in71,
    in72,
    in73,
    in74,
    in75,
    in76,
    in77,
    in78,
    in79,
    in8,
    in80,
    in81,
    in82,
    in83,
    in84,
    in85,
    in86,
    in87,
    in88,
    in89,
    in9,
    in90,
    in91,
    in92,
    in93,
    in94,
    in95,
    in96,
    in97,
    in98,
    in99,
    out0,
    out1,
    out10,
    out11,
    out12,
    out13,
    out14,
    out15,
    out16,
    out17,
    out18,
    out19,
    out2,
    out20,
    out21,
    out22,
    out23,
    out24,
    out25,
    out26,
    out27,
    out28,
    out29,
    out3,
    out30,
    out31,
    out32,
    out33,
    out34,
    out35,
    out36,
    out37,
    out38,
    out39,
    out4,
    out40,
    out41,
    out42,
    out43,
    out44,
    out45,
    out46,
    out47,
    out48,
    out49,
    out5,
    out50,
    out51,
    out52,
    out53,
    out54,
    out55,
    out56,
    out57,
    out58,
    out59,
    out6,
    out60,
    out61,
    out62,
    out63,
    out64,
    out65,
    out66,
    out67,
    out68,
    out69,
    out7,
    out70,
    out71,
    out72,
    out73,
    out74,
    out75,
    out76,
    out77,
    out78,
    out79,
    out8,
    out80,
    out81,
    out82,
    out83,
    out84,
    out85,
    out86,
    out87,
    out88,
    out89,
    out9,
    out90,
    out91,
    out92,
    out93,
    out94,
    out95,
    out96,
    out97,
    out98,
    out99,
    rst);
 input clk;
 input in0;
 input in1;
 input in10;
 input in11;
 input in12;
 input in13;
 input in14;
 input in15;
 input in16;
 input in17;
 input in18;
 input in19;
 input in2;
 input in20;
 input in21;
 input in22;
 input in23;
 input in24;
 input in25;
 input in26;
 input in27;
 input in28;
 input in29;
 input in3;
 input in30;
 input in31;
 input in32;
 input in33;
 input in34;
 input in35;
 input in36;
 input in37;
 input in38;
 input in39;
 input in4;
 input in40;
 input in41;
 input in42;
 input in43;
 input in44;
 input in45;
 input in46;
 input in47;
 input in48;
 input in49;
 input in5;
 input in50;
 input in51;
 input in52;
 input in53;
 input in54;
 input in55;
 input in56;
 input in57;
 input in58;
 input in59;
 input in6;
 input in60;
 input in61;
 input in62;
 input in63;
 input in64;
 input in65;
 input in66;
 input in67;
 input in68;
 input in69;
 input in7;
 input in70;
 input in71;
 input in72;
 input in73;
 input in74;
 input in75;
 input in76;
 input in77;
 input in78;
 input in79;
 input in8;
 input in80;
 input in81;
 input in82;
 input in83;
 input in84;
 input in85;
 input in86;
 input in87;
 input in88;
 input in89;
 input in9;
 input in90;
 input in91;
 input in92;
 input in93;
 input in94;
 input in95;
 input in96;
 input in97;
 input in98;
 input in99;
 output out0;
 output out1;
 output out10;
 output out11;
 output out12;
 output out13;
 output out14;
 output out15;
 output out16;
 output out17;
 output out18;
 output out19;
 output out2;
 output out20;
 output out21;
 output out22;
 output out23;
 output out24;
 output out25;
 output out26;
 output out27;
 output out28;
 output out29;
 output out3;
 output out30;
 output out31;
 output out32;
 output out33;
 output out34;
 output out35;
 output out36;
 output out37;
 output out38;
 output out39;
 output out4;
 output out40;
 output out41;
 output out42;
 output out43;
 output out44;
 output out45;
 output out46;
 output out47;
 output out48;
 output out49;
 output out5;
 output out50;
 output out51;
 output out52;
 output out53;
 output out54;
 output out55;
 output out56;
 output out57;
 output out58;
 output out59;
 output out6;
 output out60;
 output out61;
 output out62;
 output out63;
 output out64;
 output out65;
 output out66;
 output out67;
 output out68;
 output out69;
 output out7;
 output out70;
 output out71;
 output out72;
 output out73;
 output out74;
 output out75;
 output out76;
 output out77;
 output out78;
 output out79;
 output out8;
 output out80;
 output out81;
 output out82;
 output out83;
 output out84;
 output out85;
 output out86;
 output out87;
 output out88;
 output out89;
 output out9;
 output out90;
 output out91;
 output out92;
 output out93;
 output out94;
 output out95;
 output out96;
 output out97;
 output out98;
 output out99;
 input rst;

 wire net0;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net63;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net64;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net65;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net66;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net67;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net68;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net69;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net7;
 wire net70;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net71;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net72;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net73;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net74;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net75;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net76;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net77;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net84;
 wire net254;
 wire net481;
 wire net608;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_0_net766;
 wire clknet_1_0__leaf_net766;
 wire clknet_1_1__leaf_net766;
 wire clknet_0_net535;
 wire clknet_1_0__leaf_net535;
 wire clknet_1_1__leaf_net535;
 wire clknet_0_net677;
 wire clknet_1_0__leaf_net677;
 wire clknet_1_1__leaf_net677;
 wire clknet_0_net402;
 wire clknet_1_0__leaf_net402;
 wire clknet_1_1__leaf_net402;
 wire clknet_0_net501;
 wire clknet_1_0__leaf_net501;
 wire clknet_1_1__leaf_net501;
 wire clknet_0_net512;
 wire clknet_1_0__leaf_net512;
 wire clknet_1_1__leaf_net512;
 wire clknet_0_net517;
 wire clknet_1_0__leaf_net517;
 wire clknet_1_1__leaf_net517;
 wire clknet_0_net522;
 wire clknet_1_0__leaf_net522;
 wire clknet_1_1__leaf_net522;
 wire clknet_0_net526;
 wire clknet_1_0__leaf_net526;
 wire clknet_1_1__leaf_net526;
 wire clknet_0_net532;
 wire clknet_1_0__leaf_net532;
 wire clknet_1_1__leaf_net532;
 wire clknet_0_net527;
 wire clknet_1_0__leaf_net527;
 wire clknet_1_1__leaf_net527;
 wire clknet_0_net525;
 wire clknet_1_0__leaf_net525;
 wire clknet_1_1__leaf_net525;
 wire clknet_0_net565;
 wire clknet_1_0__leaf_net565;
 wire clknet_1_1__leaf_net565;
 wire clknet_0_net584;
 wire clknet_1_0__leaf_net584;
 wire clknet_1_1__leaf_net584;
 wire clknet_0_net578;
 wire clknet_1_0__leaf_net578;
 wire clknet_1_1__leaf_net578;
 wire clknet_0_net573;
 wire clknet_1_0__leaf_net573;
 wire clknet_1_1__leaf_net573;
 wire clknet_0_net571;
 wire clknet_1_0__leaf_net571;
 wire clknet_1_1__leaf_net571;
 wire clknet_0_net675;
 wire clknet_1_0__leaf_net675;
 wire clknet_1_1__leaf_net675;
 wire clknet_0_net556;
 wire clknet_1_0__leaf_net556;
 wire clknet_1_1__leaf_net556;
 wire clknet_0_net559;
 wire clknet_1_0__leaf_net559;
 wire clknet_1_1__leaf_net559;
 wire clknet_0_net562;
 wire clknet_1_0__leaf_net562;
 wire clknet_1_1__leaf_net562;
 wire clknet_0_net564;
 wire clknet_1_0__leaf_net564;
 wire clknet_1_1__leaf_net564;
 wire clknet_0_net566;
 wire clknet_1_0__leaf_net566;
 wire clknet_1_1__leaf_net566;
 wire clknet_0_net560;
 wire clknet_1_0__leaf_net560;
 wire clknet_1_1__leaf_net560;
 wire clknet_0_net555;
 wire clknet_1_0__leaf_net555;
 wire clknet_1_1__leaf_net555;
 wire clknet_0_net541;
 wire clknet_1_0__leaf_net541;
 wire clknet_1_1__leaf_net541;
 wire clknet_0_net540;
 wire clknet_1_0__leaf_net540;
 wire clknet_1_1__leaf_net540;
 wire clknet_0_net550;
 wire clknet_1_0__leaf_net550;
 wire clknet_1_1__leaf_net550;
 wire clknet_0_net531;
 wire clknet_1_0__leaf_net531;
 wire clknet_1_1__leaf_net531;
 wire clknet_0_net524;
 wire clknet_1_0__leaf_net524;
 wire clknet_1_1__leaf_net524;
 wire clknet_0_net523;
 wire clknet_1_0__leaf_net523;
 wire clknet_1_1__leaf_net523;
 wire clknet_0_net515;
 wire clknet_1_0__leaf_net515;
 wire clknet_1_1__leaf_net515;
 wire clknet_0_net514;
 wire clknet_1_0__leaf_net514;
 wire clknet_1_1__leaf_net514;
 wire clknet_0_net513;
 wire clknet_1_0__leaf_net513;
 wire clknet_1_1__leaf_net513;
 wire clknet_0_net510;
 wire clknet_1_0__leaf_net510;
 wire clknet_1_1__leaf_net510;
 wire clknet_0_net509;
 wire clknet_1_0__leaf_net509;
 wire clknet_1_1__leaf_net509;
 wire clknet_0_net511;
 wire clknet_1_0__leaf_net511;
 wire clknet_1_1__leaf_net511;
 wire clknet_0_net508;
 wire clknet_1_0__leaf_net508;
 wire clknet_1_1__leaf_net508;
 wire clknet_0_net521;
 wire clknet_1_0__leaf_net521;
 wire clknet_1_1__leaf_net521;
 wire clknet_0_net518;
 wire clknet_1_0__leaf_net518;
 wire clknet_1_1__leaf_net518;
 wire clknet_0_net520;
 wire clknet_1_0__leaf_net520;
 wire clknet_1_1__leaf_net520;
 wire clknet_0_net519;
 wire clknet_1_0__leaf_net519;
 wire clknet_1_1__leaf_net519;
 wire clknet_0_net507;
 wire clknet_1_0__leaf_net507;
 wire clknet_1_1__leaf_net507;
 wire clknet_0_net506;
 wire clknet_1_0__leaf_net506;
 wire clknet_1_1__leaf_net506;
 wire clknet_0_net505;
 wire clknet_1_0__leaf_net505;
 wire clknet_1_1__leaf_net505;
 wire clknet_0_net504;
 wire clknet_1_0__leaf_net504;
 wire clknet_1_1__leaf_net504;
 wire clknet_0_net503;
 wire clknet_1_0__leaf_net503;
 wire clknet_1_1__leaf_net503;
 wire clknet_0_net502;
 wire clknet_1_0__leaf_net502;
 wire clknet_1_1__leaf_net502;
 wire clknet_0_net765;
 wire clknet_1_0__leaf_net765;
 wire clknet_1_1__leaf_net765;
 wire clknet_0_net878;
 wire clknet_1_0__leaf_net878;
 wire clknet_1_1__leaf_net878;
 wire clknet_0_net595;
 wire clknet_1_0__leaf_net595;
 wire clknet_1_1__leaf_net595;
 wire clknet_0_net604;
 wire clknet_1_0__leaf_net604;
 wire clknet_1_1__leaf_net604;
 wire clknet_0_net707;
 wire clknet_1_0__leaf_net707;
 wire clknet_1_1__leaf_net707;
 wire clknet_0_net601;
 wire clknet_1_0__leaf_net601;
 wire clknet_1_1__leaf_net601;
 wire clknet_0_net888;
 wire clknet_1_0__leaf_net888;
 wire clknet_1_1__leaf_net888;
 wire clknet_0_net600;
 wire clknet_1_0__leaf_net600;
 wire clknet_1_1__leaf_net600;
 wire clknet_0_net599;
 wire clknet_1_0__leaf_net599;
 wire clknet_1_1__leaf_net599;
 wire clknet_0_net598;
 wire clknet_1_0__leaf_net598;
 wire clknet_1_1__leaf_net598;
 wire clknet_0_net597;
 wire clknet_1_0__leaf_net597;
 wire clknet_1_1__leaf_net597;
 wire clknet_0_net596;
 wire clknet_1_0__leaf_net596;
 wire clknet_1_1__leaf_net596;
 wire clknet_0_net593;
 wire clknet_1_0__leaf_net593;
 wire clknet_1_1__leaf_net593;
 wire clknet_0_net594;
 wire clknet_1_0__leaf_net594;
 wire clknet_1_1__leaf_net594;
 wire clknet_0_net592;
 wire clknet_1_0__leaf_net592;
 wire clknet_1_1__leaf_net592;
 wire clknet_0_net488;
 wire clknet_1_0__leaf_net488;
 wire clknet_1_1__leaf_net488;
 wire clknet_0_net491;
 wire clknet_1_0__leaf_net491;
 wire clknet_1_1__leaf_net491;
 wire clknet_0_net492;
 wire clknet_1_0__leaf_net492;
 wire clknet_1_1__leaf_net492;
 wire clknet_0_net490;
 wire clknet_1_0__leaf_net490;
 wire clknet_1_1__leaf_net490;
 wire clknet_0_net489;
 wire clknet_1_0__leaf_net489;
 wire clknet_1_1__leaf_net489;
 wire clknet_0_net877;
 wire clknet_1_0__leaf_net877;
 wire clknet_1_1__leaf_net877;
 wire clknet_0_net486;
 wire clknet_1_0__leaf_net486;
 wire clknet_1_1__leaf_net486;
 wire clknet_0_net487;
 wire clknet_1_0__leaf_net487;
 wire clknet_1_1__leaf_net487;
 wire clknet_0_net880;
 wire clknet_1_0__leaf_net880;
 wire clknet_1_1__leaf_net880;
 wire clknet_0_net484;
 wire clknet_1_0__leaf_net484;
 wire clknet_1_1__leaf_net484;
 wire clknet_0_net483;
 wire clknet_1_0__leaf_net483;
 wire clknet_1_1__leaf_net483;
 wire clknet_0_net764;
 wire clknet_1_0__leaf_net764;
 wire clknet_1_1__leaf_net764;
 wire clknet_0_net884;
 wire clknet_1_0__leaf_net884;
 wire clknet_1_1__leaf_net884;
 wire clknet_0_net473;
 wire clknet_1_0__leaf_net473;
 wire clknet_1_1__leaf_net473;
 wire clknet_0_net628;
 wire clknet_1_0__leaf_net628;
 wire clknet_1_1__leaf_net628;
 wire clknet_0_net747;
 wire clknet_1_0__leaf_net747;
 wire clknet_1_1__leaf_net747;
 wire clknet_0_net746;
 wire clknet_1_0__leaf_net746;
 wire clknet_1_1__leaf_net746;
 wire clknet_0_net327;
 wire clknet_1_0__leaf_net327;
 wire clknet_1_1__leaf_net327;
 wire clknet_0_net891;
 wire clknet_1_0__leaf_net891;
 wire clknet_1_1__leaf_net891;
 wire clknet_0_net729;
 wire clknet_1_0__leaf_net729;
 wire clknet_1_1__leaf_net729;
 wire clknet_0_net219;
 wire clknet_1_0__leaf_net219;
 wire clknet_1_1__leaf_net219;
 wire clknet_0_net451;
 wire clknet_1_0__leaf_net451;
 wire clknet_1_1__leaf_net451;
 wire clknet_0_net453;
 wire clknet_1_0__leaf_net453;
 wire clknet_1_1__leaf_net453;
 wire clknet_0_net452;
 wire clknet_1_0__leaf_net452;
 wire clknet_1_1__leaf_net452;
 wire clknet_0_net468;
 wire clknet_1_0__leaf_net468;
 wire clknet_1_1__leaf_net468;
 wire clknet_0_net462;
 wire clknet_1_0__leaf_net462;
 wire clknet_1_1__leaf_net462;
 wire clknet_0_net247;
 wire clknet_1_0__leaf_net247;
 wire clknet_1_1__leaf_net247;
 wire clknet_0_net256;
 wire clknet_1_0__leaf_net256;
 wire clknet_1_1__leaf_net256;
 wire clknet_0_net711;
 wire clknet_1_0__leaf_net711;
 wire clknet_1_1__leaf_net711;
 wire clknet_0_net259;
 wire clknet_1_0__leaf_net259;
 wire clknet_1_1__leaf_net259;
 wire clknet_0_net654;
 wire clknet_1_0__leaf_net654;
 wire clknet_1_1__leaf_net654;
 wire clknet_0_net676;
 wire clknet_1_0__leaf_net676;
 wire clknet_1_1__leaf_net676;
 wire clknet_0_net117;
 wire clknet_1_0__leaf_net117;
 wire clknet_1_1__leaf_net117;
 wire clknet_0_net116;
 wire clknet_1_0__leaf_net116;
 wire clknet_1_1__leaf_net116;
 wire clknet_0_net889;
 wire clknet_1_0__leaf_net889;
 wire clknet_1_1__leaf_net889;
 wire clknet_0_net344;
 wire clknet_1_0__leaf_net344;
 wire clknet_1_1__leaf_net344;
 wire clknet_0_net356;
 wire clknet_1_0__leaf_net356;
 wire clknet_1_1__leaf_net356;
 wire clknet_0_net360;
 wire clknet_1_0__leaf_net360;
 wire clknet_1_1__leaf_net360;
 wire clknet_0_net370;
 wire clknet_1_0__leaf_net370;
 wire clknet_1_1__leaf_net370;
 wire clknet_0_net369;
 wire clknet_1_0__leaf_net369;
 wire clknet_1_1__leaf_net369;
 wire clknet_0_net376;
 wire clknet_1_0__leaf_net376;
 wire clknet_1_1__leaf_net376;
 wire clknet_0_net367;
 wire clknet_1_0__leaf_net367;
 wire clknet_1_1__leaf_net367;
 wire clknet_0_net366;
 wire clknet_1_0__leaf_net366;
 wire clknet_1_1__leaf_net366;
 wire clknet_0_net365;
 wire clknet_1_0__leaf_net365;
 wire clknet_1_1__leaf_net365;
 wire clknet_0_net364;
 wire clknet_1_0__leaf_net364;
 wire clknet_1_1__leaf_net364;
 wire clknet_0_net363;
 wire clknet_1_0__leaf_net363;
 wire clknet_1_1__leaf_net363;
 wire clknet_0_net362;
 wire clknet_1_0__leaf_net362;
 wire clknet_1_1__leaf_net362;
 wire clknet_0_net361;
 wire clknet_1_0__leaf_net361;
 wire clknet_1_1__leaf_net361;
 wire clknet_0_net883;
 wire clknet_1_0__leaf_net883;
 wire clknet_1_1__leaf_net883;
 wire clknet_0_net354;
 wire clknet_1_0__leaf_net354;
 wire clknet_1_1__leaf_net354;
 wire clknet_0_net357;
 wire clknet_1_0__leaf_net357;
 wire clknet_1_1__leaf_net357;
 wire clknet_0_net355;
 wire clknet_1_0__leaf_net355;
 wire clknet_1_1__leaf_net355;
 wire clknet_0_net351;
 wire clknet_1_0__leaf_net351;
 wire clknet_1_1__leaf_net351;
 wire clknet_0_net353;
 wire clknet_1_0__leaf_net353;
 wire clknet_1_1__leaf_net353;
 wire clknet_0_net352;
 wire clknet_1_0__leaf_net352;
 wire clknet_1_1__leaf_net352;
 wire clknet_0_net346;
 wire clknet_1_0__leaf_net346;
 wire clknet_1_1__leaf_net346;
 wire clknet_0_net887;
 wire clknet_1_0__leaf_net887;
 wire clknet_1_1__leaf_net887;
 wire clknet_0_net350;
 wire clknet_1_0__leaf_net350;
 wire clknet_1_1__leaf_net350;
 wire clknet_0_net349;
 wire clknet_1_0__leaf_net349;
 wire clknet_1_1__leaf_net349;
 wire clknet_0_net348;
 wire clknet_1_0__leaf_net348;
 wire clknet_1_1__leaf_net348;
 wire clknet_0_net347;
 wire clknet_1_0__leaf_net347;
 wire clknet_1_1__leaf_net347;
 wire clknet_0_net345;
 wire clknet_1_0__leaf_net345;
 wire clknet_1_1__leaf_net345;
 wire clknet_0_net220;
 wire clknet_1_0__leaf_net220;
 wire clknet_1_1__leaf_net220;
 wire clknet_0_net233;
 wire clknet_1_0__leaf_net233;
 wire clknet_1_1__leaf_net233;
 wire clknet_0_net243;
 wire clknet_1_0__leaf_net243;
 wire clknet_1_1__leaf_net243;
 wire clknet_0_net248;
 wire clknet_1_0__leaf_net248;
 wire clknet_1_1__leaf_net248;
 wire clknet_0_net246;
 wire clknet_1_0__leaf_net246;
 wire clknet_1_1__leaf_net246;
 wire clknet_0_net249;
 wire clknet_1_0__leaf_net249;
 wire clknet_1_1__leaf_net249;
 wire clknet_0_net244;
 wire clknet_1_0__leaf_net244;
 wire clknet_1_1__leaf_net244;
 wire clknet_0_net236;
 wire clknet_1_0__leaf_net236;
 wire clknet_1_1__leaf_net236;
 wire clknet_0_net238;
 wire clknet_1_0__leaf_net238;
 wire clknet_1_1__leaf_net238;
 wire clknet_0_net234;
 wire clknet_1_0__leaf_net234;
 wire clknet_1_1__leaf_net234;
 wire clknet_0_net235;
 wire clknet_1_0__leaf_net235;
 wire clknet_1_1__leaf_net235;
 wire clknet_0_net231;
 wire clknet_1_0__leaf_net231;
 wire clknet_1_1__leaf_net231;
 wire clknet_0_net232;
 wire clknet_1_0__leaf_net232;
 wire clknet_1_1__leaf_net232;
 wire clknet_0_net230;
 wire clknet_1_0__leaf_net230;
 wire clknet_1_1__leaf_net230;
 wire clknet_0_net229;
 wire clknet_1_0__leaf_net229;
 wire clknet_1_1__leaf_net229;
 wire clknet_0_net228;
 wire clknet_1_0__leaf_net228;
 wire clknet_1_1__leaf_net228;
 wire clknet_0_net227;
 wire clknet_1_0__leaf_net227;
 wire clknet_1_1__leaf_net227;
 wire clknet_0_net226;
 wire clknet_1_0__leaf_net226;
 wire clknet_1_1__leaf_net226;
 wire clknet_0_net225;
 wire clknet_1_0__leaf_net225;
 wire clknet_1_1__leaf_net225;
 wire clknet_0_net224;
 wire clknet_1_0__leaf_net224;
 wire clknet_1_1__leaf_net224;
 wire clknet_0_net223;
 wire clknet_1_0__leaf_net223;
 wire clknet_1_1__leaf_net223;
 wire clknet_0_net222;
 wire clknet_1_0__leaf_net222;
 wire clknet_1_1__leaf_net222;
 wire clknet_0_net221;
 wire clknet_1_0__leaf_net221;
 wire clknet_1_1__leaf_net221;
 wire clknet_0_net218;
 wire clknet_1_0__leaf_net218;
 wire clknet_1_1__leaf_net218;
 wire clknet_0_net217;
 wire clknet_1_0__leaf_net217;
 wire clknet_1_1__leaf_net217;
 wire clknet_0_net127;
 wire clknet_1_0__leaf_net127;
 wire clknet_1_1__leaf_net127;
 wire clknet_0_net137;
 wire clknet_1_0__leaf_net137;
 wire clknet_1_1__leaf_net137;
 wire clknet_0_net142;
 wire clknet_1_0__leaf_net142;
 wire clknet_1_1__leaf_net142;
 wire clknet_0_net138;
 wire clknet_1_0__leaf_net138;
 wire clknet_1_1__leaf_net138;
 wire clknet_0_net139;
 wire clknet_1_0__leaf_net139;
 wire clknet_1_1__leaf_net139;
 wire clknet_0_net135;
 wire clknet_1_0__leaf_net135;
 wire clknet_1_1__leaf_net135;
 wire clknet_0_net133;
 wire clknet_1_0__leaf_net133;
 wire clknet_1_1__leaf_net133;
 wire clknet_0_net136;
 wire clknet_1_0__leaf_net136;
 wire clknet_1_1__leaf_net136;
 wire clknet_0_net134;
 wire clknet_1_0__leaf_net134;
 wire clknet_1_1__leaf_net134;
 wire clknet_0_net129;
 wire clknet_1_0__leaf_net129;
 wire clknet_1_1__leaf_net129;
 wire clknet_0_net132;
 wire clknet_1_0__leaf_net132;
 wire clknet_1_1__leaf_net132;
 wire clknet_0_net894;
 wire clknet_1_0__leaf_net894;
 wire clknet_1_1__leaf_net894;
 wire clknet_0_net901;
 wire clknet_1_0__leaf_net901;
 wire clknet_1_1__leaf_net901;
 wire clknet_0_net898;
 wire clknet_1_0__leaf_net898;
 wire clknet_1_1__leaf_net898;
 wire clknet_0_net895;
 wire clknet_1_0__leaf_net895;
 wire clknet_1_1__leaf_net895;
 wire clknet_0_net131;
 wire clknet_1_0__leaf_net131;
 wire clknet_1_1__leaf_net131;
 wire clknet_0_net130;
 wire clknet_1_0__leaf_net130;
 wire clknet_1_1__leaf_net130;
 wire clknet_0_net128;
 wire clknet_1_0__leaf_net128;
 wire clknet_1_1__leaf_net128;
 wire clknet_0_net890;
 wire clknet_1_0__leaf_net890;
 wire clknet_1_1__leaf_net890;
 wire clknet_0_net125;
 wire clknet_1_0__leaf_net125;
 wire clknet_1_1__leaf_net125;
 wire clknet_0_net126;
 wire clknet_1_0__leaf_net126;
 wire clknet_1_1__leaf_net126;
 wire clknet_0_net124;
 wire clknet_1_0__leaf_net124;
 wire clknet_1_1__leaf_net124;
 wire clknet_0_net123;
 wire clknet_1_0__leaf_net123;
 wire clknet_1_1__leaf_net123;
 wire clknet_0_net122;
 wire clknet_1_0__leaf_net122;
 wire clknet_1_1__leaf_net122;
 wire clknet_0_net108;
 wire clknet_1_0__leaf_net108;
 wire clknet_1_1__leaf_net108;
 wire clknet_0_net710;
 wire clknet_1_0__leaf_net710;
 wire clknet_1_1__leaf_net710;
 wire clknet_0_net207;
 wire clknet_1_0__leaf_net207;
 wire clknet_1_1__leaf_net207;
 wire clknet_0_net209;
 wire clknet_1_0__leaf_net209;
 wire clknet_1_1__leaf_net209;
 wire clknet_0_net208;
 wire clknet_1_0__leaf_net208;
 wire clknet_1_1__leaf_net208;
 wire clknet_0_net212;
 wire clknet_1_0__leaf_net212;
 wire clknet_1_1__leaf_net212;
 wire clknet_0_net166;
 wire clknet_1_0__leaf_net166;
 wire clknet_1_1__leaf_net166;
 wire clknet_0_net164;
 wire clknet_1_0__leaf_net164;
 wire clknet_1_1__leaf_net164;
 wire clknet_0_net709;
 wire clknet_1_0__leaf_net709;
 wire clknet_1_1__leaf_net709;
 wire clknet_0_net181;
 wire clknet_1_0__leaf_net181;
 wire clknet_1_1__leaf_net181;
 wire clknet_0_net189;
 wire clknet_1_0__leaf_net189;
 wire clknet_1_1__leaf_net189;
 wire clknet_0_net194;
 wire clknet_1_0__leaf_net194;
 wire clknet_1_1__leaf_net194;
 wire clknet_0_net191;
 wire clknet_1_0__leaf_net191;
 wire clknet_1_1__leaf_net191;
 wire clknet_0_net193;
 wire clknet_1_0__leaf_net193;
 wire clknet_1_1__leaf_net193;
 wire clknet_0_net292;
 wire clknet_1_0__leaf_net292;
 wire clknet_1_1__leaf_net292;
 wire clknet_0_net197;
 wire clknet_1_0__leaf_net197;
 wire clknet_1_1__leaf_net197;
 wire clknet_0_net188;
 wire clknet_1_0__leaf_net188;
 wire clknet_1_1__leaf_net188;
 wire clknet_0_net187;
 wire clknet_1_0__leaf_net187;
 wire clknet_1_1__leaf_net187;
 wire clknet_0_net186;
 wire clknet_1_0__leaf_net186;
 wire clknet_1_1__leaf_net186;
 wire clknet_0_net185;
 wire clknet_1_0__leaf_net185;
 wire clknet_1_1__leaf_net185;
 wire clknet_0_net184;
 wire clknet_1_0__leaf_net184;
 wire clknet_1_1__leaf_net184;
 wire clknet_0_net183;
 wire clknet_1_0__leaf_net183;
 wire clknet_1_1__leaf_net183;
 wire clknet_0_net182;
 wire clknet_1_0__leaf_net182;
 wire clknet_1_1__leaf_net182;
 wire clknet_0_net180;
 wire clknet_1_0__leaf_net180;
 wire clknet_1_1__leaf_net180;
 wire clknet_0_net179;
 wire clknet_1_0__leaf_net179;
 wire clknet_1_1__leaf_net179;
 wire clknet_0_net178;
 wire clknet_1_0__leaf_net178;
 wire clknet_1_1__leaf_net178;
 wire clknet_0_net177;
 wire clknet_1_0__leaf_net177;
 wire clknet_1_1__leaf_net177;
 wire clknet_0_net160;
 wire clknet_1_0__leaf_net160;
 wire clknet_1_1__leaf_net160;
 wire clknet_0_net159;
 wire clknet_1_0__leaf_net159;
 wire clknet_1_1__leaf_net159;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;

 sky130_fd_sc_hd__mux4_2 c100 (.A0(net870),
    .A1(net862),
    .A2(net865),
    .A3(net866),
    .S0(net859),
    .S1(net867),
    .X(net0));
 sky130_fd_sc_hd__mux4_1 c101 (.A0(net873),
    .A1(net871),
    .A2(net868),
    .A3(net866),
    .S0(net861),
    .S1(net853),
    .X(net1));
 sky130_fd_sc_hd__mux4_1 c102 (.A0(net872),
    .A1(net867),
    .A2(net844),
    .A3(net854),
    .S0(net862),
    .S1(net866),
    .X(net2));
 sky130_fd_sc_hd__mux4_1 c103 (.A0(net1),
    .A1(net2),
    .A2(net871),
    .A3(net857),
    .S0(net846),
    .S1(net866),
    .X(net3));
 sky130_fd_sc_hd__mux4_2 c104 (.A0(net861),
    .A1(net864),
    .A2(net867),
    .A3(net873),
    .S0(net868),
    .S1(net3),
    .X(net4));
 sky130_fd_sc_hd__mux4_1 c105 (.A0(net869),
    .A1(net0),
    .A2(net867),
    .A3(net861),
    .S0(net866),
    .S1(net873),
    .X(net5));
 sky130_fd_sc_hd__mux4_1 c106 (.A0(net866),
    .A1(net5),
    .A2(net1),
    .A3(net872),
    .S0(net845),
    .S1(net864),
    .X(net6));
 sky130_fd_sc_hd__mux4_1 c107 (.A0(net6),
    .A1(net4),
    .A2(net873),
    .A3(net5),
    .S0(net867),
    .S1(net838),
    .X(net7));
 sky130_fd_sc_hd__mux4_1 c108 (.A0(net3),
    .A1(net868),
    .A2(net871),
    .A3(net6),
    .S0(net7),
    .S1(net5),
    .X(net8));
 sky130_fd_sc_hd__mux4_1 c109 (.A0(net7),
    .A1(net8),
    .A2(net1),
    .A3(net843),
    .S0(net865),
    .S1(net6),
    .X(net9));
 sky130_fd_sc_hd__a41o_1 c110 (.A1(net9),
    .A2(net865),
    .A3(net857),
    .A4(net4),
    .B1(net0),
    .X(net10));
 sky130_fd_sc_hd__a41o_1 c111 (.A1(net916),
    .A2(net9),
    .A3(net844),
    .A4(net839),
    .B1(net865),
    .X(net11));
 sky130_fd_sc_hd__a41o_1 c112 (.A1(net914),
    .A2(net916),
    .A3(net842),
    .A4(net4),
    .B1(net870),
    .X(net12));
 sky130_fd_sc_hd__a41o_1 c113 (.A1(net916),
    .A2(net914),
    .A3(net12),
    .A4(net870),
    .B1(net865),
    .X(net13));
 sky130_fd_sc_hd__a41o_2 c114 (.A1(net865),
    .A2(net13),
    .A3(net914),
    .A4(net12),
    .B1(net916),
    .X(net14));
 sky130_fd_sc_hd__a41o_1 c115 (.A1(net12),
    .A2(net916),
    .A3(net14),
    .A4(net914),
    .B1(net13),
    .X(net15));
 sky130_fd_sc_hd__mux4_2 c116 (.A0(net916),
    .A1(net914),
    .A2(net12),
    .A3(net14),
    .S0(net13),
    .S1(net15),
    .X(net16));
 sky130_fd_sc_hd__mux4_2 c117 (.A0(net14),
    .A1(net15),
    .A2(net914),
    .A3(net16),
    .S0(net916),
    .S1(net12),
    .X(net17));
 sky130_fd_sc_hd__mux4_2 c118 (.A0(net14),
    .A1(net15),
    .A2(net16),
    .A3(net17),
    .S0(net916),
    .S1(net914),
    .X(net18));
 sky130_fd_sc_hd__mux4_2 c119 (.A0(net15),
    .A1(net18),
    .A2(net16),
    .A3(net12),
    .S0(net914),
    .S1(net916),
    .X(net19));
 sky130_fd_sc_hd__mux4_2 c120 (.A0(net842),
    .A1(net19),
    .A2(net16),
    .A3(net18),
    .S0(net14),
    .S1(net10),
    .X(net20));
 sky130_fd_sc_hd__mux4_2 c121 (.A0(net18),
    .A1(net913),
    .A2(net19),
    .A3(net11),
    .S0(net16),
    .S1(net14),
    .X(net21));
 sky130_fd_sc_hd__mux4_1 c122 (.A0(net16),
    .A1(net19),
    .A2(net18),
    .A3(net14),
    .S0(net913),
    .S1(net17),
    .X(net22));
 sky130_fd_sc_hd__mux4_1 c123 (.A0(net13),
    .A1(net19),
    .A2(net21),
    .A3(net18),
    .S0(net913),
    .S1(net16),
    .X(net23));
 sky130_fd_sc_hd__mux4_1 c124 (.A0(net22),
    .A1(net21),
    .A2(net23),
    .A3(net914),
    .S0(net16),
    .S1(net18),
    .X(net24));
 sky130_fd_sc_hd__mux4_2 c125 (.A0(net17),
    .A1(net23),
    .A2(net24),
    .A3(net14),
    .S0(net19),
    .S1(net21),
    .X(net25));
 sky130_fd_sc_hd__mux4_1 c126 (.A0(net19),
    .A1(net913),
    .A2(net25),
    .A3(net24),
    .S0(net18),
    .S1(net22),
    .X(net26));
 sky130_fd_sc_hd__mux4_1 c127 (.A0(net25),
    .A1(net24),
    .A2(net21),
    .A3(net18),
    .S0(net19),
    .S1(net660),
    .X(net27));
 sky130_fd_sc_hd__mux4_1 c128 (.A0(net24),
    .A1(net21),
    .A2(net25),
    .A3(net19),
    .S0(net660),
    .S1(net692),
    .X(net28));
 sky130_fd_sc_hd__mux4_1 c129 (.A0(net916),
    .A1(net21),
    .A2(net25),
    .A3(net636),
    .S0(net660),
    .S1(net692),
    .X(net29));
 sky130_fd_sc_hd__mux4_1 c130 (.A0(net913),
    .A1(net25),
    .A2(net16),
    .A3(net636),
    .S0(net660),
    .S1(net692),
    .X(net30));
 sky130_fd_sc_hd__a41o_1 c131 (.A1(net17),
    .A2(net16),
    .A3(net914),
    .A4(net636),
    .B1(net692),
    .X(net893));
 sky130_fd_sc_hd__mux4_2 c132 (.A0(net797),
    .A1(net782),
    .A2(net784),
    .A3(net781),
    .S0(net778),
    .S1(net863),
    .X(net31));
 sky130_fd_sc_hd__mux4_1 c133 (.A0(net819),
    .A1(net31),
    .A2(net778),
    .A3(net852),
    .S0(net787),
    .S1(net779),
    .X(net32));
 sky130_fd_sc_hd__mux4_2 c134 (.A0(net31),
    .A1(net919),
    .A2(net783),
    .A3(net780),
    .S0(net481),
    .S1(net788),
    .X(net33));
 sky130_fd_sc_hd__mux4_2 c135 (.A0(net919),
    .A1(net33),
    .A2(net779),
    .A3(net31),
    .S0(net852),
    .S1(net786),
    .X(net34));
 sky130_fd_sc_hd__mux4_2 c136 (.A0(net781),
    .A1(net780),
    .A2(net919),
    .A3(net33),
    .S0(net31),
    .S1(net34),
    .X(net35));
 sky130_fd_sc_hd__mux4_2 c137 (.A0(net917),
    .A1(net33),
    .A2(net788),
    .A3(net919),
    .S0(net31),
    .S1(net34),
    .X(net36));
 sky130_fd_sc_hd__mux4_2 c138 (.A0(net917),
    .A1(net34),
    .A2(net919),
    .A3(net254),
    .S0(net784),
    .S1(net36),
    .X(net37));
 sky130_fd_sc_hd__mux4_1 c139 (.A0(net34),
    .A1(net36),
    .A2(net785),
    .A3(net917),
    .S0(net33),
    .S1(net919),
    .X(net38));
 sky130_fd_sc_hd__mux4_1 c140 (.A0(net481),
    .A1(net33),
    .A2(net34),
    .A3(net36),
    .S0(net32),
    .S1(net917),
    .X(net39));
 sky130_fd_sc_hd__mux4_2 c141 (.A0(net37),
    .A1(net38),
    .A2(net36),
    .A3(net31),
    .S0(net919),
    .S1(net33),
    .X(net40));
 sky130_fd_sc_hd__mux4_2 c142 (.A0(net36),
    .A1(net40),
    .A2(net919),
    .A3(net38),
    .S0(net35),
    .S1(net33),
    .X(net41));
 sky130_fd_sc_hd__mux4_2 c143 (.A0(net36),
    .A1(net41),
    .A2(net37),
    .A3(net917),
    .S0(net919),
    .S1(net33),
    .X(net42));
 sky130_fd_sc_hd__mux4_2 c144 (.A0(net33),
    .A1(net917),
    .A2(net841),
    .A3(net36),
    .S0(net608),
    .S1(net42),
    .X(net43));
 sky130_fd_sc_hd__mux4_2 c145 (.A0(net31),
    .A1(net39),
    .A2(net42),
    .A3(net36),
    .S0(net33),
    .S1(net41),
    .X(net44));
 sky130_fd_sc_hd__mux4_2 c146 (.A0(net44),
    .A1(net42),
    .A2(net917),
    .A3(net808),
    .S0(net40),
    .S1(net36),
    .X(net45));
 sky130_fd_sc_hd__mux4_1 c147 (.A0(net863),
    .A1(net44),
    .A2(net42),
    .A3(net45),
    .S0(net917),
    .S1(net919),
    .X(net46));
 sky130_fd_sc_hd__mux4_2 c148 (.A0(net40),
    .A1(net45),
    .A2(net46),
    .A3(net41),
    .S0(net830),
    .S1(net36),
    .X(net47));
 sky130_fd_sc_hd__mux4_1 c149 (.A0(net41),
    .A1(net47),
    .A2(net44),
    .A3(net84),
    .S0(net45),
    .S1(net917),
    .X(net48));
 sky130_fd_sc_hd__mux4_1 c150 (.A0(net45),
    .A1(net48),
    .A2(net38),
    .A3(net47),
    .S0(net42),
    .S1(net917),
    .X(net49));
 sky130_fd_sc_hd__mux4_1 c151 (.A0(net39),
    .A1(net49),
    .A2(net48),
    .A3(net47),
    .S0(net37),
    .S1(net45),
    .X(net50));
 sky130_fd_sc_hd__mux4_2 c152 (.A0(net38),
    .A1(net46),
    .A2(net43),
    .A3(net37),
    .S0(net44),
    .S1(net47),
    .X(net51));
 sky130_fd_sc_hd__mux4_2 c153 (.A0(net50),
    .A1(net47),
    .A2(net39),
    .A3(net51),
    .S0(net49),
    .S1(net48),
    .X(net52));
 sky130_fd_sc_hd__mux4_2 c154 (.A0(net52),
    .A1(net799),
    .A2(net51),
    .A3(net791),
    .S0(net804),
    .S1(net812),
    .X(net53));
 sky130_fd_sc_hd__mux4_1 c155 (.A0(net812),
    .A1(net53),
    .A2(net792),
    .A3(net789),
    .S0(net795),
    .S1(net800),
    .X(net54));
 sky130_fd_sc_hd__mux4_2 c156 (.A0(net53),
    .A1(net811),
    .A2(net910),
    .A3(net798),
    .S0(net809),
    .S1(net807),
    .X(net55));
 sky130_fd_sc_hd__sdfbbn_1 c157 (.CLK_N(clknet_4_4_0_clk),
    .D(net55),
    .RESET_B(net792),
    .SCD(net796),
    .SCE(net53),
    .SET_B(net910),
    .Q(net57),
    .Q_N(net56));
 sky130_fd_sc_hd__mux4_1 c158 (.A0(net57),
    .A1(net804),
    .A2(net55),
    .A3(net910),
    .S0(net52),
    .S1(net53),
    .X(net58));
 sky130_fd_sc_hd__a41o_1 c159 (.A1(net910),
    .A2(net57),
    .A3(net55),
    .A4(net53),
    .B1(net942),
    .X(net59));
 sky130_fd_sc_hd__mux4_2 c160 (.A0(net53),
    .A1(net802),
    .A2(net798),
    .A3(net910),
    .S0(net693),
    .S1(net715),
    .X(net60));
 sky130_fd_sc_hd__mux4_1 c161 (.A0(net60),
    .A1(net55),
    .A2(net56),
    .A3(net910),
    .S0(net693),
    .S1(net715),
    .X(net61));
 sky130_fd_sc_hd__mux4_1 c162 (.A0(net55),
    .A1(net794),
    .A2(net54),
    .A3(net693),
    .S0(net706),
    .X(net62));
 sky130_fd_sc_hd__mux4_1 c163 (.A0(net55),
    .A1(net801),
    .A2(net800),
    .A3(net56),
    .S0(net706),
    .S1(net715),
    .X(net63));
 sky130_fd_sc_hd__a41o_1 c164 (.A1(net60),
    .A2(net56),
    .A3(net910),
    .A4(net715),
    .B1(net946),
    .X(net64));
 sky130_fd_sc_hd__sdfbbn_2 c165 (.CLK_N(clknet_4_1_0_clk),
    .D(net60),
    .RESET_B(net642),
    .SCD(net694),
    .SCE(net715),
    .SET_B(net723),
    .Q(net66),
    .Q_N(net65));
 sky130_fd_sc_hd__mux4_2 c166 (.A0(net910),
    .A1(net57),
    .A2(net66),
    .A3(net803),
    .S0(net790),
    .S1(net722),
    .X(net67));
 sky130_fd_sc_hd__mux4_1 c167 (.A0(net66),
    .A1(net60),
    .A2(net67),
    .A3(net642),
    .S0(net715),
    .S1(net722),
    .X(net68));
 sky130_fd_sc_hd__mux4_2 c168 (.A0(net66),
    .A1(net56),
    .A2(net642),
    .A3(net715),
    .S0(net723),
    .S1(net724),
    .X(net69));
 sky130_fd_sc_hd__mux4_1 c169 (.A0(net910),
    .A1(net69),
    .A2(net67),
    .A3(net807),
    .S0(net65),
    .S1(net945),
    .X(net70));
 sky130_fd_sc_hd__mux4_1 c170 (.A0(net51),
    .A1(net69),
    .A2(net66),
    .A3(net643),
    .S0(net715),
    .S1(net725),
    .X(net71));
 sky130_fd_sc_hd__mux4_1 c171 (.A0(net57),
    .A1(net66),
    .A2(net71),
    .A3(net643),
    .S0(net722),
    .S1(net725),
    .X(net72));
 sky130_fd_sc_hd__mux4_2 c172 (.A0(net57),
    .A1(net69),
    .A2(net910),
    .A3(net643),
    .S0(net723),
    .S1(net724),
    .X(net73));
 sky130_fd_sc_hd__mux4_1 c173 (.A0(net908),
    .A1(net791),
    .A2(net55),
    .A3(net809),
    .S0(net65),
    .S1(net643),
    .X(net74));
 sky130_fd_sc_hd__mux4_1 c174 (.A0(net72),
    .A1(net71),
    .A2(net69),
    .A3(net908),
    .S0(net65),
    .S1(net715),
    .X(net75));
 sky130_fd_sc_hd__mux4_1 c175 (.A0(net69),
    .A1(net908),
    .A2(net789),
    .A3(net787),
    .S0(net65),
    .S1(net706),
    .X(net76));
 sky130_fd_sc_hd__mux4_2 c176 (.A0(net836),
    .A1(net829),
    .A2(net810),
    .A3(net816),
    .S0(net831),
    .S1(net642),
    .X(net77));
 sky130_fd_sc_hd__a41o_2 c177 (.A1(net821),
    .A2(net77),
    .A3(net833),
    .A4(net815),
    .B1(net643),
    .X(net78));
 sky130_fd_sc_hd__mux4_1 c178 (.A0(net77),
    .A1(net831),
    .A2(net78),
    .A3(net836),
    .S0(net908),
    .S1(net820),
    .X(net79));
 sky130_fd_sc_hd__mux4_1 c179 (.A0(net78),
    .A1(net77),
    .A2(net908),
    .A3(net826),
    .S0(net814),
    .S1(net941),
    .X(net80));
 sky130_fd_sc_hd__mux4_1 c180 (.A0(net78),
    .A1(net815),
    .A2(net835),
    .A3(net77),
    .S0(net618),
    .S1(net932),
    .X(net81));
 sky130_fd_sc_hd__mux4_1 c181 (.A0(net813),
    .A1(net78),
    .A2(net805),
    .A3(net908),
    .S0(net77),
    .S1(net932),
    .X(net82));
 sky130_fd_sc_hd__mux4_2 c182 (.A0(net834),
    .A1(net78),
    .A2(net77),
    .A3(net619),
    .S0(net932),
    .S1(net930),
    .X(net83));
 sky130_fd_sc_hd__mux4_2 c183 (.A0(net83),
    .A1(net817),
    .A2(net78),
    .A3(net73),
    .S1(net932),
    .X(net618));
 sky130_fd_sc_hd__mux4_1 c184 (.A0(net81),
    .A1(net83),
    .A2(net823),
    .A3(net619),
    .S0(net932),
    .S1(net930),
    .X(net85));
 sky130_fd_sc_hd__mux4_2 c185 (.A0(net827),
    .A1(net83),
    .A2(net78),
    .A3(net85),
    .S0(net619),
    .S1(net932),
    .X(net86));
 sky130_fd_sc_hd__mux4_1 c186 (.A0(net83),
    .A1(net77),
    .A2(net86),
    .A3(net78),
    .S0(net726),
    .S1(net930),
    .X(net87));
 sky130_fd_sc_hd__mux4_1 c187 (.A0(net77),
    .A1(net86),
    .A2(net83),
    .A3(net824),
    .S0(net619),
    .S1(net930),
    .X(net88));
 sky130_fd_sc_hd__mux4_2 c188 (.A0(net87),
    .A1(net88),
    .A2(net83),
    .A3(net86),
    .S0(net618),
    .S1(net932),
    .X(net89));
 sky130_fd_sc_hd__mux4_2 c189 (.A0(net88),
    .A1(net87),
    .A2(net89),
    .A3(net83),
    .S0(net86),
    .S1(net618),
    .X(net90));
 sky130_fd_sc_hd__mux4_2 c190 (.A0(net89),
    .A1(net90),
    .A2(net822),
    .A3(net86),
    .S0(net83),
    .S1(net930),
    .X(net91));
 sky130_fd_sc_hd__mux4_2 c191 (.A0(net90),
    .A1(net91),
    .A2(net828),
    .A3(net89),
    .S0(net619),
    .S1(net932),
    .X(net92));
 sky130_fd_sc_hd__mux4_1 c192 (.A0(net85),
    .A1(net91),
    .A2(net89),
    .A3(net86),
    .S0(net92),
    .S1(net618),
    .X(net93));
 sky130_fd_sc_hd__mux4_1 c193 (.A0(net93),
    .A1(net81),
    .A2(net87),
    .A3(net86),
    .S0(net820),
    .S1(net90),
    .X(net94));
 sky130_fd_sc_hd__mux4_1 c194 (.A0(net92),
    .A1(net90),
    .A2(net94),
    .A3(net833),
    .S0(net825),
    .S1(net93),
    .X(net95));
 sky130_fd_sc_hd__mux4_1 c195 (.A0(net86),
    .A1(net91),
    .A2(net85),
    .A3(net94),
    .S0(net89),
    .S1(net930),
    .X(net96));
 sky130_fd_sc_hd__mux4_2 c196 (.A0(net94),
    .A1(net95),
    .A2(net93),
    .A3(net96),
    .S0(net91),
    .S1(net932),
    .X(net97));
 sky130_fd_sc_hd__mux4_2 c197 (.A0(net96),
    .A1(net97),
    .A2(net95),
    .A3(net93),
    .S0(net92),
    .S1(net619),
    .X(net98));
 sky130_fd_sc_hd__mux4_2 c198 (.A0(net98),
    .A1(net850),
    .A2(net845),
    .A3(net858),
    .S0(net847),
    .S1(net837),
    .X(net99));
 sky130_fd_sc_hd__a41o_2 c199 (.A1(net99),
    .A2(net847),
    .A3(net98),
    .A4(net853),
    .B1(net855),
    .X(net100));
 sky130_fd_sc_hd__sdfbbp_1 c200 (.CLK(clknet_4_2_0_clk),
    .D(net837),
    .RESET_B(net849),
    .SCD(net99),
    .SCE(net73),
    .SET_B(net100),
    .Q(net102),
    .Q_N(net101));
 sky130_fd_sc_hd__mux4_2 c201 (.A0(net100),
    .A1(net99),
    .A2(net101),
    .A3(net860),
    .S0(net854),
    .S1(net930),
    .X(net103));
 sky130_fd_sc_hd__mux4_2 c202 (.A0(net851),
    .A1(net99),
    .A2(net814),
    .A3(net103),
    .S0(net101),
    .S1(net100),
    .X(net104));
 sky130_fd_sc_hd__mux4_2 c203 (.A0(net103),
    .A1(net848),
    .A2(net99),
    .A3(net102),
    .S0(net104),
    .S1(net930),
    .X(net105));
 sky130_fd_sc_hd__mux4_2 c204 (.A0(net103),
    .A1(net832),
    .A2(net105),
    .A3(net104),
    .S0(net935),
    .S1(net99),
    .X(net106));
 sky130_fd_sc_hd__mux4_1 c205 (.A0(net106),
    .A1(net102),
    .A2(net104),
    .A3(net105),
    .S0(net103),
    .S1(net99),
    .X(net107));
 sky130_fd_sc_hd__mux4_1 c206 (.A0(net99),
    .A1(net103),
    .A2(net102),
    .A3(net105),
    .S0(net104),
    .S1(clknet_1_0__leaf_net711),
    .X(net108));
 sky130_fd_sc_hd__mux4_1 c207 (.A0(net105),
    .A1(net103),
    .A2(net860),
    .A3(clknet_1_0__leaf_net108),
    .S0(net106),
    .S1(clknet_1_0__leaf_net711),
    .X(net109));
 sky130_fd_sc_hd__mux4_1 c208 (.A0(net100),
    .A1(net106),
    .A2(clknet_1_0__leaf_net108),
    .A3(net105),
    .S0(clknet_1_0__leaf_net711),
    .S1(net728),
    .X(net110));
 sky130_fd_sc_hd__mux4_1 c209 (.A0(clknet_1_0__leaf_net108),
    .A1(net105),
    .A2(net640),
    .A3(clknet_1_0__leaf_net711),
    .S0(net930),
    .S1(net728),
    .X(net111));
 sky130_fd_sc_hd__mux4_1 c210 (.A0(net102),
    .A1(net856),
    .A2(clknet_1_1__leaf_net108),
    .A3(net645),
    .S0(net930),
    .S1(net728),
    .X(net112));
 sky130_fd_sc_hd__mux4_1 c211 (.A0(net105),
    .A1(clknet_1_1__leaf_net108),
    .A2(net106),
    .A3(net639),
    .S0(clknet_1_0__leaf_net711),
    .S1(net728),
    .X(net113));
 sky130_fd_sc_hd__a41o_1 c212 (.A1(clknet_1_1__leaf_net108),
    .A2(net106),
    .A3(net640),
    .A4(net645),
    .B1(clknet_1_0__leaf_net711),
    .X(net114));
 sky130_fd_sc_hd__mux4_1 c213 (.A0(clknet_1_1__leaf_net108),
    .A1(net102),
    .A2(net639),
    .A3(clknet_1_0__leaf_net676),
    .S0(net682),
    .S1(net728),
    .X(net115));
 sky130_fd_sc_hd__mux4_1 c214 (.A0(net100),
    .A1(net99),
    .A2(clknet_1_0__leaf_net676),
    .A3(net682),
    .S0(net728),
    .S1(clknet_1_0__leaf_net889),
    .X(net116));
 sky130_fd_sc_hd__a41o_1 c215 (.A1(net105),
    .A2(net640),
    .A3(clknet_1_0__leaf_net676),
    .A4(net682),
    .B1(clknet_1_0__leaf_net889),
    .X(net117));
 sky130_fd_sc_hd__mux4_1 c216 (.A0(net104),
    .A1(net106),
    .A2(clknet_1_0__leaf_net117),
    .A3(clknet_1_0__leaf_net116),
    .S0(net100),
    .S1(net682),
    .X(net118));
 sky130_fd_sc_hd__mux4_1 c217 (.A0(clknet_1_0__leaf_net116),
    .A1(clknet_1_0__leaf_net117),
    .A2(net855),
    .A3(net639),
    .S0(clknet_1_0__leaf_net676),
    .S1(clknet_1_0__leaf_net729),
    .X(net119));
 sky130_fd_sc_hd__mux4_1 c218 (.A0(net858),
    .A1(clknet_1_1__leaf_net116),
    .A2(clknet_1_1__leaf_net117),
    .S0(clknet_1_0__leaf_net676),
    .S1(net682),
    .X(net120));
 sky130_fd_sc_hd__a41o_1 c219 (.A1(clknet_1_1__leaf_net117),
    .A2(clknet_1_1__leaf_net116),
    .A3(net645),
    .A4(clknet_1_0__leaf_net889),
    .B1(clknet_1_0__leaf_net729),
    .X(net121));
 sky130_fd_sc_hd__a41o_1 c220 (.A1(net840),
    .A2(net935),
    .A3(net637),
    .A4(net645),
    .B1(clknet_1_1__leaf_net889),
    .X(net122));
 sky130_fd_sc_hd__a41o_1 c221 (.A1(clknet_1_1__leaf_net122),
    .A2(net102),
    .A3(net832),
    .A4(net0),
    .B1(clknet_1_1__leaf_net889),
    .X(net123));
 sky130_fd_sc_hd__a41o_1 c222 (.A1(clknet_1_0__leaf_net123),
    .A2(net818),
    .A3(net9),
    .A4(clknet_1_0__leaf_net122),
    .B1(clknet_1_1__leaf_net889),
    .X(net124));
 sky130_fd_sc_hd__a41o_1 c223 (.A1(clknet_1_0__leaf_net124),
    .A2(clknet_1_0__leaf_net123),
    .A3(clknet_1_1__leaf_net122),
    .A4(net637),
    .B1(clknet_1_1__leaf_net889),
    .X(net125));
 sky130_fd_sc_hd__a41o_1 c224 (.A1(clknet_1_1__leaf_net122),
    .A2(clknet_1_0__leaf_net124),
    .A3(clknet_1_0__leaf_net125),
    .A4(clknet_1_0__leaf_net123),
    .B1(clknet_1_1__leaf_net729),
    .X(net126));
 sky130_fd_sc_hd__mux4_1 c225 (.A0(clknet_1_0__leaf_net126),
    .A1(clknet_1_0__leaf_net125),
    .A2(clknet_1_0__leaf_net124),
    .A3(clknet_1_0__leaf_net123),
    .S0(clknet_1_0__leaf_net122),
    .S1(clknet_1_1__leaf_net889),
    .X(net127));
 sky130_fd_sc_hd__mux4_1 c226 (.A0(clknet_1_1__leaf_net122),
    .A1(clknet_1_0__leaf_net123),
    .A2(clknet_1_0__leaf_net124),
    .A3(clknet_1_0__leaf_net125),
    .S0(clknet_1_0__leaf_net127),
    .S1(net645),
    .X(net128));
 sky130_fd_sc_hd__mux4_1 c227 (.A0(clknet_1_0__leaf_net128),
    .A1(clknet_1_0__leaf_net127),
    .A2(clknet_1_0__leaf_net124),
    .A3(clknet_1_0__leaf_net125),
    .S0(net935),
    .S1(clknet_1_0__leaf_net123),
    .X(net129));
 sky130_fd_sc_hd__mux4_1 c228 (.A0(clknet_1_0__leaf_net123),
    .A1(clknet_1_0__leaf_net126),
    .A2(clknet_1_0__leaf_net124),
    .A3(clknet_1_0__leaf_net125),
    .S0(clknet_1_0__leaf_net128),
    .S1(clknet_1_0__leaf_net122),
    .X(net890));
 sky130_fd_sc_hd__mux4_1 c229 (.A0(clknet_1_0__leaf_net129),
    .A1(clknet_1_0__leaf_net128),
    .A2(clknet_1_1__leaf_net125),
    .A3(clknet_1_0__leaf_net890),
    .S0(clknet_1_1__leaf_net123),
    .S1(clknet_1_1__leaf_net124),
    .X(net130));
 sky130_fd_sc_hd__mux4_1 c230 (.A0(clknet_1_1__leaf_net123),
    .A1(clknet_1_0__leaf_net129),
    .A2(clknet_1_0__leaf_net128),
    .A3(clknet_1_1__leaf_net125),
    .S0(clknet_1_0__leaf_net130),
    .S1(clknet_1_1__leaf_net124),
    .X(net131));
 sky130_fd_sc_hd__mux4_1 c231 (.A0(clknet_1_1__leaf_net124),
    .A1(clknet_1_0__leaf_net130),
    .A2(clknet_1_0__leaf_net131),
    .A3(clknet_1_1__leaf_net129),
    .S0(clknet_1_1__leaf_net123),
    .S1(clknet_1_0__leaf_net890),
    .X(net132));
 sky130_fd_sc_hd__mux4_1 c232 (.A0(clknet_1_1__leaf_net130),
    .A1(clknet_1_0__leaf_net132),
    .A2(clknet_1_1__leaf_net127),
    .A3(clknet_1_0__leaf_net131),
    .S0(clknet_1_1__leaf_net123),
    .S1(clknet_1_1__leaf_net124),
    .X(net133));
 sky130_fd_sc_hd__mux4_1 c233 (.A0(clknet_1_0__leaf_net133),
    .A1(clknet_1_1__leaf_net131),
    .A2(clknet_1_1__leaf_net130),
    .A3(clknet_1_1__leaf_net123),
    .S0(clknet_1_1__leaf_net128),
    .S1(clknet_1_0__leaf_net132),
    .X(net134));
 sky130_fd_sc_hd__mux4_1 c234 (.A0(clknet_1_0__leaf_net132),
    .A1(clknet_1_1__leaf_net133),
    .A2(clknet_1_1__leaf_net127),
    .A3(clknet_1_1__leaf_net134),
    .S0(clknet_1_1__leaf_net130),
    .S1(clknet_1_1__leaf_net123),
    .X(net135));
 sky130_fd_sc_hd__mux4_1 c235 (.A0(clknet_1_1__leaf_net131),
    .A1(clknet_1_1__leaf_net130),
    .A2(clknet_1_1__leaf_net134),
    .A3(clknet_1_1__leaf_net124),
    .S0(clknet_1_0__leaf_net133),
    .S1(clknet_1_1__leaf_net128),
    .X(net136));
 sky130_fd_sc_hd__mux4_1 c236 (.A0(clknet_1_0__leaf_net127),
    .A1(clknet_1_0__leaf_net135),
    .A2(clknet_1_0__leaf_net136),
    .A3(clknet_1_0__leaf_net130),
    .S0(clknet_1_1__leaf_net126),
    .S1(clknet_1_0__leaf_net134),
    .X(net137));
 sky130_fd_sc_hd__mux4_1 c237 (.A0(clknet_1_0__leaf_net125),
    .A1(clknet_1_0__leaf_net135),
    .A2(clknet_1_0__leaf_net132),
    .A3(clknet_1_0__leaf_net137),
    .S0(clknet_1_1__leaf_net126),
    .S1(clknet_1_0__leaf_net123),
    .X(net138));
 sky130_fd_sc_hd__mux4_1 c238 (.A0(clknet_1_0__leaf_net138),
    .A1(clknet_1_1__leaf_net135),
    .A2(clknet_1_0__leaf_net124),
    .A3(clknet_1_0__leaf_net136),
    .S0(clknet_1_0__leaf_net134),
    .S1(clknet_1_1__leaf_net729),
    .X(net139));
 sky130_fd_sc_hd__mux4_1 c239 (.A0(clknet_1_0__leaf_net139),
    .A1(clknet_1_0__leaf_net134),
    .A2(clknet_1_0__leaf_net137),
    .A3(clknet_1_1__leaf_net136),
    .S0(clknet_1_0__leaf_net138),
    .S1(clknet_1_0__leaf_net132),
    .X(net140));
 sky130_fd_sc_hd__mux4_1 c240 (.A0(clknet_1_0__leaf_net128),
    .A1(clknet_1_1__leaf_net136),
    .A2(clknet_1_1__leaf_net138),
    .A3(clknet_1_1__leaf_net139),
    .S0(clknet_1_0__leaf_net130),
    .S1(net681),
    .X(net141));
 sky130_fd_sc_hd__a41o_1 c241 (.A1(clknet_1_1__leaf_net137),
    .A2(clknet_1_1__leaf_net125),
    .A3(clknet_1_1__leaf_net138),
    .A4(clknet_1_1__leaf_net134),
    .B1(net681),
    .X(net142));
 sky130_fd_sc_hd__a41o_1 c256 (.A1(net893),
    .A2(net913),
    .A3(clknet_1_1__leaf_net132),
    .A4(clknet_1_1__leaf_net890),
    .B1(net681),
    .X(net895));
 sky130_fd_sc_hd__sdfbbn_1 c257 (.CLK_N(clknet_4_10_0_clk),
    .D(clknet_1_1__leaf_net142),
    .RESET_B(clknet_1_1__leaf_net895),
    .SCD(net913),
    .SCE(clknet_1_1__leaf_net132),
    .SET_B(clknet_1_1__leaf_net890),
    .Q(net899),
    .Q_N(net143));
 sky130_fd_sc_hd__a41o_1 c258 (.A1(clknet_1_0__leaf_net895),
    .A2(net899),
    .A3(clknet_1_1__leaf_net132),
    .A4(net913),
    .B1(net692),
    .X(net898));
 sky130_fd_sc_hd__a41o_1 c259 (.A1(clknet_1_0__leaf_net898),
    .A2(net143),
    .A3(clknet_1_0__leaf_net895),
    .A4(net913),
    .B1(clknet_1_1__leaf_net132),
    .X(net894));
 sky130_fd_sc_hd__a41o_1 c260 (.A1(net899),
    .A2(clknet_1_0__leaf_net894),
    .A3(clknet_1_0__leaf_net898),
    .A4(clknet_1_0__leaf_net895),
    .B1(net913),
    .X(net901));
 sky130_fd_sc_hd__mux4_1 c261 (.A0(clknet_1_0__leaf_net898),
    .A1(clknet_1_0__leaf_net901),
    .A2(clknet_1_0__leaf_net894),
    .A3(net143),
    .S0(clknet_1_1__leaf_net895),
    .S1(net20),
    .X(net144));
 sky130_fd_sc_hd__mux4_1 c262 (.A0(net20),
    .A1(clknet_1_0__leaf_net901),
    .A2(net143),
    .A3(clknet_1_1__leaf_net898),
    .S0(clknet_1_0__leaf_net894),
    .S1(net900),
    .X(net145));
 sky130_fd_sc_hd__mux4_1 c263 (.A0(clknet_1_1__leaf_net901),
    .A1(clknet_1_1__leaf_net898),
    .A2(clknet_1_0__leaf_net894),
    .S0(net681),
    .S1(clknet_1_0__leaf_net891),
    .X(net146));
 sky130_fd_sc_hd__a41o_1 c264 (.A1(net786),
    .A2(net52),
    .A3(net254),
    .A4(net50),
    .B1(net43),
    .X(net147));
 sky130_fd_sc_hd__a41o_1 c265 (.A1(net911),
    .A2(net782),
    .A3(net43),
    .A4(net819),
    .B1(net841),
    .X(net148));
 sky130_fd_sc_hd__a31o_2 c266 (.A1(net909),
    .A2(net911),
    .A3(net50),
    .B1(net43),
    .X(net149));
 sky130_fd_sc_hd__a31o_1 c267 (.A1(net911),
    .A2(net909),
    .A3(net149),
    .B1(net43),
    .X(net150));
 sky130_fd_sc_hd__sdfbbn_1 c268 (.CLK_N(clknet_4_1_0_clk),
    .D(net909),
    .RESET_B(net911),
    .SCD(net149),
    .SCE(net43),
    .SET_B(net933),
    .Q(net152),
    .Q_N(net151));
 sky130_fd_sc_hd__a41o_1 c269 (.A1(net909),
    .A2(net911),
    .A3(net152),
    .A4(net149),
    .B1(net933),
    .X(net153));
 sky130_fd_sc_hd__mux4_1 c270 (.A0(net911),
    .A1(net152),
    .A2(net909),
    .A3(net149),
    .S1(net933),
    .X(net154));
 sky130_fd_sc_hd__a41o_1 c271 (.A1(net152),
    .A2(net911),
    .A3(net909),
    .A4(net149),
    .B1(net674),
    .X(net155));
 sky130_fd_sc_hd__mux4_1 c272 (.A0(net151),
    .A1(net147),
    .A2(net148),
    .A3(net149),
    .S0(net674),
    .S1(clknet_1_1__leaf_net709),
    .X(net156));
 sky130_fd_sc_hd__mux4_1 c273 (.A0(net149),
    .A1(net152),
    .A2(net147),
    .A3(net674),
    .S0(clknet_1_1__leaf_net709),
    .S1(net933),
    .X(net157));
 sky130_fd_sc_hd__mux4_1 c274 (.A0(net149),
    .A1(net911),
    .A2(net909),
    .A3(net151),
    .S0(net669),
    .S1(net718),
    .X(net158));
 sky130_fd_sc_hd__mux4_1 c275 (.A0(net911),
    .A1(net151),
    .A2(net674),
    .A3(clknet_1_1__leaf_net709),
    .S0(net718),
    .S1(net730),
    .X(net159));
 sky130_fd_sc_hd__mux4_1 c276 (.A0(clknet_1_0__leaf_net159),
    .A1(net911),
    .A2(net151),
    .A3(clknet_1_1__leaf_net709),
    .S0(net718),
    .S1(net731),
    .X(net160));
 sky130_fd_sc_hd__mux4_1 c277 (.A0(clknet_1_0__leaf_net160),
    .A1(clknet_1_1__leaf_net159),
    .A2(net152),
    .A3(net909),
    .S0(clknet_1_1__leaf_net709),
    .S1(net730),
    .X(net161));
 sky130_fd_sc_hd__mux4_1 c278 (.A0(clknet_1_1__leaf_net160),
    .A1(net148),
    .A2(net647),
    .A3(net674),
    .S0(net718),
    .S1(net731),
    .X(net162));
 sky130_fd_sc_hd__mux4_1 c279 (.A0(net152),
    .A1(net149),
    .A2(clknet_1_1__leaf_net159),
    .A3(net147),
    .S0(net647),
    .S1(clknet_1_1__leaf_net710),
    .X(net163));
 sky130_fd_sc_hd__mux4_1 c280 (.A0(clknet_1_0__leaf_net159),
    .A1(net909),
    .A2(net151),
    .A3(net669),
    .S0(net683),
    .S1(clknet_1_1__leaf_net710),
    .X(net164));
 sky130_fd_sc_hd__mux4_1 c281 (.A0(clknet_1_0__leaf_net164),
    .A1(net909),
    .A2(clknet_1_0__leaf_net159),
    .A3(net683),
    .S0(clknet_1_1__leaf_net710),
    .S1(net718),
    .X(net165));
 sky130_fd_sc_hd__mux4_1 c282 (.A0(net84),
    .A1(net151),
    .A2(clknet_1_0__leaf_net159),
    .A3(net674),
    .S0(clknet_1_0__leaf_net710),
    .S1(net730),
    .X(net166));
 sky130_fd_sc_hd__mux4_1 c283 (.A0(clknet_1_1__leaf_net164),
    .A1(clknet_1_1__leaf_net159),
    .A2(net647),
    .A3(net683),
    .S0(clknet_1_1__leaf_net710),
    .S1(net731),
    .X(net167));
 sky130_fd_sc_hd__a41o_1 c284 (.A1(clknet_1_0__leaf_net166),
    .A2(net149),
    .A3(net669),
    .A4(net683),
    .B1(net694),
    .X(net168));
 sky130_fd_sc_hd__mux4_1 c285 (.A0(clknet_1_1__leaf_net159),
    .A1(clknet_1_0__leaf_net166),
    .A2(net648),
    .A3(net669),
    .S0(net933),
    .S1(net718),
    .X(net169));
 sky130_fd_sc_hd__sdfbbp_1 c286 (.CLK(clknet_4_1_0_clk),
    .D(net71),
    .RESET_B(net795),
    .SCD(net908),
    .SCE(net794),
    .SET_B(net943),
    .Q(net171),
    .Q_N(net170));
 sky130_fd_sc_hd__sdfbbn_2 c287 (.CLK_N(clknet_4_1_0_clk),
    .D(net170),
    .RESET_B(net908),
    .SCD(net803),
    .SCE(net694),
    .SET_B(net706),
    .Q(net173),
    .Q_N(net172));
 sky130_fd_sc_hd__sdfbbn_2 c288 (.CLK_N(clknet_4_0_0_clk),
    .D(net173),
    .RESET_B(net171),
    .SCD(net805),
    .SCE(net908),
    .SET_B(net643),
    .Q(net175),
    .Q_N(net174));
 sky130_fd_sc_hd__a41o_1 c289 (.A1(net175),
    .A2(net170),
    .A3(net172),
    .A4(net908),
    .B1(net642),
    .X(net176));
 sky130_fd_sc_hd__a41o_1 c290 (.A1(net175),
    .A2(net170),
    .A3(net172),
    .A4(clknet_1_0__leaf_net709),
    .B1(net725),
    .X(net177));
 sky130_fd_sc_hd__mux4_1 c291 (.A0(net793),
    .A1(clknet_1_1__leaf_net177),
    .A2(net173),
    .A3(net175),
    .S0(net170),
    .S1(clknet_1_0__leaf_net709),
    .X(net178));
 sky130_fd_sc_hd__mux4_1 c292 (.A0(net171),
    .A1(clknet_1_0__leaf_net177),
    .A2(net175),
    .A3(net172),
    .S0(clknet_1_0__leaf_net178),
    .S1(clknet_1_0__leaf_net709),
    .X(net179));
 sky130_fd_sc_hd__mux4_1 c293 (.A0(clknet_1_0__leaf_net179),
    .A1(clknet_1_0__leaf_net177),
    .A2(net174),
    .A3(net172),
    .S0(clknet_1_0__leaf_net709),
    .S1(net724),
    .X(net180));
 sky130_fd_sc_hd__mux4_1 c294 (.A0(net173),
    .A1(clknet_1_1__leaf_net178),
    .A2(net170),
    .A3(clknet_1_1__leaf_net179),
    .S0(net642),
    .S1(clknet_1_0__leaf_net709),
    .X(net181));
 sky130_fd_sc_hd__mux4_1 c295 (.A0(clknet_1_0__leaf_net178),
    .A1(net171),
    .A2(clknet_1_0__leaf_net181),
    .A3(clknet_1_0__leaf_net179),
    .S0(net175),
    .S1(clknet_1_0__leaf_net180),
    .X(net182));
 sky130_fd_sc_hd__mux4_1 c296 (.A0(net43),
    .A1(net173),
    .A2(clknet_1_0__leaf_net181),
    .A3(clknet_1_0__leaf_net180),
    .S0(clknet_1_0__leaf_net179),
    .S1(net174),
    .X(net183));
 sky130_fd_sc_hd__mux4_1 c297 (.A0(clknet_1_0__leaf_net181),
    .A1(clknet_1_0__leaf_net182),
    .A2(clknet_1_0__leaf_net179),
    .A3(net173),
    .S0(clknet_1_0__leaf_net183),
    .S1(clknet_1_1__leaf_net180),
    .X(net184));
 sky130_fd_sc_hd__mux4_1 c298 (.A0(clknet_1_1__leaf_net182),
    .A1(clknet_1_1__leaf_net184),
    .A2(clknet_1_0__leaf_net181),
    .A3(clknet_1_0__leaf_net179),
    .S0(net172),
    .S1(clknet_1_1__leaf_net180),
    .X(net185));
 sky130_fd_sc_hd__mux4_1 c299 (.A0(clknet_1_1__leaf_net180),
    .A1(clknet_1_0__leaf_net185),
    .A2(clknet_1_0__leaf_net181),
    .A3(clknet_1_0__leaf_net179),
    .S0(net172),
    .S1(clknet_1_0__leaf_net184),
    .X(net186));
 sky130_fd_sc_hd__mux4_1 c300 (.A0(clknet_1_0__leaf_net186),
    .A1(clknet_1_0__leaf_net183),
    .A2(clknet_1_0__leaf_net185),
    .A3(net173),
    .S0(clknet_1_1__leaf_net184),
    .S1(clknet_1_1__leaf_net181),
    .X(net187));
 sky130_fd_sc_hd__mux4_1 c301 (.A0(clknet_1_1__leaf_net179),
    .A1(clknet_1_1__leaf_net181),
    .A2(clknet_1_0__leaf_net187),
    .A3(clknet_1_0__leaf_net186),
    .S0(clknet_1_0__leaf_net185),
    .S1(clknet_1_0__leaf_net184),
    .X(net188));
 sky130_fd_sc_hd__mux4_1 c302 (.A0(clknet_1_0__leaf_net188),
    .A1(clknet_1_0__leaf_net186),
    .A2(clknet_1_1__leaf_net179),
    .A3(clknet_1_0__leaf_net185),
    .S0(net173),
    .S1(clknet_1_1__leaf_net181),
    .X(net189));
 sky130_fd_sc_hd__mux4_1 c303 (.A0(clknet_1_0__leaf_net166),
    .A1(clknet_1_1__leaf_net187),
    .A2(clknet_1_1__leaf_net185),
    .A3(net175),
    .S0(clknet_1_0__leaf_net189),
    .S1(clknet_1_1__leaf_net181),
    .X(net190));
 sky130_fd_sc_hd__mux4_1 c304 (.A0(clknet_1_1__leaf_net183),
    .A1(clknet_1_1__leaf_net188),
    .A2(clknet_1_1__leaf_net185),
    .A3(clknet_1_1__leaf_net179),
    .S0(clknet_1_0__leaf_net189),
    .S1(net680),
    .X(net191));
 sky130_fd_sc_hd__mux4_1 c305 (.A0(net73),
    .A1(clknet_1_1__leaf_net191),
    .A2(clknet_1_1__leaf_net186),
    .A3(net171),
    .S0(clknet_1_1__leaf_net185),
    .S1(net680),
    .X(net192));
 sky130_fd_sc_hd__a41o_1 c306 (.A1(clknet_1_1__leaf_net185),
    .A2(net171),
    .A3(clknet_1_0__leaf_net191),
    .A4(clknet_1_1__leaf_net186),
    .B1(net680),
    .X(net193));
 sky130_fd_sc_hd__mux4_1 c307 (.A0(clknet_1_1__leaf_net189),
    .A1(clknet_1_0__leaf_net191),
    .A2(clknet_1_1__leaf_net193),
    .A3(clknet_1_1__leaf_net186),
    .S0(clknet_1_1__leaf_net185),
    .S1(net680),
    .X(net194));
 sky130_fd_sc_hd__mux4_1 c308 (.A0(net97),
    .A1(clknet_1_0__leaf_net194),
    .A2(clknet_1_0__leaf_net193),
    .A3(net174),
    .S0(net73),
    .S1(net931),
    .X(net195));
 sky130_fd_sc_hd__a41o_1 c309 (.A1(net97),
    .A2(net98),
    .A3(net174),
    .A4(net931),
    .B1(net733),
    .X(net196));
 sky130_fd_sc_hd__mux4_1 c310 (.A0(clknet_1_0__leaf_net193),
    .A1(net902),
    .A2(net813),
    .A3(net97),
    .S0(net931),
    .S1(net733),
    .X(net197));
 sky130_fd_sc_hd__mux4_1 c311 (.A0(net81),
    .A1(net826),
    .A2(net902),
    .A3(clknet_1_0__leaf_net197),
    .S0(net97),
    .S1(net732),
    .X(net198));
 sky130_fd_sc_hd__mux4_1 c312 (.A0(net902),
    .A1(clknet_1_0__leaf_net197),
    .A2(clknet_1_0__leaf_net193),
    .A3(net696),
    .S0(net931),
    .S1(net733),
    .X(net199));
 sky130_fd_sc_hd__mux4_1 c313 (.A0(clknet_1_0__leaf_net184),
    .A1(clknet_1_0__leaf_net197),
    .A2(net902),
    .A3(net696),
    .S0(net732),
    .S1(net734),
    .X(net200));
 sky130_fd_sc_hd__mux4_1 c314 (.A0(net902),
    .A1(clknet_1_0__leaf_net197),
    .A2(net696),
    .A3(net732),
    .S0(net734),
    .S1(net929),
    .X(net201));
 sky130_fd_sc_hd__mux4_1 c315 (.A0(net67),
    .A1(net97),
    .A2(net902),
    .A3(clknet_1_1__leaf_net197),
    .S0(net701),
    .S1(net929),
    .X(net202));
 sky130_fd_sc_hd__mux4_1 c316 (.A0(net196),
    .A1(clknet_1_0__leaf_net197),
    .A2(net701),
    .A3(net732),
    .S0(net735),
    .S1(net929),
    .X(net203));
 sky130_fd_sc_hd__mux4_2 c317 (.A0(net902),
    .A1(net649),
    .A2(net670),
    .A3(net701),
    .S0(net735),
    .S1(net929),
    .X(net204));
 sky130_fd_sc_hd__mux4_1 c318 (.A0(net204),
    .A1(net902),
    .A2(net649),
    .A3(net701),
    .S0(net734),
    .S1(net929),
    .X(net205));
 sky130_fd_sc_hd__mux4_1 c319 (.A0(net205),
    .A1(net196),
    .A2(clknet_1_0__leaf_net197),
    .A3(net696),
    .S0(net734),
    .S1(net929),
    .X(net206));
 sky130_fd_sc_hd__mux4_1 c320 (.A0(net204),
    .A1(net205),
    .A2(clknet_1_1__leaf_net710),
    .A3(net733),
    .S0(net929),
    .S1(net928),
    .X(net207));
 sky130_fd_sc_hd__mux4_1 c321 (.A0(net175),
    .A1(clknet_1_0__leaf_net207),
    .A2(net97),
    .A3(net735),
    .S0(net929),
    .S1(net928),
    .X(net208));
 sky130_fd_sc_hd__mux4_1 c322 (.A0(clknet_1_0__leaf_net208),
    .A1(clknet_1_0__leaf_net207),
    .A2(net650),
    .A3(net670),
    .S0(net929),
    .S1(net928),
    .X(net209));
 sky130_fd_sc_hd__mux4_1 c323 (.A0(net205),
    .A1(clknet_1_0__leaf_net208),
    .A2(clknet_1_0__leaf_net209),
    .A3(clknet_1_1__leaf_net197),
    .S0(net670),
    .S1(net931),
    .X(net210));
 sky130_fd_sc_hd__mux4_1 c324 (.A0(clknet_1_1__leaf_net207),
    .A1(clknet_1_1__leaf_net209),
    .A2(clknet_1_1__leaf_net208),
    .A3(net204),
    .S0(net902),
    .S1(net706),
    .X(net211));
 sky130_fd_sc_hd__mux4_1 c325 (.A0(clknet_1_1__leaf_net208),
    .A1(net902),
    .A2(net683),
    .A3(net701),
    .S0(net706),
    .S1(net929),
    .X(net212));
 sky130_fd_sc_hd__mux4_1 c326 (.A0(clknet_1_1__leaf_net212),
    .A1(clknet_1_0__leaf_net209),
    .A2(net683),
    .A3(net706),
    .S0(net735),
    .S1(net736),
    .X(net213));
 sky130_fd_sc_hd__mux4_1 c327 (.A0(clknet_1_1__leaf_net212),
    .A1(net670),
    .A2(net683),
    .A3(net686),
    .S0(net706),
    .S1(net928),
    .X(net214));
 sky130_fd_sc_hd__mux4_1 c328 (.A0(clknet_1_1__leaf_net197),
    .A1(clknet_1_0__leaf_net212),
    .A2(net683),
    .A3(net686),
    .S0(net706),
    .S1(net735),
    .X(net215));
 sky130_fd_sc_hd__a41o_1 c329 (.A1(net204),
    .A2(clknet_1_0__leaf_net212),
    .A3(net686),
    .A4(net696),
    .B1(net733),
    .X(net216));
 sky130_fd_sc_hd__mux4_1 c330 (.A0(net816),
    .A1(net935),
    .A2(net838),
    .A3(clknet_1_0__leaf_net889),
    .S0(clknet_1_1__leaf_net729),
    .S1(net928),
    .X(net217));
 sky130_fd_sc_hd__a41o_1 c331 (.A1(net839),
    .A2(clknet_1_1__leaf_net217),
    .A3(net843),
    .A4(clknet_1_1__leaf_net889),
    .B1(net928),
    .X(net218));
 sky130_fd_sc_hd__a41o_1 c332 (.A1(clknet_1_0__leaf_net218),
    .A2(clknet_1_0__leaf_net217),
    .A3(net175),
    .A4(net645),
    .B1(clknet_1_0__leaf_net729),
    .X(net219));
 sky130_fd_sc_hd__a41o_1 c333 (.A1(clknet_1_1__leaf_net217),
    .A2(clknet_1_0__leaf_net219),
    .A3(clknet_1_1__leaf_net218),
    .A4(net935),
    .B1(clknet_1_0__leaf_net889),
    .X(net220));
 sky130_fd_sc_hd__mux4_1 c334 (.A0(clknet_1_0__leaf_net219),
    .A1(clknet_1_0__leaf_net220),
    .A2(net102),
    .A3(clknet_1_0__leaf_net217),
    .S0(clknet_1_0__leaf_net218),
    .S1(net928),
    .X(net221));
 sky130_fd_sc_hd__mux4_1 c335 (.A0(clknet_1_0__leaf_net221),
    .A1(clknet_1_0__leaf_net219),
    .A2(clknet_1_0__leaf_net220),
    .A3(clknet_1_0__leaf_net217),
    .S0(clknet_1_0__leaf_net218),
    .S1(net928),
    .X(net222));
 sky130_fd_sc_hd__mux4_1 c336 (.A0(clknet_1_0__leaf_net221),
    .A1(clknet_1_0__leaf_net222),
    .A2(clknet_1_0__leaf_net219),
    .A3(clknet_1_0__leaf_net220),
    .S0(clknet_1_0__leaf_net217),
    .S1(clknet_1_0__leaf_net218),
    .X(net223));
 sky130_fd_sc_hd__mux4_1 c337 (.A0(clknet_1_0__leaf_net217),
    .A1(clknet_1_0__leaf_net219),
    .A2(clknet_1_0__leaf_net222),
    .A3(clknet_1_1__leaf_net221),
    .S0(clknet_1_0__leaf_net220),
    .S1(clknet_1_0__leaf_net223),
    .X(net224));
 sky130_fd_sc_hd__mux4_1 c338 (.A0(net102),
    .A1(clknet_1_0__leaf_net224),
    .A2(clknet_1_1__leaf_net223),
    .A3(clknet_1_1__leaf_net222),
    .S0(clknet_1_0__leaf_net219),
    .S1(clknet_1_1__leaf_net220),
    .X(net225));
 sky130_fd_sc_hd__mux4_1 c339 (.A0(clknet_1_0__leaf_net222),
    .A1(clknet_1_0__leaf_net217),
    .A2(clknet_1_0__leaf_net223),
    .A3(clknet_1_1__leaf_net220),
    .S0(clknet_1_0__leaf_net219),
    .S1(clknet_1_1__leaf_net221),
    .X(net226));
 sky130_fd_sc_hd__mux4_1 c340 (.A0(clknet_1_0__leaf_net226),
    .A1(clknet_1_0__leaf_net223),
    .A2(clknet_1_0__leaf_net225),
    .A3(clknet_1_0__leaf_net219),
    .S0(clknet_1_1__leaf_net221),
    .S1(clknet_1_1__leaf_net220),
    .X(net227));
 sky130_fd_sc_hd__mux4_1 c341 (.A0(clknet_1_1__leaf_net218),
    .A1(clknet_1_0__leaf_net227),
    .A2(clknet_1_0__leaf_net226),
    .A3(clknet_1_1__leaf_net222),
    .S0(clknet_1_0__leaf_net220),
    .S1(clknet_1_0__leaf_net225),
    .X(net228));
 sky130_fd_sc_hd__mux4_1 c342 (.A0(clknet_1_1__leaf_net223),
    .A1(clknet_1_0__leaf_net226),
    .A2(clknet_1_0__leaf_net228),
    .A3(clknet_1_0__leaf_net222),
    .S0(clknet_1_1__leaf_net220),
    .S1(clknet_1_0__leaf_net227),
    .X(net229));
 sky130_fd_sc_hd__mux4_1 c343 (.A0(clknet_1_1__leaf_net224),
    .A1(clknet_1_0__leaf_net229),
    .A2(clknet_1_1__leaf_net226),
    .A3(clknet_1_0__leaf_net228),
    .S0(clknet_1_1__leaf_net220),
    .S1(clknet_1_1__leaf_net225),
    .X(net230));
 sky130_fd_sc_hd__mux4_1 c344 (.A0(clknet_1_1__leaf_net230),
    .A1(clknet_1_0__leaf_net226),
    .A2(clknet_1_1__leaf_net222),
    .A3(clknet_1_1__leaf_net228),
    .S0(clknet_1_1__leaf_net220),
    .S1(clknet_1_0__leaf_net227),
    .X(net231));
 sky130_fd_sc_hd__mux4_1 c345 (.A0(clknet_1_1__leaf_net229),
    .A1(clknet_1_1__leaf_net223),
    .A2(clknet_1_0__leaf_net228),
    .A3(clknet_1_1__leaf_net230),
    .S0(clknet_1_1__leaf_net231),
    .S1(clknet_1_1__leaf_net226),
    .X(net232));
 sky130_fd_sc_hd__mux4_1 c346 (.A0(clknet_1_0__leaf_net220),
    .A1(clknet_1_0__leaf_net230),
    .A2(clknet_1_1__leaf_net217),
    .A3(clknet_1_0__leaf_net232),
    .S0(clknet_1_0__leaf_net219),
    .S1(clknet_1_0__leaf_net228),
    .X(net233));
 sky130_fd_sc_hd__mux4_1 c347 (.A0(clknet_1_0__leaf_net231),
    .A1(clknet_1_0__leaf_net233),
    .A2(clknet_1_0__leaf_net232),
    .A3(clknet_1_0__leaf_net230),
    .S0(clknet_1_1__leaf_net222),
    .S1(net637),
    .X(net234));
 sky130_fd_sc_hd__mux4_1 c348 (.A0(clknet_1_0__leaf_net234),
    .A1(clknet_1_1__leaf_net228),
    .A2(clknet_1_1__leaf_net218),
    .A3(clknet_1_0__leaf_net231),
    .S0(clknet_1_0__leaf_net232),
    .S1(clknet_1_1__leaf_net226),
    .X(net235));
 sky130_fd_sc_hd__mux4_1 c349 (.A0(clknet_1_1__leaf_net225),
    .A1(clknet_1_0__leaf_net235),
    .A2(clknet_1_0__leaf_net233),
    .A3(clknet_1_0__leaf_net234),
    .S0(clknet_1_1__leaf_net226),
    .S1(clknet_1_1__leaf_net231),
    .X(net236));
 sky130_fd_sc_hd__mux4_1 c350 (.A0(clknet_1_1__leaf_net227),
    .A1(clknet_1_0__leaf_net236),
    .A2(clknet_1_1__leaf_net232),
    .A3(clknet_1_1__leaf_net234),
    .S0(clknet_1_1__leaf_net230),
    .S1(clknet_1_1__leaf_net228),
    .X(net237));
 sky130_fd_sc_hd__mux4_1 c351 (.A0(clknet_1_1__leaf_net232),
    .A1(net237),
    .A2(clknet_1_1__leaf_net227),
    .A3(clknet_1_1__leaf_net235),
    .S0(clknet_1_1__leaf_net236),
    .S1(clknet_1_1__leaf_net228),
    .X(net238));
 sky130_fd_sc_hd__sdfbbp_1 c352 (.CLK(clknet_4_8_0_clk),
    .D(clknet_1_0__leaf_net132),
    .RESET_B(clknet_1_0__leaf_net890),
    .SCD(clknet_1_0__leaf_net142),
    .SCE(clknet_1_1__leaf_net219),
    .SET_B(net681),
    .Q(net240),
    .Q_N(net239));
 sky130_fd_sc_hd__sdfbbn_1 c353 (.CLK_N(clknet_4_8_0_clk),
    .D(net240),
    .RESET_B(clknet_1_1__leaf_net132),
    .SCD(clknet_1_1__leaf_net219),
    .SCE(clknet_1_0__leaf_net142),
    .SET_B(clknet_1_1__leaf_net889),
    .Q(net242),
    .Q_N(net241));
 sky130_fd_sc_hd__a41o_1 c354 (.A1(clknet_1_1__leaf_net233),
    .A2(net240),
    .A3(net242),
    .A4(clknet_1_0__leaf_net132),
    .B1(clknet_1_1__leaf_net219),
    .X(net243));
 sky130_fd_sc_hd__a41o_1 c355 (.A1(net240),
    .A2(clknet_1_1__leaf_net219),
    .A3(net241),
    .A4(clknet_1_1__leaf_net243),
    .B1(clknet_1_0__leaf_net132),
    .X(net244));
 sky130_fd_sc_hd__mux4_1 c356 (.A0(clknet_1_1__leaf_net243),
    .A1(clknet_1_1__leaf_net244),
    .A2(net239),
    .A3(clknet_1_1__leaf_net219),
    .S0(net241),
    .S1(clknet_1_1__leaf_net238),
    .X(net245));
 sky130_fd_sc_hd__a41o_1 c357 (.A1(clknet_1_1__leaf_net244),
    .A2(clknet_1_1__leaf_net243),
    .A3(net239),
    .A4(net241),
    .B1(net671),
    .X(net246));
 sky130_fd_sc_hd__mux4_1 c358 (.A0(clknet_1_1__leaf_net219),
    .A1(clknet_1_0__leaf_net246),
    .A2(clknet_1_0__leaf_net244),
    .A3(net239),
    .S0(net241),
    .S1(net671),
    .X(net247));
 sky130_fd_sc_hd__mux4_1 c359 (.A0(clknet_1_0__leaf_net890),
    .A1(clknet_1_0__leaf_net244),
    .A2(clknet_1_1__leaf_net247),
    .A3(clknet_1_0__leaf_net246),
    .S0(net239),
    .S1(clknet_1_0__leaf_net243),
    .X(net248));
 sky130_fd_sc_hd__mux4_1 c360 (.A0(clknet_1_0__leaf_net246),
    .A1(clknet_1_1__leaf_net247),
    .A2(net242),
    .A3(net97),
    .S0(clknet_1_0__leaf_net244),
    .S1(net239),
    .X(net249));
 sky130_fd_sc_hd__mux4_1 c361 (.A0(net242),
    .A1(clknet_1_1__leaf_net246),
    .A2(clknet_1_0__leaf_net247),
    .A3(clknet_1_1__leaf_net244),
    .S0(net240),
    .S1(clknet_1_1__leaf_net248),
    .X(net250));
 sky130_fd_sc_hd__mux4_1 c362 (.A0(net240),
    .A1(clknet_1_1__leaf_net246),
    .A2(clknet_1_1__leaf_net247),
    .A3(clknet_1_1__leaf_net248),
    .S0(clknet_1_1__leaf_net249),
    .S1(net671),
    .X(net251));
 sky130_fd_sc_hd__mux4_1 c363 (.A0(clknet_1_1__leaf_net247),
    .A1(clknet_1_1__leaf_net249),
    .A2(clknet_1_0__leaf_net244),
    .A3(clknet_1_0__leaf_net654),
    .S0(net671),
    .S1(net927),
    .X(net252));
 sky130_fd_sc_hd__mux4_1 c364 (.A0(clknet_1_0__leaf_net248),
    .A1(clknet_1_0__leaf_net243),
    .A2(clknet_1_0__leaf_net249),
    .A3(net240),
    .S0(clknet_1_0__leaf_net654),
    .S1(clknet_1_1__leaf_net711),
    .X(net253));
 sky130_fd_sc_hd__mux4_1 c365 (.A0(clknet_1_0__leaf_net243),
    .A1(clknet_1_0__leaf_net248),
    .A3(clknet_1_1__leaf_net676),
    .S0(clknet_1_1__leaf_net711),
    .S1(net927),
    .X(net654));
 sky130_fd_sc_hd__mux4_1 c366 (.A0(clknet_1_0__leaf_net249),
    .A1(clknet_1_0__leaf_net247),
    .A2(clknet_1_0__leaf_net132),
    .A3(net653),
    .S0(clknet_1_1__leaf_net676),
    .S1(clknet_1_1__leaf_net711),
    .X(net255));
 sky130_fd_sc_hd__mux4_1 c367 (.A0(clknet_1_0__leaf_net247),
    .A1(clknet_1_0__leaf_net132),
    .A2(net650),
    .A3(net653),
    .S0(clknet_1_1__leaf_net676),
    .S1(clknet_1_1__leaf_net711),
    .X(net256));
 sky130_fd_sc_hd__mux4_1 c368 (.A0(clknet_1_0__leaf_net256),
    .A1(net242),
    .A2(clknet_1_1__leaf_net248),
    .A3(clknet_1_1__leaf_net246),
    .S0(clknet_1_1__leaf_net676),
    .S1(clknet_1_1__leaf_net711),
    .X(net257));
 sky130_fd_sc_hd__a41o_1 c369 (.A1(clknet_1_0__leaf_net256),
    .A2(net650),
    .A3(clknet_1_1__leaf_net654),
    .A4(net927),
    .B1(net892),
    .X(net258));
 sky130_fd_sc_hd__mux4_1 c370 (.A0(net650),
    .A1(net653),
    .A2(net661),
    .A3(clknet_1_1__leaf_net676),
    .S0(clknet_1_1__leaf_net711),
    .S1(net892),
    .X(net259));
 sky130_fd_sc_hd__mux4_1 c371 (.A0(clknet_1_1__leaf_net244),
    .A1(clknet_1_0__leaf_net259),
    .A2(clknet_1_1__leaf_net249),
    .A3(clknet_1_1__leaf_net256),
    .S0(net661),
    .S1(net892),
    .X(net260));
 sky130_fd_sc_hd__mux4_1 c372 (.A0(clknet_1_0__leaf_net259),
    .A1(clknet_1_1__leaf_net256),
    .A2(net242),
    .A3(net661),
    .S0(net670),
    .S1(net892),
    .X(net261));
 sky130_fd_sc_hd__a41o_1 c373 (.A1(clknet_1_1__leaf_net256),
    .A2(clknet_1_1__leaf_net259),
    .A3(net661),
    .A4(net670),
    .B1(net671),
    .X(net262));
 sky130_fd_sc_hd__dfbbn_2 c396 (.CLK_N(clknet_4_4_0_clk),
    .D(clknet_1_1__leaf_net166),
    .RESET_B(net694),
    .SET_B(clknet_1_0__leaf_net710),
    .Q(net264),
    .Q_N(net263));
 sky130_fd_sc_hd__a41o_1 c397 (.A1(net264),
    .A2(clknet_1_1__leaf_net166),
    .A3(net648),
    .A4(net694),
    .B1(clknet_1_0__leaf_net710),
    .X(net265));
 sky130_fd_sc_hd__sdfrbp_2 c398 (.CLK(clknet_4_4_0_clk),
    .D(net264),
    .RESET_B(clknet_1_1__leaf_net166),
    .SCD(net613),
    .SCE(clknet_1_0__leaf_net710),
    .Q(net267),
    .Q_N(net266));
 sky130_fd_sc_hd__a41o_1 c399 (.A1(net264),
    .A2(net267),
    .A3(clknet_1_1__leaf_net166),
    .B1(clknet_1_0__leaf_net710),
    .X(net268));
 sky130_fd_sc_hd__a31o_1 c400 (.A1(net263),
    .A2(net267),
    .A3(net613),
    .B1(net648),
    .X(net269));
 sky130_fd_sc_hd__a31o_1 c401 (.A1(net918),
    .A2(net263),
    .A3(net267),
    .B1(net612),
    .X(net270));
 sky130_fd_sc_hd__a41o_1 c402 (.A1(net270),
    .A2(net918),
    .A3(net263),
    .A4(net267),
    .B1(net613),
    .X(net271));
 sky130_fd_sc_hd__a41o_2 c403 (.A1(net918),
    .A2(net271),
    .A3(net263),
    .A4(net270),
    .B1(net613),
    .X(net272));
 sky130_fd_sc_hd__a41o_1 c404 (.A1(net271),
    .A2(net272),
    .A3(net263),
    .A4(net918),
    .B1(net613),
    .X(net273));
 sky130_fd_sc_hd__mux4_1 c405 (.A0(net264),
    .A1(net270),
    .A2(net273),
    .A3(net918),
    .S0(net272),
    .S1(net612),
    .X(net274));
 sky130_fd_sc_hd__mux4_2 c406 (.A0(net274),
    .A1(net918),
    .A2(net273),
    .A3(net263),
    .S0(net272),
    .S1(net613),
    .X(net275));
 sky130_fd_sc_hd__mux4_2 c407 (.A0(net275),
    .A1(net270),
    .A2(net263),
    .A3(net271),
    .S0(net267),
    .S1(net269),
    .X(net276));
 sky130_fd_sc_hd__mux4_2 c408 (.A0(net273),
    .A1(net276),
    .A2(net918),
    .A3(net275),
    .S0(net271),
    .S1(net613),
    .X(net277));
 sky130_fd_sc_hd__mux4_2 c409 (.A0(net277),
    .A1(net274),
    .A2(net918),
    .A3(net264),
    .S0(net272),
    .S1(net612),
    .X(net278));
 sky130_fd_sc_hd__mux4_1 c410 (.A0(net267),
    .A1(net276),
    .A2(net278),
    .A3(net277),
    .S0(net264),
    .S1(net612),
    .X(net279));
 sky130_fd_sc_hd__mux4_1 c411 (.A0(net278),
    .A1(net275),
    .A2(net279),
    .A3(net918),
    .S0(net277),
    .S1(net612),
    .X(net280));
 sky130_fd_sc_hd__mux4_1 c412 (.A0(net279),
    .A1(net274),
    .A2(net277),
    .A3(net278),
    .S0(net264),
    .S1(net612),
    .X(net281));
 sky130_fd_sc_hd__mux4_2 c413 (.A0(net272),
    .A1(net278),
    .A2(net271),
    .A3(net277),
    .S0(net275),
    .S1(net612),
    .X(net282));
 sky130_fd_sc_hd__mux4_1 c414 (.A0(net281),
    .A1(net280),
    .A2(net282),
    .A3(net918),
    .S0(net277),
    .S1(net612),
    .X(net283));
 sky130_fd_sc_hd__mux4_2 c415 (.A0(net283),
    .A1(net269),
    .A2(net280),
    .A3(net282),
    .S0(net278),
    .S1(net613),
    .X(net284));
 sky130_fd_sc_hd__mux4_1 c416 (.A0(net280),
    .A1(net282),
    .A2(net283),
    .A3(net277),
    .S0(net284),
    .S1(net278),
    .X(net285));
 sky130_fd_sc_hd__mux4_2 c417 (.A0(net276),
    .A1(net285),
    .A2(net283),
    .A3(net284),
    .S0(net267),
    .S1(net282),
    .X(net286));
 sky130_fd_sc_hd__sdfbbn_1 c418 (.CLK_N(clknet_4_5_0_clk),
    .D(net267),
    .RESET_B(net806),
    .SCD(clknet_1_1__leaf_net194),
    .SCE(net174),
    .SET_B(clknet_1_1__leaf_net193),
    .Q(net288),
    .Q_N(net287));
 sky130_fd_sc_hd__sdfbbp_1 c419 (.CLK(clknet_4_4_0_clk),
    .D(clknet_1_0__leaf_net194),
    .RESET_B(net288),
    .SCD(net174),
    .SCE(net284),
    .SET_B(net266),
    .Q(net290),
    .Q_N(net289));
 sky130_fd_sc_hd__a41o_2 c420 (.A1(net284),
    .A2(net290),
    .A3(net288),
    .A4(net266),
    .B1(net174),
    .X(net291));
 sky130_fd_sc_hd__mux4_1 c421 (.A0(net290),
    .A1(net284),
    .A2(net291),
    .A3(net287),
    .S0(clknet_1_1__leaf_net193),
    .S1(net286),
    .X(net292));
 sky130_fd_sc_hd__sdfbbn_1 c422 (.CLK_N(clknet_4_4_0_clk),
    .D(clknet_1_0__leaf_net292),
    .RESET_B(net290),
    .SCD(net291),
    .SCE(net286),
    .SET_B(net944),
    .Q(net294),
    .Q_N(net293));
 sky130_fd_sc_hd__mux4_1 c423 (.A0(net291),
    .A1(net293),
    .A2(net286),
    .A3(net289),
    .S0(net287),
    .S1(clknet_1_1__leaf_net292),
    .X(net295));
 sky130_fd_sc_hd__mux4_1 c424 (.A0(net291),
    .A1(clknet_1_1__leaf_net292),
    .A2(net289),
    .A3(net293),
    .S0(net287),
    .S1(net738),
    .X(net296));
 sky130_fd_sc_hd__mux4_1 c425 (.A0(clknet_1_1__leaf_net292),
    .A1(net293),
    .A2(net289),
    .A3(net291),
    .S0(net713),
    .S1(net738),
    .X(net297));
 sky130_fd_sc_hd__mux4_1 c426 (.A0(clknet_1_0__leaf_net292),
    .A1(net289),
    .A2(net291),
    .A3(net293),
    .S0(net713),
    .S1(net740),
    .X(net298));
 sky130_fd_sc_hd__mux4_2 c427 (.A0(net290),
    .A1(net287),
    .A2(net291),
    .A3(net713),
    .S0(net740),
    .S1(net741),
    .X(net299));
 sky130_fd_sc_hd__mux4_1 c428 (.A0(net299),
    .A1(net288),
    .A2(clknet_1_1__leaf_net292),
    .A3(net713),
    .S0(net738),
    .S1(net739),
    .X(net300));
 sky130_fd_sc_hd__mux4_2 c429 (.A0(net294),
    .A1(net299),
    .A2(net690),
    .A3(net738),
    .S0(net739),
    .S1(net742),
    .X(net301));
 sky130_fd_sc_hd__mux4_1 c430 (.A0(net288),
    .A1(net301),
    .A2(net299),
    .A3(net690),
    .S0(net739),
    .S1(net741),
    .X(net302));
 sky130_fd_sc_hd__mux4_1 c431 (.A0(net294),
    .A1(net302),
    .A2(net299),
    .A3(net713),
    .S0(net740),
    .S1(net742),
    .X(net303));
 sky130_fd_sc_hd__mux4_1 c432 (.A0(net303),
    .A1(net294),
    .A2(net301),
    .A3(net290),
    .S0(net690),
    .S1(net740),
    .X(net304));
 sky130_fd_sc_hd__mux4_1 c433 (.A0(net301),
    .A1(net303),
    .A2(net906),
    .A3(net299),
    .S0(clknet_1_0__leaf_net292),
    .S1(net742),
    .X(net305));
 sky130_fd_sc_hd__mux4_1 c434 (.A0(net291),
    .A1(net906),
    .A2(net301),
    .A3(net303),
    .S0(net690),
    .S1(net738),
    .X(net306));
 sky130_fd_sc_hd__mux4_1 c435 (.A0(net294),
    .A1(net906),
    .A2(net306),
    .A3(net303),
    .S0(net669),
    .S1(net741),
    .X(net307));
 sky130_fd_sc_hd__mux4_1 c436 (.A0(net306),
    .A1(net302),
    .A2(net906),
    .A3(net299),
    .S0(net669),
    .S1(net739),
    .X(net308));
 sky130_fd_sc_hd__mux4_1 c437 (.A0(net301),
    .A1(net291),
    .A2(net907),
    .A3(net662),
    .S0(net669),
    .S1(net699),
    .X(net309));
 sky130_fd_sc_hd__mux4_1 c438 (.A0(net309),
    .A1(net907),
    .A2(net662),
    .A3(net699),
    .S0(net738),
    .S1(net742),
    .X(net310));
 sky130_fd_sc_hd__mux4_1 c439 (.A0(net302),
    .A1(net309),
    .A2(net301),
    .A3(net907),
    .S0(net662),
    .S1(net699),
    .X(net311));
 sky130_fd_sc_hd__a41o_1 c440 (.A1(net906),
    .A2(net97),
    .A3(net649),
    .A4(net686),
    .B1(net928),
    .X(net312));
 sky130_fd_sc_hd__sdfbbn_1 c441 (.CLK_N(clknet_4_3_0_clk),
    .D(net906),
    .RESET_B(net903),
    .SCD(net284),
    .SCE(net695),
    .SET_B(net928),
    .Q(net314),
    .Q_N(net313));
 sky130_fd_sc_hd__sdfrbp_2 c442 (.CLK(clknet_4_6_0_clk),
    .D(net314),
    .RESET_B(net903),
    .SCD(net695),
    .SCE(net737),
    .Q(net316),
    .Q_N(net315));
 sky130_fd_sc_hd__a41o_1 c443 (.A1(net314),
    .A2(net316),
    .A3(net903),
    .A4(net695),
    .B1(net737),
    .X(net317));
 sky130_fd_sc_hd__a41o_1 c444 (.A1(net316),
    .A2(net312),
    .A3(net313),
    .A4(net881),
    .B1(net737),
    .X(net318));
 sky130_fd_sc_hd__mux4_1 c445 (.A0(net903),
    .A1(net314),
    .A2(net315),
    .A3(net881),
    .S0(net934),
    .S1(net737),
    .X(net319));
 sky130_fd_sc_hd__mux4_1 c446 (.A0(net903),
    .A1(net313),
    .A2(net315),
    .A3(net881),
    .S0(net934),
    .S1(net926),
    .X(net320));
 sky130_fd_sc_hd__mux4_1 c447 (.A0(net314),
    .A1(net903),
    .A2(net315),
    .A3(net668),
    .S0(net881),
    .S1(net926),
    .X(net321));
 sky130_fd_sc_hd__mux4_1 c448 (.A0(net903),
    .A1(net315),
    .A2(net313),
    .A3(net934),
    .S0(net719),
    .S1(net925),
    .X(net322));
 sky130_fd_sc_hd__mux4_1 c449 (.A0(net315),
    .A1(net312),
    .A2(net700),
    .A3(net934),
    .S0(net925),
    .S1(net744),
    .X(net323));
 sky130_fd_sc_hd__mux4_1 c450 (.A0(net315),
    .A1(net903),
    .A2(net668),
    .A3(net719),
    .S0(net925),
    .S1(net745),
    .X(net324));
 sky130_fd_sc_hd__mux4_1 c451 (.A0(net315),
    .A1(net903),
    .A2(net934),
    .A3(net925),
    .S0(net744),
    .S1(net745),
    .X(net325));
 sky130_fd_sc_hd__mux4_1 c452 (.A0(net316),
    .A1(net906),
    .A2(net312),
    .A3(net744),
    .S0(net745),
    .S1(clknet_1_0__leaf_net746),
    .X(net326));
 sky130_fd_sc_hd__mux4_1 c453 (.A0(net906),
    .A1(net315),
    .A2(net926),
    .A3(net744),
    .S0(net745),
    .S1(clknet_1_0__leaf_net746),
    .X(net327));
 sky130_fd_sc_hd__mux4_1 c454 (.A0(net316),
    .A1(clknet_1_1__leaf_net327),
    .A2(net700),
    .A3(net744),
    .S0(net745),
    .S1(clknet_1_1__leaf_net746),
    .X(net328));
 sky130_fd_sc_hd__mux4_1 c455 (.A0(clknet_1_0__leaf_net327),
    .A1(net668),
    .A2(net934),
    .A3(net925),
    .S0(net745),
    .S1(clknet_1_1__leaf_net746),
    .X(net329));
 sky130_fd_sc_hd__mux4_1 c456 (.A0(clknet_1_1__leaf_net327),
    .A1(net316),
    .A2(net687),
    .A3(net745),
    .S0(clknet_1_1__leaf_net746),
    .S1(clknet_1_1__leaf_net747),
    .X(net330));
 sky130_fd_sc_hd__mux4_1 c457 (.A0(net312),
    .A1(net316),
    .A2(clknet_1_1__leaf_net327),
    .A3(net700),
    .S0(net745),
    .S1(clknet_1_1__leaf_net747),
    .X(net331));
 sky130_fd_sc_hd__mux4_1 c458 (.A0(clknet_1_1__leaf_net327),
    .A1(net903),
    .A2(net687),
    .A3(net701),
    .S0(net745),
    .S1(clknet_1_1__leaf_net747),
    .X(net332));
 sky130_fd_sc_hd__mux4_1 c459 (.A0(net313),
    .A1(clknet_1_0__leaf_net327),
    .A2(net719),
    .A3(net744),
    .S0(clknet_1_1__leaf_net746),
    .S1(clknet_1_0__leaf_net747),
    .X(net333));
 sky130_fd_sc_hd__mux4_1 c460 (.A0(net316),
    .A1(net679),
    .A2(net701),
    .A3(net744),
    .S0(clknet_1_0__leaf_net746),
    .S1(clknet_1_0__leaf_net747),
    .X(net334));
 sky130_fd_sc_hd__mux4_1 c461 (.A0(net334),
    .A1(clknet_1_0__leaf_net327),
    .A2(net316),
    .A3(net679),
    .S0(net925),
    .S1(clknet_1_0__leaf_net747),
    .X(net335));
 sky130_fd_sc_hd__sdfbbp_1 c462 (.CLK(clknet_4_8_0_clk),
    .D(clknet_1_0__leaf_net238),
    .RESET_B(clknet_1_1__leaf_net219),
    .SCD(net935),
    .SCE(clknet_1_1__leaf_net889),
    .SET_B(net925),
    .Q(net337),
    .Q_N(net336));
 sky130_fd_sc_hd__a41o_1 c463 (.A1(net337),
    .A2(clknet_1_1__leaf_net219),
    .A3(clknet_1_0__leaf_net238),
    .A4(net719),
    .B1(net925),
    .X(net338));
 sky130_fd_sc_hd__a41o_1 c464 (.A1(net337),
    .A2(clknet_1_1__leaf_net238),
    .A3(clknet_1_1__leaf_net219),
    .B1(net925),
    .X(net339));
 sky130_fd_sc_hd__sdfrtn_1 c465 (.CLK_N(clknet_4_8_0_clk),
    .D(clknet_1_0__leaf_net238),
    .RESET_B(net337),
    .SCD(net632),
    .SCE(net925),
    .Q(net340));
 sky130_fd_sc_hd__sdfrtp_4 c466 (.CLK(clknet_4_8_0_clk),
    .D(net340),
    .RESET_B(net337),
    .SCD(clknet_1_0__leaf_net238),
    .SCE(net632),
    .Q(net341));
 sky130_fd_sc_hd__a31o_1 c467 (.A1(net341),
    .A2(net337),
    .A3(net340),
    .B1(net632),
    .X(net342));
 sky130_fd_sc_hd__a41o_1 c468 (.A1(net342),
    .A2(net336),
    .A3(net340),
    .A4(net341),
    .B1(net632),
    .X(net343));
 sky130_fd_sc_hd__mux4_1 c469 (.A0(net341),
    .A1(net340),
    .A2(net336),
    .A3(net342),
    .S0(net632),
    .S1(clknet_1_1__leaf_net889),
    .X(net344));
 sky130_fd_sc_hd__a41o_1 c470 (.A1(net343),
    .A2(clknet_1_0__leaf_net344),
    .A3(net336),
    .A4(net342),
    .B1(net632),
    .X(net345));
 sky130_fd_sc_hd__mux4_1 c471 (.A0(net342),
    .A1(clknet_1_0__leaf_net344),
    .A2(clknet_1_0__leaf_net345),
    .A3(net343),
    .S0(net340),
    .S1(net336),
    .X(net346));
 sky130_fd_sc_hd__mux4_1 c472 (.A0(clknet_1_0__leaf_net346),
    .A1(clknet_1_0__leaf_net345),
    .A2(net343),
    .A3(net341),
    .S0(net336),
    .S1(net340),
    .X(net347));
 sky130_fd_sc_hd__mux4_1 c473 (.A0(net340),
    .A1(clknet_1_1__leaf_net346),
    .A2(clknet_1_0__leaf_net347),
    .A3(net342),
    .S0(clknet_1_1__leaf_net345),
    .S1(net336),
    .X(net348));
 sky130_fd_sc_hd__mux4_1 c474 (.A0(clknet_1_0__leaf_net347),
    .A1(clknet_1_1__leaf_net346),
    .A2(clknet_1_1__leaf_net345),
    .A3(net336),
    .S0(net341),
    .S1(net340),
    .X(net349));
 sky130_fd_sc_hd__mux4_1 c475 (.A0(net343),
    .A1(net337),
    .A2(clknet_1_1__leaf_net347),
    .A3(net340),
    .S0(clknet_1_0__leaf_net346),
    .S1(net632),
    .X(net887));
 sky130_fd_sc_hd__mux4_1 c476 (.A0(net337),
    .A1(clknet_1_0__leaf_net887),
    .A2(net343),
    .A3(clknet_1_1__leaf_net347),
    .S0(net341),
    .S1(clknet_1_0__leaf_net349),
    .X(net350));
 sky130_fd_sc_hd__a41o_1 c477 (.A1(clknet_1_1__leaf_net344),
    .A2(clknet_1_0__leaf_net350),
    .A3(net342),
    .A4(net341),
    .B1(net632),
    .X(net351));
 sky130_fd_sc_hd__mux4_1 c478 (.A0(clknet_1_1__leaf_net345),
    .A1(clknet_1_0__leaf_net349),
    .A2(clknet_1_0__leaf_net347),
    .A3(clknet_1_0__leaf_net351),
    .S0(net340),
    .S1(net341),
    .X(net352));
 sky130_fd_sc_hd__mux4_1 c479 (.A0(clknet_1_0__leaf_net352),
    .A1(net342),
    .A2(clknet_1_1__leaf_net351),
    .A3(clknet_1_1__leaf_net346),
    .S0(clknet_1_1__leaf_net349),
    .S1(clknet_1_1__leaf_net887),
    .X(net353));
 sky130_fd_sc_hd__mux4_1 c480 (.A0(net341),
    .A1(clknet_1_1__leaf_net350),
    .A2(clknet_1_0__leaf_net346),
    .A3(clknet_1_0__leaf_net887),
    .S0(clknet_1_1__leaf_net344),
    .S1(clknet_1_0__leaf_net351),
    .X(net354));
 sky130_fd_sc_hd__mux4_1 c481 (.A0(clknet_1_1__leaf_net348),
    .A1(clknet_1_0__leaf_net353),
    .A2(clknet_1_0__leaf_net354),
    .A3(clknet_1_1__leaf_net349),
    .S0(clknet_1_1__leaf_net352),
    .S1(clknet_1_1__leaf_net351),
    .X(net355));
 sky130_fd_sc_hd__mux4_1 c482 (.A0(clknet_1_1__leaf_net349),
    .A1(clknet_1_0__leaf_net351),
    .A2(clknet_1_0__leaf_net355),
    .A3(clknet_1_0__leaf_net348),
    .S0(clknet_1_1__leaf_net344),
    .S1(clknet_1_0__leaf_net354),
    .X(net356));
 sky130_fd_sc_hd__mux4_1 c483 (.A0(clknet_1_1__leaf_net355),
    .A1(clknet_1_1__leaf_net354),
    .A2(clknet_1_1__leaf_net353),
    .A3(clknet_1_1__leaf_net351),
    .S0(clknet_1_1__leaf_net887),
    .S1(net719),
    .X(net357));
 sky130_fd_sc_hd__a41o_1 c484 (.A1(clknet_1_1__leaf_net887),
    .A2(clknet_1_1__leaf_net357),
    .A3(clknet_1_1__leaf_net356),
    .A4(net896),
    .B1(net927),
    .X(net883));
 sky130_fd_sc_hd__sdfbbn_1 c485 (.CLK_N(clknet_4_10_0_clk),
    .D(clknet_1_0__leaf_net883),
    .RESET_B(clknet_1_1__leaf_net142),
    .SCD(clknet_1_1__leaf_net887),
    .SCE(net896),
    .SET_B(net927),
    .Q(net359),
    .Q_N(net358));
 sky130_fd_sc_hd__a41o_1 c486 (.A1(net359),
    .A2(clknet_1_0__leaf_net883),
    .A3(clknet_1_0__leaf_net356),
    .A4(clknet_1_1__leaf_net887),
    .B1(net927),
    .X(net360));
 sky130_fd_sc_hd__mux4_1 c487 (.A0(clknet_1_1__leaf_net360),
    .A1(clknet_1_1__leaf_net883),
    .A2(net359),
    .A3(clknet_1_1__leaf_net887),
    .S0(net927),
    .S1(net892),
    .X(net361));
 sky130_fd_sc_hd__a41o_1 c488 (.A1(clknet_1_0__leaf_net883),
    .A2(net359),
    .A3(clknet_1_0__leaf_net361),
    .A4(clknet_1_1__leaf_net357),
    .B1(clknet_1_1__leaf_net360),
    .X(net362));
 sky130_fd_sc_hd__a41o_1 c489 (.A1(clknet_1_0__leaf_net361),
    .A2(clknet_1_1__leaf_net362),
    .A3(clknet_1_0__leaf_net360),
    .A4(clknet_1_0__leaf_net883),
    .B1(net358),
    .X(net363));
 sky130_fd_sc_hd__mux4_1 c490 (.A0(clknet_1_1__leaf_net361),
    .A1(clknet_1_1__leaf_net883),
    .A2(clknet_1_1__leaf_net360),
    .A3(net358),
    .S0(clknet_1_1__leaf_net363),
    .S1(net927),
    .X(net364));
 sky130_fd_sc_hd__mux4_1 c491 (.A0(net359),
    .A1(clknet_1_1__leaf_net361),
    .A2(clknet_1_0__leaf_net363),
    .A3(clknet_1_0__leaf_net883),
    .S0(clknet_1_0__leaf_net362),
    .S1(clknet_1_0__leaf_net360),
    .X(net365));
 sky130_fd_sc_hd__mux4_1 c492 (.A0(clknet_1_1__leaf_net365),
    .A1(clknet_1_1__leaf_net361),
    .A2(clknet_1_1__leaf_net360),
    .A3(net358),
    .S0(net927),
    .S1(net892),
    .X(net366));
 sky130_fd_sc_hd__mux4_1 c493 (.A0(clknet_1_0__leaf_net360),
    .A1(clknet_1_0__leaf_net363),
    .A2(clknet_1_1__leaf_net366),
    .A3(clknet_1_0__leaf_net364),
    .S0(clknet_1_0__leaf_net361),
    .S1(clknet_1_1__leaf_net365),
    .X(net367));
 sky130_fd_sc_hd__mux4_1 c494 (.A0(net359),
    .A1(clknet_1_0__leaf_net360),
    .A2(clknet_1_0__leaf_net364),
    .A3(clknet_1_0__leaf_net366),
    .S0(clknet_1_0__leaf_net365),
    .S1(clknet_1_0__leaf_net883),
    .X(net368));
 sky130_fd_sc_hd__mux4_1 c495 (.A0(clknet_1_0__leaf_net362),
    .A1(clknet_1_1__leaf_net360),
    .A2(clknet_1_1__leaf_net366),
    .A3(clknet_1_1__leaf_net361),
    .S0(clknet_1_1__leaf_net890),
    .S1(net358),
    .X(net369));
 sky130_fd_sc_hd__mux4_1 c496 (.A0(clknet_1_1__leaf_net364),
    .A1(clknet_1_1__leaf_net366),
    .A2(clknet_1_1__leaf_net369),
    .A3(net358),
    .S0(clknet_1_1__leaf_net360),
    .S1(clknet_1_1__leaf_net365),
    .X(net370));
 sky130_fd_sc_hd__mux4_1 c497 (.A0(clknet_1_1__leaf_net369),
    .A1(clknet_1_1__leaf_net367),
    .A2(clknet_1_1__leaf_net370),
    .A3(clknet_1_1__leaf_net361),
    .S0(clknet_1_1__leaf_net366),
    .S1(clknet_1_1__leaf_net360),
    .X(net371));
 sky130_fd_sc_hd__mux4_1 c498 (.A0(clknet_1_1__leaf_net363),
    .A1(clknet_1_1__leaf_net365),
    .A2(clknet_1_1__leaf_net366),
    .A3(clknet_1_1__leaf_net369),
    .S0(clknet_1_1__leaf_net370),
    .S1(clknet_1_0__leaf_net884),
    .X(net372));
 sky130_fd_sc_hd__mux4_1 c499 (.A0(clknet_1_0__leaf_net367),
    .A1(clknet_1_0__leaf_net369),
    .A2(clknet_1_0__leaf_net360),
    .A3(clknet_1_0__leaf_net370),
    .S0(clknet_1_0__leaf_net365),
    .S1(clknet_1_0__leaf_net884),
    .X(net373));
 sky130_fd_sc_hd__mux4_1 c500 (.A0(clknet_1_0__leaf_net366),
    .A1(clknet_1_0__leaf_net369),
    .A2(clknet_1_0__leaf_net370),
    .A3(clknet_1_0__leaf_net360),
    .S0(net671),
    .S1(net692),
    .X(net374));
 sky130_fd_sc_hd__mux4_1 c501 (.A0(clknet_1_0__leaf_net370),
    .A1(clknet_1_0__leaf_net365),
    .A2(clknet_1_0__leaf_net361),
    .A3(net671),
    .S0(net692),
    .S1(net933),
    .X(net375));
 sky130_fd_sc_hd__mux4_1 c502 (.A0(clknet_1_0__leaf_net366),
    .A1(clknet_1_0__leaf_net367),
    .A2(clknet_1_0__leaf_net369),
    .A3(net667),
    .S0(net692),
    .S1(net933),
    .X(net376));
 sky130_fd_sc_hd__mux4_1 c503 (.A0(net368),
    .A1(clknet_1_0__leaf_net376),
    .A2(clknet_1_0__leaf_net370),
    .A3(clknet_1_0__leaf_net369),
    .S0(net667),
    .S1(clknet_1_0__leaf_net884),
    .X(net377));
 sky130_fd_sc_hd__mux4_1 c504 (.A0(net359),
    .A1(clknet_1_0__leaf_net376),
    .A2(clknet_1_0__leaf_net366),
    .A3(net667),
    .S0(net670),
    .S1(net692),
    .X(net378));
 sky130_fd_sc_hd__mux4_1 c505 (.A0(clknet_1_1__leaf_net376),
    .A1(clknet_1_0__leaf_net370),
    .A2(net667),
    .A3(net670),
    .S0(net692),
    .S1(net933),
    .X(net379));
 sky130_fd_sc_hd__a31o_1 c528 (.A1(net286),
    .A2(net284),
    .A3(net266),
    .B1(net43),
    .X(net380));
 sky130_fd_sc_hd__a31o_2 c529 (.A1(net912),
    .A2(net286),
    .A3(net267),
    .B1(net284),
    .X(net381));
 sky130_fd_sc_hd__a41o_2 c530 (.A1(net912),
    .A2(net381),
    .A3(net284),
    .A4(net266),
    .B1(net286),
    .X(net382));
 sky130_fd_sc_hd__a41o_1 c531 (.A1(net382),
    .A2(net381),
    .A3(net912),
    .A4(net266),
    .B1(net284),
    .X(net383));
 sky130_fd_sc_hd__a41o_1 c532 (.A1(net381),
    .A2(net912),
    .A3(net382),
    .A4(net905),
    .B1(net266),
    .X(net384));
 sky130_fd_sc_hd__sdfbbn_2 c533 (.CLK_N(clknet_4_5_0_clk),
    .D(net384),
    .RESET_B(net382),
    .SCD(net912),
    .SCE(net905),
    .SET_B(net381),
    .Q(net386),
    .Q_N(net385));
 sky130_fd_sc_hd__mux4_1 c534 (.A0(net383),
    .A1(net386),
    .A2(net384),
    .A3(net381),
    .S0(net912),
    .S1(net382),
    .X(net387));
 sky130_fd_sc_hd__mux4_2 c535 (.A0(net382),
    .A1(net386),
    .A2(net381),
    .A3(net912),
    .S0(net905),
    .S1(net689),
    .X(net388));
 sky130_fd_sc_hd__mux4_2 c536 (.A0(net905),
    .A1(net386),
    .A2(net912),
    .A3(net381),
    .S0(net382),
    .S1(net689),
    .X(net389));
 sky130_fd_sc_hd__mux4_1 c537 (.A0(net384),
    .A1(net389),
    .A2(net912),
    .A3(net385),
    .S0(net381),
    .S1(net689),
    .X(net390));
 sky130_fd_sc_hd__mux4_1 c538 (.A0(net389),
    .A1(net386),
    .A2(net905),
    .A3(net912),
    .S0(net689),
    .S1(net749),
    .X(net391));
 sky130_fd_sc_hd__mux4_1 c539 (.A0(net381),
    .A1(net384),
    .A2(net386),
    .A3(net905),
    .S0(net380),
    .S1(net947),
    .X(net392));
 sky130_fd_sc_hd__mux4_1 c540 (.A0(net386),
    .A1(net389),
    .A2(net381),
    .A3(net668),
    .S0(net749),
    .S1(net750),
    .X(net393));
 sky130_fd_sc_hd__mux4_1 c541 (.A0(net384),
    .A1(net905),
    .A2(net385),
    .A3(net704),
    .S0(net748),
    .S1(net751),
    .X(net394));
 sky130_fd_sc_hd__mux4_1 c542 (.A0(net386),
    .A1(net904),
    .A2(net389),
    .A3(net704),
    .S0(net751),
    .S1(net752),
    .X(net395));
 sky130_fd_sc_hd__mux4_1 c543 (.A0(net905),
    .A1(net668),
    .A2(net748),
    .A3(net750),
    .S0(net752),
    .S1(net924),
    .X(net396));
 sky130_fd_sc_hd__mux4_1 c544 (.A0(net905),
    .A1(net382),
    .A2(net704),
    .A3(net749),
    .S0(net750),
    .S1(net752),
    .X(net397));
 sky130_fd_sc_hd__mux4_1 c545 (.A0(net397),
    .A1(net396),
    .A2(net748),
    .A3(net751),
    .S0(net752),
    .S1(net924),
    .X(net398));
 sky130_fd_sc_hd__mux4_1 c546 (.A0(net388),
    .A1(net397),
    .A2(net703),
    .A3(net704),
    .S0(net752),
    .S1(net924),
    .X(net399));
 sky130_fd_sc_hd__mux4_1 c547 (.A0(net396),
    .A1(net386),
    .A2(net397),
    .A3(clknet_1_0__leaf_net677),
    .S0(net703),
    .S1(net752),
    .X(net400));
 sky130_fd_sc_hd__a41o_1 c548 (.A1(net397),
    .A2(net389),
    .A3(net905),
    .A4(clknet_1_0__leaf_net677),
    .B1(net924),
    .X(net401));
 sky130_fd_sc_hd__a41o_1 c549 (.A1(net668),
    .A2(clknet_1_0__leaf_net677),
    .A3(net751),
    .A4(net752),
    .B1(net924),
    .X(net402));
 sky130_fd_sc_hd__mux4_1 c550 (.A0(clknet_1_0__leaf_net402),
    .A1(net907),
    .A2(net266),
    .A3(net385),
    .S0(net904),
    .S1(net923),
    .X(net403));
 sky130_fd_sc_hd__sdfbbp_1 c551 (.CLK(clknet_4_5_0_clk),
    .D(net907),
    .RESET_B(clknet_1_1__leaf_net184),
    .SCD(net904),
    .SCE(net923),
    .SET_B(net922),
    .Q(net405),
    .Q_N(net404));
 sky130_fd_sc_hd__sdfbbn_1 c552 (.CLK_N(clknet_4_7_0_clk),
    .D(net404),
    .RESET_B(net385),
    .SCD(net904),
    .SCE(net923),
    .SET_B(net922),
    .Q(net407),
    .Q_N(net406));
 sky130_fd_sc_hd__mux4_1 c553 (.A0(net407),
    .A1(net404),
    .A2(net385),
    .A3(net904),
    .S0(net923),
    .S1(net922),
    .X(net408));
 sky130_fd_sc_hd__mux4_1 c554 (.A0(net407),
    .A1(net404),
    .A2(clknet_1_0__leaf_net402),
    .A3(net904),
    .S0(net712),
    .S1(net922),
    .X(net409));
 sky130_fd_sc_hd__mux4_2 c555 (.A0(net407),
    .A1(net404),
    .A2(net699),
    .A3(net702),
    .S0(net712),
    .S1(net754),
    .X(net410));
 sky130_fd_sc_hd__mux4_1 c556 (.A0(net405),
    .A1(net407),
    .A2(net907),
    .A3(net410),
    .S0(net712),
    .S1(net922),
    .X(net411));
 sky130_fd_sc_hd__mux4_1 c557 (.A0(net411),
    .A1(net405),
    .A2(net410),
    .A3(net406),
    .S0(net949),
    .S1(net922),
    .X(net412));
 sky130_fd_sc_hd__mux4_1 c558 (.A0(net407),
    .A1(net937),
    .A2(net411),
    .A3(net712),
    .S0(net922),
    .S1(net755),
    .X(net413));
 sky130_fd_sc_hd__mux4_2 c559 (.A0(net407),
    .A1(net907),
    .A2(net938),
    .A3(net713),
    .S0(net755),
    .S1(net756),
    .X(net414));
 sky130_fd_sc_hd__mux4_1 c560 (.A0(net414),
    .A1(net938),
    .A2(net406),
    .A3(net754),
    .S0(net755),
    .S1(net756),
    .X(net415));
 sky130_fd_sc_hd__mux4_1 c561 (.A0(net414),
    .A1(net404),
    .A2(net406),
    .A3(net949),
    .S0(net922),
    .S1(net756),
    .X(net416));
 sky130_fd_sc_hd__mux4_2 c562 (.A0(net410),
    .A1(net405),
    .A2(net406),
    .A3(net755),
    .S0(net756),
    .S1(net758),
    .X(net417));
 sky130_fd_sc_hd__mux4_2 c563 (.A0(net417),
    .A1(net406),
    .A2(net662),
    .A3(net755),
    .S0(net756),
    .S1(net757),
    .X(net418));
 sky130_fd_sc_hd__mux4_1 c564 (.A0(net410),
    .A1(net418),
    .A2(net417),
    .A3(net906),
    .S0(net755),
    .S1(net757),
    .X(net419));
 sky130_fd_sc_hd__mux4_1 c565 (.A0(net419),
    .A1(net418),
    .A2(net417),
    .A3(net405),
    .S0(net406),
    .S1(net757),
    .X(net420));
 sky130_fd_sc_hd__mux4_1 c566 (.A0(net419),
    .A1(net662),
    .A2(net684),
    .A3(net702),
    .S0(net922),
    .S1(net755),
    .X(net421));
 sky130_fd_sc_hd__mux4_1 c567 (.A0(net906),
    .A1(net405),
    .A2(net414),
    .A3(net418),
    .S0(net758),
    .S1(net759),
    .X(net422));
 sky130_fd_sc_hd__mux4_2 c568 (.A0(net418),
    .A1(net662),
    .A2(net922),
    .A3(net755),
    .S0(net760),
    .S1(net921),
    .X(net423));
 sky130_fd_sc_hd__mux4_1 c569 (.A0(net411),
    .A1(net417),
    .A2(net423),
    .A3(net756),
    .S0(net758),
    .S1(net760),
    .X(net424));
 sky130_fd_sc_hd__mux4_1 c570 (.A0(net414),
    .A1(net684),
    .A2(net712),
    .A3(net756),
    .S0(net760),
    .S1(net921),
    .X(net425));
 sky130_fd_sc_hd__a41o_1 c571 (.A1(net423),
    .A2(net684),
    .A3(net688),
    .A4(net758),
    .B1(net921),
    .X(net426));
 sky130_fd_sc_hd__a41o_2 c572 (.A1(net688),
    .A2(net700),
    .A3(net926),
    .A4(net923),
    .B1(net921),
    .X(net427));
 sky130_fd_sc_hd__a41o_2 c573 (.A1(net427),
    .A2(net266),
    .A3(net695),
    .A4(net926),
    .B1(net921),
    .X(net428));
 sky130_fd_sc_hd__a41o_2 c574 (.A1(net428),
    .A2(net427),
    .A3(net679),
    .A4(net688),
    .B1(net921),
    .X(net429));
 sky130_fd_sc_hd__a41o_2 c575 (.A1(net429),
    .A2(net428),
    .A3(net427),
    .A4(net679),
    .B1(net921),
    .X(net430));
 sky130_fd_sc_hd__a41o_1 c576 (.A1(net429),
    .A2(net430),
    .A3(net428),
    .A4(net427),
    .B1(net921),
    .X(net431));
 sky130_fd_sc_hd__mux4_2 c577 (.A0(net429),
    .A1(net430),
    .A2(net431),
    .A3(net428),
    .S0(net427),
    .S1(net926),
    .X(net432));
 sky130_fd_sc_hd__mux4_2 c578 (.A0(net430),
    .A1(net915),
    .A2(net429),
    .A3(net426),
    .S0(net431),
    .S1(net921),
    .X(net433));
 sky130_fd_sc_hd__mux4_2 c579 (.A0(net433),
    .A1(net430),
    .A2(net915),
    .A3(net431),
    .S0(net429),
    .S1(net427),
    .X(net434));
 sky130_fd_sc_hd__mux4_2 c580 (.A0(net431),
    .A1(net915),
    .A2(net433),
    .A3(net430),
    .S0(net428),
    .S1(net688),
    .X(net435));
 sky130_fd_sc_hd__mux4_2 c581 (.A0(net431),
    .A1(net435),
    .A2(net915),
    .A3(net430),
    .S0(net433),
    .S1(net429),
    .X(net436));
 sky130_fd_sc_hd__mux4_2 c582 (.A0(net436),
    .A1(net432),
    .A2(net429),
    .A3(net427),
    .S0(net435),
    .S1(net434),
    .X(net437));
 sky130_fd_sc_hd__mux4_2 c583 (.A0(net915),
    .A1(net435),
    .A2(net436),
    .A3(net433),
    .S0(net427),
    .S1(net437),
    .X(net438));
 sky130_fd_sc_hd__mux4_2 c584 (.A0(net430),
    .A1(net434),
    .A2(net438),
    .A3(net435),
    .S0(net915),
    .S1(net437),
    .X(net439));
 sky130_fd_sc_hd__mux4_2 c585 (.A0(net435),
    .A1(net438),
    .A2(net436),
    .A3(net437),
    .S0(net439),
    .S1(net432),
    .X(net440));
 sky130_fd_sc_hd__mux4_2 c586 (.A0(net437),
    .A1(net435),
    .A2(net439),
    .A3(net432),
    .S0(net440),
    .S1(net430),
    .X(net441));
 sky130_fd_sc_hd__mux4_2 c587 (.A0(net427),
    .A1(net439),
    .A2(net437),
    .A3(net441),
    .S0(net435),
    .S1(net915),
    .X(net442));
 sky130_fd_sc_hd__mux4_2 c588 (.A0(net429),
    .A1(net441),
    .A2(net439),
    .A3(net915),
    .S0(net440),
    .S1(net442),
    .X(net443));
 sky130_fd_sc_hd__mux4_2 c589 (.A0(net443),
    .A1(net440),
    .A2(net441),
    .A3(net438),
    .S0(net430),
    .S1(net442),
    .X(net444));
 sky130_fd_sc_hd__mux4_2 c590 (.A0(net441),
    .A1(net442),
    .A2(net443),
    .A3(net430),
    .S0(net438),
    .S1(net439),
    .X(net445));
 sky130_fd_sc_hd__mux4_2 c591 (.A0(net438),
    .A1(net443),
    .A2(net444),
    .A3(net441),
    .S0(net445),
    .S1(net915),
    .X(net446));
 sky130_fd_sc_hd__mux4_1 c592 (.A0(net428),
    .A1(net445),
    .A2(net446),
    .A3(net443),
    .S0(net439),
    .S1(net388),
    .X(net447));
 sky130_fd_sc_hd__mux4_2 c593 (.A0(net446),
    .A1(net441),
    .A2(net438),
    .A3(net915),
    .S0(net445),
    .S1(net701),
    .X(net448));
 sky130_fd_sc_hd__sdfbbn_1 c594 (.CLK_N(clknet_4_9_0_clk),
    .D(clknet_1_0__leaf_net357),
    .RESET_B(net448),
    .SCD(clknet_1_0__leaf_net887),
    .SCE(clknet_1_1__leaf_net238),
    .SET_B(net701),
    .Q(net450),
    .Q_N(net449));
 sky130_fd_sc_hd__a41o_1 c595 (.A1(clknet_1_0__leaf_net356),
    .A2(net450),
    .A3(clknet_1_0__leaf_net887),
    .A4(clknet_1_1__leaf_net219),
    .B1(clknet_1_0__leaf_net357),
    .X(net451));
 sky130_fd_sc_hd__a41o_1 c596 (.A1(net448),
    .A2(clknet_1_0__leaf_net451),
    .A3(net450),
    .A4(clknet_1_0__leaf_net887),
    .B1(net921),
    .X(net452));
 sky130_fd_sc_hd__a41o_1 c597 (.A1(clknet_1_0__leaf_net451),
    .A2(clknet_1_0__leaf_net452),
    .A3(net449),
    .A4(clknet_1_0__leaf_net887),
    .B1(net701),
    .X(net453));
 sky130_fd_sc_hd__sdfbbp_1 c598 (.CLK(clknet_4_9_0_clk),
    .D(clknet_1_0__leaf_net451),
    .RESET_B(net450),
    .SCD(clknet_1_0__leaf_net453),
    .SCE(clknet_1_0__leaf_net452),
    .SET_B(clknet_1_0__leaf_net887),
    .Q(net455),
    .Q_N(net454));
 sky130_fd_sc_hd__mux4_1 c599 (.A0(net448),
    .A1(clknet_1_0__leaf_net451),
    .A2(clknet_1_0__leaf_net452),
    .A3(net449),
    .S0(clknet_1_1__leaf_net453),
    .S1(net454),
    .X(net456));
 sky130_fd_sc_hd__mux4_1 c600 (.A0(clknet_1_1__leaf_net451),
    .A1(clknet_1_1__leaf_net453),
    .A2(clknet_1_0__leaf_net887),
    .A3(clknet_1_1__leaf_net452),
    .S0(net454),
    .S1(net762),
    .X(net457));
 sky130_fd_sc_hd__mux4_1 c601 (.A0(net455),
    .A1(net449),
    .A2(clknet_1_1__leaf_net453),
    .A3(clknet_1_1__leaf_net452),
    .S0(net762),
    .S1(net920),
    .X(net458));
 sky130_fd_sc_hd__mux4_1 c602 (.A0(net454),
    .A1(clknet_1_0__leaf_net453),
    .A2(clknet_1_0__leaf_net451),
    .A3(net933),
    .S0(net762),
    .S1(net920),
    .X(net459));
 sky130_fd_sc_hd__mux4_1 c603 (.A0(clknet_1_1__leaf_net452),
    .A1(clknet_1_1__leaf_net451),
    .A2(clknet_1_1__leaf_net453),
    .A3(net684),
    .S0(net762),
    .S1(net920),
    .X(net460));
 sky130_fd_sc_hd__mux4_1 c604 (.A0(clknet_1_1__leaf_net453),
    .A1(net455),
    .A2(clknet_1_1__leaf_net452),
    .A3(clknet_1_1__leaf_net451),
    .S0(net933),
    .S1(net762),
    .X(net461));
 sky130_fd_sc_hd__mux4_1 c605 (.A0(net455),
    .A1(clknet_1_0__leaf_net452),
    .A2(net684),
    .A3(net705),
    .S0(net762),
    .S1(net920),
    .X(net462));
 sky130_fd_sc_hd__mux4_1 c606 (.A0(clknet_1_1__leaf_net462),
    .A1(clknet_1_1__leaf_net453),
    .A2(net454),
    .A3(net717),
    .S0(net762),
    .S1(net763),
    .X(net463));
 sky130_fd_sc_hd__mux4_1 c607 (.A0(net455),
    .A1(clknet_1_1__leaf_net462),
    .A2(clknet_1_1__leaf_net453),
    .A3(clknet_1_1__leaf_net451),
    .S0(clknet_1_1__leaf_net452),
    .S1(net705),
    .X(net464));
 sky130_fd_sc_hd__mux4_1 c608 (.A0(clknet_1_0__leaf_net453),
    .A1(clknet_1_0__leaf_net462),
    .A2(clknet_1_0__leaf_net452),
    .A3(net705),
    .S0(net720),
    .S1(net920),
    .X(net465));
 sky130_fd_sc_hd__mux4_1 c609 (.A0(net450),
    .A1(clknet_1_0__leaf_net462),
    .A2(net881),
    .A3(net705),
    .S0(net720),
    .S1(net920),
    .X(net466));
 sky130_fd_sc_hd__mux4_1 c610 (.A0(clknet_1_1__leaf_net462),
    .A1(clknet_1_0__leaf_net451),
    .A2(net449),
    .A3(net881),
    .S0(net705),
    .S1(net920),
    .X(net467));
 sky130_fd_sc_hd__mux4_1 c611 (.A0(net455),
    .A1(clknet_1_0__leaf_net452),
    .A2(net684),
    .A3(net705),
    .S0(net720),
    .S1(net920),
    .X(net468));
 sky130_fd_sc_hd__mux4_1 c612 (.A0(clknet_1_1__leaf_net468),
    .A1(clknet_1_0__leaf_net462),
    .A2(clknet_1_0__leaf_net452),
    .A3(net705),
    .S0(net720),
    .S1(net920),
    .X(net469));
 sky130_fd_sc_hd__mux4_1 c613 (.A0(clknet_1_0__leaf_net468),
    .A1(clknet_1_0__leaf_net453),
    .A2(net671),
    .A3(net934),
    .S0(net720),
    .S1(net920),
    .X(net470));
 sky130_fd_sc_hd__mux4_1 c614 (.A0(clknet_1_0__leaf_net451),
    .A1(net687),
    .A2(net705),
    .A3(net716),
    .S0(net720),
    .S1(net762),
    .X(net471));
 sky130_fd_sc_hd__mux4_1 c615 (.A0(net471),
    .A1(clknet_1_0__leaf_net453),
    .A2(net671),
    .A3(net687),
    .S0(net705),
    .S1(net716),
    .X(net472));
 sky130_fd_sc_hd__a41o_1 c616 (.A1(clknet_1_1__leaf_net452),
    .A2(net719),
    .A3(net892),
    .A4(clknet_1_0__leaf_net884),
    .B1(net886),
    .X(net473));
 sky130_fd_sc_hd__sdfbbn_1 c617 (.CLK_N(clknet_4_11_0_clk),
    .D(clknet_1_0__leaf_net473),
    .RESET_B(net927),
    .SCD(clknet_1_0__leaf_net884),
    .SCE(net885),
    .SET_B(clknet_1_0__leaf_net764),
    .Q(net475),
    .Q_N(net474));
 sky130_fd_sc_hd__sdfbbn_1 c618 (.CLK_N(clknet_4_11_0_clk),
    .D(clknet_1_0__leaf_net473),
    .RESET_B(net475),
    .SCD(clknet_1_1__leaf_net884),
    .SCE(net885),
    .SET_B(clknet_1_0__leaf_net764),
    .Q(net477),
    .Q_N(net476));
 sky130_fd_sc_hd__sdfbbp_1 c619 (.CLK(clknet_4_10_0_clk),
    .D(clknet_1_0__leaf_net473),
    .RESET_B(net477),
    .SCD(net474),
    .SCE(clknet_1_1__leaf_net884),
    .SET_B(net885),
    .Q(net479),
    .Q_N(net478));
 sky130_fd_sc_hd__sdfbbn_1 c620 (.CLK_N(clknet_4_11_0_clk),
    .D(net475),
    .RESET_B(net477),
    .SCD(net479),
    .SCE(clknet_1_1__leaf_net473),
    .SET_B(clknet_1_0__leaf_net884),
    .Q(net882),
    .Q_N(net879));
 sky130_fd_sc_hd__mux4_1 c621 (.A0(net882),
    .A1(net475),
    .A2(net477),
    .A3(clknet_1_1__leaf_net473),
    .S0(net478),
    .S1(net885),
    .X(net480));
 sky130_fd_sc_hd__mux4_2 c622 (.A0(net882),
    .A1(net478),
    .A2(net476),
    .A3(net474),
    .S0(clknet_1_1__leaf_net473),
    .X(net628));
 sky130_fd_sc_hd__mux4_1 c623 (.A0(net479),
    .A1(clknet_1_1__leaf_net473),
    .A2(net879),
    .A3(net476),
    .S0(net474),
    .S1(clknet_1_1__leaf_net628),
    .X(net482));
 sky130_fd_sc_hd__mux4_2 c624 (.A0(net479),
    .A1(net474),
    .A2(net879),
    .A3(net476),
    .S0(clknet_1_1__leaf_net628),
    .S1(clknet_1_1__leaf_net765),
    .X(net483));
 sky130_fd_sc_hd__a41o_1 c625 (.A1(net479),
    .A2(net879),
    .A3(net476),
    .A4(clknet_1_1__leaf_net628),
    .B1(clknet_1_0__leaf_net765),
    .X(net484));
 sky130_fd_sc_hd__mux4_1 c626 (.A0(clknet_1_0__leaf_net483),
    .A1(clknet_1_0__leaf_net484),
    .A2(net475),
    .A3(net478),
    .S0(clknet_1_0__leaf_net473),
    .S1(clknet_1_0__leaf_net765),
    .X(net485));
 sky130_fd_sc_hd__mux4_2 c627 (.A0(net475),
    .A1(net882),
    .A2(clknet_1_0__leaf_net483),
    .A3(clknet_1_0__leaf_net484),
    .S0(net721),
    .S1(clknet_1_0__leaf_net765),
    .X(net486));
 sky130_fd_sc_hd__mux4_2 c628 (.A0(clknet_1_1__leaf_net484),
    .A1(clknet_1_0__leaf_net486),
    .A2(net477),
    .A3(clknet_1_0__leaf_net483),
    .S0(clknet_1_0__leaf_net628),
    .S1(net721),
    .X(net880));
 sky130_fd_sc_hd__mux4_2 c629 (.A0(clknet_1_0__leaf_net880),
    .A1(clknet_1_0__leaf_net486),
    .A2(net474),
    .A3(clknet_1_1__leaf_net484),
    .S0(clknet_1_0__leaf_net628),
    .S1(net721),
    .X(net487));
 sky130_fd_sc_hd__mux4_2 c630 (.A0(clknet_1_1__leaf_net487),
    .A1(clknet_1_1__leaf_net486),
    .A2(net476),
    .A3(clknet_1_1__leaf_net483),
    .S0(net721),
    .S1(clknet_1_1__leaf_net765),
    .X(net877));
 sky130_fd_sc_hd__mux4_2 c631 (.A0(clknet_1_0__leaf_net487),
    .A1(clknet_1_0__leaf_net877),
    .A2(net475),
    .A3(clknet_1_0__leaf_net486),
    .S0(clknet_1_0__leaf_net628),
    .S1(clknet_1_0__leaf_net765),
    .X(net488));
 sky130_fd_sc_hd__mux4_2 c632 (.A0(clknet_1_0__leaf_net488),
    .A1(clknet_1_0__leaf_net877),
    .A2(clknet_1_0__leaf_net487),
    .A3(clknet_1_1__leaf_net486),
    .S0(clknet_1_0__leaf_net484),
    .S1(net721),
    .X(net489));
 sky130_fd_sc_hd__mux4_2 c633 (.A0(net477),
    .A1(clknet_1_0__leaf_net880),
    .A2(clknet_1_1__leaf_net488),
    .A3(clknet_1_1__leaf_net877),
    .S0(clknet_1_0__leaf_net489),
    .S1(clknet_1_1__leaf_net484),
    .X(net490));
 sky130_fd_sc_hd__mux4_2 c634 (.A0(clknet_1_1__leaf_net486),
    .A1(net477),
    .A2(clknet_1_0__leaf_net489),
    .A3(clknet_1_1__leaf_net484),
    .S0(clknet_1_0__leaf_net488),
    .S1(clknet_1_0__leaf_net628),
    .X(net491));
 sky130_fd_sc_hd__mux4_2 c635 (.A0(clknet_1_0__leaf_net490),
    .A1(clknet_1_1__leaf_net489),
    .A2(clknet_1_0__leaf_net491),
    .A3(clknet_1_1__leaf_net483),
    .S0(clknet_1_1__leaf_net487),
    .S1(clknet_1_1__leaf_net628),
    .X(net492));
 sky130_fd_sc_hd__mux4_2 c636 (.A0(clknet_1_0__leaf_net492),
    .A1(clknet_1_0__leaf_net491),
    .A2(clknet_1_1__leaf_net489),
    .A3(clknet_1_1__leaf_net628),
    .S0(net721),
    .S1(clknet_1_1__leaf_net765),
    .X(net493));
 sky130_fd_sc_hd__mux4_2 c637 (.A0(clknet_1_1__leaf_net489),
    .A1(net493),
    .A2(clknet_1_1__leaf_net490),
    .A3(clknet_1_1__leaf_net492),
    .S0(clknet_1_1__leaf_net491),
    .S1(clknet_1_1__leaf_net887),
    .X(net878));
 sky130_fd_sc_hd__a41o_1 c660 (.A1(net904),
    .A2(net385),
    .A3(clknet_1_1__leaf_net402),
    .A4(net286),
    .B1(net923),
    .X(net494));
 sky130_fd_sc_hd__sdfbbn_1 c661 (.CLK_N(clknet_4_5_0_clk),
    .D(net904),
    .RESET_B(net385),
    .SCD(clknet_1_1__leaf_net402),
    .SCE(net626),
    .SET_B(net923),
    .Q(net496),
    .Q_N(net495));
 sky130_fd_sc_hd__a41o_1 c662 (.A1(net496),
    .A2(net385),
    .A3(net904),
    .B1(net923),
    .X(net497));
 sky130_fd_sc_hd__a31o_2 c663 (.A1(net496),
    .A2(net385),
    .A3(net626),
    .B1(net923),
    .X(net498));
 sky130_fd_sc_hd__sdfbbp_1 c664 (.CLK(clknet_4_5_0_clk),
    .D(net496),
    .RESET_B(net498),
    .SCD(net904),
    .SCE(net626),
    .SET_B(net923),
    .Q(net500),
    .Q_N(net499));
 sky130_fd_sc_hd__a41o_1 c665 (.A1(net496),
    .A2(clknet_1_1__leaf_net402),
    .A3(net498),
    .A4(net499),
    .B1(net626),
    .X(net501));
 sky130_fd_sc_hd__mux4_1 c666 (.A0(clknet_1_0__leaf_net501),
    .A1(net495),
    .A2(net386),
    .A3(net499),
    .S0(net498),
    .S1(net626),
    .X(net502));
 sky130_fd_sc_hd__mux4_1 c667 (.A0(clknet_1_0__leaf_net501),
    .A1(clknet_1_1__leaf_net502),
    .A2(net500),
    .A3(net495),
    .S0(net498),
    .S1(net626),
    .X(net503));
 sky130_fd_sc_hd__mux4_1 c668 (.A0(net500),
    .A1(clknet_1_0__leaf_net503),
    .A2(net495),
    .A3(clknet_1_0__leaf_net501),
    .S0(net498),
    .S1(net626),
    .X(net504));
 sky130_fd_sc_hd__mux4_1 c669 (.A0(net498),
    .A1(clknet_1_0__leaf_net501),
    .A2(clknet_1_0__leaf_net502),
    .A3(net495),
    .S0(net499),
    .S1(clknet_1_0__leaf_net503),
    .X(net505));
 sky130_fd_sc_hd__mux4_1 c670 (.A0(clknet_1_0__leaf_net503),
    .A1(clknet_1_1__leaf_net502),
    .A2(clknet_1_1__leaf_net504),
    .A3(clknet_1_0__leaf_net505),
    .S0(net495),
    .S1(clknet_1_0__leaf_net501),
    .X(net506));
 sky130_fd_sc_hd__mux4_1 c671 (.A0(clknet_1_1__leaf_net504),
    .A1(clknet_1_0__leaf_net505),
    .A2(clknet_1_1__leaf_net502),
    .A3(clknet_1_1__leaf_net503),
    .S0(clknet_1_1__leaf_net501),
    .S1(clknet_1_0__leaf_net506),
    .X(net507));
 sky130_fd_sc_hd__mux4_1 c672 (.A0(clknet_1_0__leaf_net507),
    .A1(clknet_1_0__leaf_net506),
    .A2(clknet_1_1__leaf_net504),
    .A3(clknet_1_1__leaf_net501),
    .S0(clknet_1_1__leaf_net503),
    .S1(clknet_1_0__leaf_net505),
    .X(net508));
 sky130_fd_sc_hd__mux4_1 c673 (.A0(net500),
    .A1(clknet_1_0__leaf_net506),
    .A2(clknet_1_1__leaf_net501),
    .A3(clknet_1_0__leaf_net507),
    .S0(clknet_1_0__leaf_net505),
    .S1(clknet_1_1__leaf_net503),
    .X(net509));
 sky130_fd_sc_hd__mux4_1 c674 (.A0(clknet_1_1__leaf_net501),
    .A1(clknet_1_0__leaf_net504),
    .A2(net498),
    .A3(clknet_1_0__leaf_net508),
    .S0(clknet_1_0__leaf_net506),
    .S1(clknet_1_0__leaf_net509),
    .X(net510));
 sky130_fd_sc_hd__mux4_1 c675 (.A0(clknet_1_0__leaf_net503),
    .A1(clknet_1_0__leaf_net504),
    .A2(clknet_1_0__leaf_net509),
    .A3(net496),
    .S0(clknet_1_0__leaf_net506),
    .S1(net626),
    .X(net511));
 sky130_fd_sc_hd__mux4_1 c676 (.A0(clknet_1_0__leaf_net502),
    .A1(clknet_1_0__leaf_net510),
    .A2(clknet_1_0__leaf_net509),
    .A3(clknet_1_0__leaf_net508),
    .S0(clknet_1_1__leaf_net501),
    .S1(clknet_1_0__leaf_net511),
    .X(net512));
 sky130_fd_sc_hd__mux4_1 c677 (.A0(clknet_1_1__leaf_net509),
    .A1(clknet_1_0__leaf_net512),
    .A2(clknet_1_0__leaf_net508),
    .A3(clknet_1_1__leaf_net507),
    .S0(clknet_1_0__leaf_net510),
    .S1(clknet_1_1__leaf_net503),
    .X(net513));
 sky130_fd_sc_hd__mux4_1 c678 (.A0(clknet_1_0__leaf_net513),
    .A1(clknet_1_0__leaf_net512),
    .A2(clknet_1_1__leaf_net511),
    .A3(clknet_1_1__leaf_net510),
    .S0(clknet_1_1__leaf_net507),
    .S1(clknet_1_0__leaf_net505),
    .X(net514));
 sky130_fd_sc_hd__mux4_1 c679 (.A0(net386),
    .A1(net498),
    .A2(clknet_1_1__leaf_net512),
    .A3(clknet_1_0__leaf_net513),
    .S0(clknet_1_0__leaf_net514),
    .S1(clknet_1_1__leaf_net509),
    .X(net515));
 sky130_fd_sc_hd__mux4_1 c680 (.A0(clknet_1_0__leaf_net514),
    .A1(clknet_1_0__leaf_net515),
    .A2(clknet_1_0__leaf_net505),
    .A3(clknet_1_1__leaf_net512),
    .S0(clknet_1_1__leaf_net510),
    .S1(clknet_1_1__leaf_net508),
    .X(net516));
 sky130_fd_sc_hd__mux4_1 c681 (.A0(clknet_1_0__leaf_net511),
    .A1(net516),
    .A2(clknet_1_1__leaf_net514),
    .A3(clknet_1_1__leaf_net515),
    .S0(clknet_1_1__leaf_net513),
    .S1(clknet_1_1__leaf_net512),
    .X(net517));
 sky130_fd_sc_hd__mux4_1 c682 (.A0(clknet_1_1__leaf_net505),
    .A1(net385),
    .A2(clknet_1_1__leaf_net506),
    .A3(clknet_1_1__leaf_net508),
    .S0(net760),
    .S1(net761),
    .X(net518));
 sky130_fd_sc_hd__mux4_1 c683 (.A0(clknet_1_0__leaf_net518),
    .A1(net426),
    .A2(clknet_1_1__leaf_net506),
    .A3(clknet_1_1__leaf_net505),
    .S0(net759),
    .S1(net761),
    .X(net519));
 sky130_fd_sc_hd__mux4_1 c684 (.A0(clknet_1_1__leaf_net518),
    .A1(clknet_1_0__leaf_net519),
    .A2(clknet_1_1__leaf_net506),
    .A3(clknet_1_1__leaf_net505),
    .S0(net759),
    .S1(net761),
    .X(net520));
 sky130_fd_sc_hd__mux4_1 c685 (.A0(clknet_1_1__leaf_net508),
    .A1(clknet_1_0__leaf_net518),
    .A2(clknet_1_0__leaf_net520),
    .A3(clknet_1_0__leaf_net519),
    .S0(clknet_1_0__leaf_net506),
    .S1(clknet_1_1__leaf_net505),
    .X(net521));
 sky130_fd_sc_hd__mux4_1 c686 (.A0(clknet_1_1__leaf_net519),
    .A1(clknet_1_0__leaf_net520),
    .A2(clknet_1_1__leaf_net521),
    .A3(clknet_1_1__leaf_net517),
    .S0(clknet_1_0__leaf_net518),
    .S1(clknet_1_1__leaf_net506),
    .X(net522));
 sky130_fd_sc_hd__mux4_1 c687 (.A0(clknet_1_0__leaf_net518),
    .A1(clknet_1_0__leaf_net520),
    .A2(clknet_1_0__leaf_net522),
    .A3(clknet_1_1__leaf_net521),
    .S0(clknet_1_1__leaf_net519),
    .S1(clknet_1_1__leaf_net505),
    .X(net523));
 sky130_fd_sc_hd__mux4_1 c688 (.A0(clknet_1_0__leaf_net523),
    .A1(clknet_1_1__leaf_net505),
    .A2(clknet_1_0__leaf_net520),
    .A3(clknet_1_1__leaf_net521),
    .S0(clknet_1_0__leaf_net522),
    .S1(clknet_1_1__leaf_net519),
    .X(net524));
 sky130_fd_sc_hd__mux4_1 c689 (.A0(clknet_1_1__leaf_net520),
    .A1(clknet_1_1__leaf_net522),
    .A2(clknet_1_0__leaf_net523),
    .A3(clknet_1_0__leaf_net521),
    .S0(clknet_1_0__leaf_net524),
    .S1(clknet_1_1__leaf_net518),
    .X(net525));
 sky130_fd_sc_hd__mux4_1 c690 (.A0(clknet_1_0__leaf_net524),
    .A1(clknet_1_1__leaf_net525),
    .A2(clknet_1_1__leaf_net521),
    .A3(clknet_1_1__leaf_net518),
    .S0(clknet_1_1__leaf_net520),
    .S1(clknet_1_1__leaf_net522),
    .X(net526));
 sky130_fd_sc_hd__mux4_1 c691 (.A0(clknet_1_1__leaf_net505),
    .A1(clknet_1_0__leaf_net526),
    .A2(clknet_1_1__leaf_net508),
    .A3(clknet_1_0__leaf_net520),
    .S0(clknet_1_1__leaf_net525),
    .S1(clknet_1_1__leaf_net521),
    .X(net527));
 sky130_fd_sc_hd__mux4_1 c692 (.A0(clknet_1_0__leaf_net521),
    .A1(clknet_1_1__leaf_net526),
    .A2(clknet_1_1__leaf_net527),
    .A3(clknet_1_1__leaf_net524),
    .S0(clknet_1_1__leaf_net525),
    .S1(clknet_1_1__leaf_net520),
    .X(net528));
 sky130_fd_sc_hd__mux4_1 c693 (.A0(clknet_1_0__leaf_net527),
    .A1(clknet_1_0__leaf_net521),
    .A2(clknet_1_1__leaf_net525),
    .A3(clknet_1_1__leaf_net520),
    .S0(clknet_1_1__leaf_net522),
    .S1(net703),
    .X(net529));
 sky130_fd_sc_hd__mux4_1 c694 (.A0(clknet_1_0__leaf_net522),
    .A1(clknet_1_0__leaf_net527),
    .A2(clknet_1_0__leaf_net520),
    .A3(clknet_1_1__leaf_net521),
    .S0(clknet_1_1__leaf_net505),
    .S1(clknet_1_0__leaf_net766),
    .X(net530));
 sky130_fd_sc_hd__mux4_1 c695 (.A0(clknet_1_1__leaf_net525),
    .A1(clknet_1_0__leaf_net520),
    .A2(clknet_1_1__leaf_net523),
    .A3(net698),
    .S0(net703),
    .S1(clknet_1_0__leaf_net766),
    .X(net531));
 sky130_fd_sc_hd__mux4_1 c696 (.A0(clknet_1_1__leaf_net526),
    .A1(clknet_1_1__leaf_net523),
    .A2(clknet_1_1__leaf_net525),
    .A3(clknet_1_1__leaf_net520),
    .S0(net698),
    .S1(net703),
    .X(net532));
 sky130_fd_sc_hd__mux4_1 c697 (.A0(clknet_1_1__leaf_net531),
    .A1(clknet_1_1__leaf_net532),
    .A2(clknet_1_1__leaf_net525),
    .A3(clknet_1_1__leaf_net520),
    .S0(net698),
    .S1(clknet_1_1__leaf_net766),
    .X(net533));
 sky130_fd_sc_hd__mux4_1 c698 (.A0(clknet_1_0__leaf_net532),
    .A1(clknet_1_1__leaf_net520),
    .A2(clknet_1_1__leaf_net525),
    .A3(net703),
    .S0(clknet_1_1__leaf_net766),
    .S1(net768),
    .X(net534));
 sky130_fd_sc_hd__mux4_1 c699 (.A0(clknet_1_0__leaf_net526),
    .A1(net426),
    .A2(net690),
    .A3(net698),
    .S0(clknet_1_0__leaf_net766),
    .S1(net767),
    .X(net535));
 sky130_fd_sc_hd__mux4_1 c700 (.A0(clknet_1_0__leaf_net531),
    .A1(clknet_1_0__leaf_net521),
    .A2(clknet_1_0__leaf_net535),
    .A3(clknet_1_1__leaf_net525),
    .S0(net690),
    .S1(net768),
    .X(net536));
 sky130_fd_sc_hd__mux4_1 c701 (.A0(clknet_1_1__leaf_net535),
    .A1(clknet_1_0__leaf_net521),
    .A2(clknet_1_0__leaf_net525),
    .A3(clknet_1_1__leaf_net677),
    .S0(net690),
    .S1(net768),
    .X(net537));
 sky130_fd_sc_hd__mux4_1 c702 (.A0(clknet_1_1__leaf_net506),
    .A1(clknet_1_1__leaf_net535),
    .A2(clknet_1_1__leaf_net677),
    .A3(net703),
    .S0(clknet_1_1__leaf_net766),
    .S1(net768),
    .X(net538));
 sky130_fd_sc_hd__a41o_1 c703 (.A1(clknet_1_0__leaf_net535),
    .A2(clknet_1_0__leaf_net531),
    .A3(clknet_1_1__leaf_net677),
    .A4(net690),
    .B1(net703),
    .X(net539));
 sky130_fd_sc_hd__a41o_1 c704 (.A1(net434),
    .A2(clknet_1_1__leaf_net506),
    .A3(clknet_1_0__leaf_net525),
    .A4(net697),
    .B1(net767),
    .X(net540));
 sky130_fd_sc_hd__a41o_1 c705 (.A1(clknet_1_0__leaf_net540),
    .A2(clknet_1_0__leaf_net525),
    .A3(net434),
    .A4(net697),
    .B1(net767),
    .X(net541));
 sky130_fd_sc_hd__mux4_1 c706 (.A0(clknet_1_0__leaf_net517),
    .A1(clknet_1_0__leaf_net540),
    .A2(net936),
    .A3(clknet_1_0__leaf_net541),
    .S0(clknet_1_0__leaf_net525),
    .S1(net767),
    .X(net542));
 sky130_fd_sc_hd__sdfbbn_2 c707 (.CLK_N(clknet_4_12_0_clk),
    .D(clknet_1_0__leaf_net540),
    .RESET_B(clknet_1_0__leaf_net541),
    .SCD(clknet_1_0__leaf_net525),
    .SCE(net767),
    .SET_B(net769),
    .Q(net544),
    .Q_N(net543));
 sky130_fd_sc_hd__sdfbbn_2 c708 (.CLK_N(clknet_4_13_0_clk),
    .D(net544),
    .RESET_B(clknet_1_1__leaf_net540),
    .SCD(clknet_1_0__leaf_net541),
    .SCE(net697),
    .SET_B(net770),
    .Q(net546),
    .Q_N(net545));
 sky130_fd_sc_hd__mux4_1 c709 (.A0(clknet_1_0__leaf_net525),
    .A1(net544),
    .A2(net546),
    .A3(clknet_1_0__leaf_net540),
    .S0(clknet_1_0__leaf_net541),
    .S1(net769),
    .X(net547));
 sky130_fd_sc_hd__mux4_1 c710 (.A0(net546),
    .A1(clknet_1_1__leaf_net540),
    .A2(net543),
    .A3(clknet_1_0__leaf_net541),
    .S0(net896),
    .S1(net770),
    .X(net548));
 sky130_fd_sc_hd__mux4_1 c711 (.A0(clknet_1_0__leaf_net541),
    .A1(net546),
    .A2(net543),
    .A3(clknet_1_1__leaf_net540),
    .S0(net704),
    .S1(net896),
    .X(net549));
 sky130_fd_sc_hd__mux4_1 c712 (.A0(clknet_1_1__leaf_net540),
    .A1(net543),
    .A2(net545),
    .A3(net704),
    .S0(net896),
    .S1(net772),
    .X(net550));
 sky130_fd_sc_hd__mux4_1 c713 (.A0(clknet_1_0__leaf_net550),
    .A1(clknet_1_0__leaf_net540),
    .A2(net543),
    .A3(net545),
    .S0(net896),
    .S1(net771),
    .X(net551));
 sky130_fd_sc_hd__mux4_1 c714 (.A0(clknet_1_1__leaf_net541),
    .A1(clknet_1_1__leaf_net550),
    .A2(net543),
    .A3(net896),
    .S0(net770),
    .S1(net771),
    .X(net552));
 sky130_fd_sc_hd__mux4_1 c715 (.A0(clknet_1_0__leaf_net550),
    .A1(clknet_1_0__leaf_net540),
    .A2(net543),
    .A3(clknet_1_1__leaf_net675),
    .S0(net769),
    .S1(net771),
    .X(net553));
 sky130_fd_sc_hd__mux4_1 c716 (.A0(net544),
    .A1(clknet_1_1__leaf_net550),
    .A2(net546),
    .A3(clknet_1_1__leaf_net540),
    .S0(clknet_1_1__leaf_net541),
    .S1(net772),
    .X(net554));
 sky130_fd_sc_hd__mux4_1 c717 (.A0(net544),
    .A1(clknet_1_1__leaf_net675),
    .A2(net896),
    .A3(net770),
    .S0(net771),
    .S1(net773),
    .X(net555));
 sky130_fd_sc_hd__mux4_1 c718 (.A0(clknet_1_0__leaf_net555),
    .A1(net543),
    .A2(clknet_1_1__leaf_net675),
    .A3(net702),
    .S0(net771),
    .S1(net773),
    .X(net556));
 sky130_fd_sc_hd__mux4_1 c719 (.A0(clknet_1_1__leaf_net556),
    .A1(clknet_1_1__leaf_net550),
    .A2(net544),
    .A3(net768),
    .S0(net772),
    .S1(net773),
    .X(net557));
 sky130_fd_sc_hd__mux4_1 c720 (.A0(clknet_1_0__leaf_net556),
    .A1(clknet_1_1__leaf_net550),
    .A2(net697),
    .A3(net708),
    .S0(net772),
    .S1(net773),
    .X(net558));
 sky130_fd_sc_hd__mux4_1 c721 (.A0(clknet_1_0__leaf_net556),
    .A1(net691),
    .A2(net702),
    .A3(net704),
    .S0(net708),
    .S1(net773),
    .X(net559));
 sky130_fd_sc_hd__mux4_1 c722 (.A0(clknet_1_0__leaf_net559),
    .A1(net545),
    .A2(net691),
    .A3(net702),
    .S0(net772),
    .S1(net773),
    .X(net560));
 sky130_fd_sc_hd__mux4_1 c723 (.A0(clknet_1_0__leaf_net560),
    .A1(clknet_1_0__leaf_net550),
    .A2(clknet_1_1__leaf_net559),
    .A3(clknet_1_1__leaf_net541),
    .S0(net544),
    .S1(net708),
    .X(net561));
 sky130_fd_sc_hd__mux4_1 c724 (.A0(clknet_1_1__leaf_net555),
    .A1(clknet_1_0__leaf_net559),
    .A2(clknet_1_1__leaf_net560),
    .A3(net544),
    .S0(net691),
    .S1(net708),
    .X(net562));
 sky130_fd_sc_hd__mux4_1 c725 (.A0(clknet_1_1__leaf_net562),
    .A1(clknet_1_1__leaf_net541),
    .A2(clknet_1_0__leaf_net550),
    .A3(net544),
    .S0(net691),
    .S1(net949),
    .X(net563));
 sky130_fd_sc_hd__a41o_1 c726 (.A1(net444),
    .A2(net546),
    .A3(clknet_1_0__leaf_net562),
    .A4(net708),
    .B1(clknet_1_1__leaf_net764),
    .X(net564));
 sky130_fd_sc_hd__a41o_1 c727 (.A1(net546),
    .A2(clknet_1_0__leaf_net564),
    .A3(clknet_1_0__leaf_net525),
    .A4(net708),
    .B1(clknet_1_1__leaf_net764),
    .X(net565));
 sky130_fd_sc_hd__a41o_1 c728 (.A1(clknet_1_0__leaf_net565),
    .A2(clknet_1_0__leaf_net564),
    .A3(net545),
    .A4(net708),
    .B1(clknet_1_1__leaf_net764),
    .X(net566));
 sky130_fd_sc_hd__sdfbbp_1 c729 (.CLK(clknet_4_12_0_clk),
    .D(clknet_1_0__leaf_net565),
    .RESET_B(clknet_1_0__leaf_net564),
    .SCD(clknet_1_0__leaf_net566),
    .SCE(net545),
    .SET_B(clknet_1_0__leaf_net764),
    .Q(net568),
    .Q_N(net567));
 sky130_fd_sc_hd__mux4_1 c730 (.A0(clknet_1_0__leaf_net564),
    .A1(net568),
    .A2(net546),
    .A3(clknet_1_0__leaf_net566),
    .S0(clknet_1_1__leaf_net565),
    .S1(clknet_1_0__leaf_net764),
    .X(net569));
 sky130_fd_sc_hd__mux4_1 c731 (.A0(clknet_1_0__leaf_net566),
    .A1(net567),
    .A2(clknet_1_0__leaf_net565),
    .A3(clknet_1_1__leaf_net564),
    .S0(net545),
    .S1(net774),
    .X(net570));
 sky130_fd_sc_hd__mux4_1 c732 (.A0(net568),
    .A1(clknet_1_0__leaf_net565),
    .A2(clknet_1_1__leaf_net564),
    .A3(net708),
    .S0(net774),
    .S1(net775),
    .X(net571));
 sky130_fd_sc_hd__mux4_1 c733 (.A0(clknet_1_0__leaf_net566),
    .A1(net568),
    .A2(clknet_1_1__leaf_net564),
    .A3(clknet_1_0__leaf_net565),
    .S0(net774),
    .S1(net775),
    .X(net572));
 sky130_fd_sc_hd__mux4_1 c734 (.A0(net568),
    .A1(clknet_1_1__leaf_net564),
    .A2(clknet_1_0__leaf_net565),
    .A3(net774),
    .S0(net775),
    .S1(net776),
    .X(net573));
 sky130_fd_sc_hd__mux4_1 c735 (.A0(clknet_1_1__leaf_net564),
    .A1(clknet_1_1__leaf_net566),
    .A2(clknet_1_0__leaf_net573),
    .A3(net567),
    .S0(net775),
    .S1(net776),
    .X(net574));
 sky130_fd_sc_hd__mux4_1 c736 (.A0(clknet_1_0__leaf_net573),
    .A1(clknet_1_0__leaf_net571),
    .A2(net567),
    .A3(net774),
    .S0(net776),
    .S1(net777),
    .X(net575));
 sky130_fd_sc_hd__mux4_1 c737 (.A0(clknet_1_1__leaf_net573),
    .A1(net685),
    .A2(net774),
    .A3(net775),
    .S0(net776),
    .S1(net777),
    .X(net576));
 sky130_fd_sc_hd__mux4_1 c738 (.A0(clknet_1_1__leaf_net571),
    .A1(net567),
    .A2(net685),
    .A3(net714),
    .S0(net776),
    .S1(net777),
    .X(net577));
 sky130_fd_sc_hd__mux4_1 c739 (.A0(clknet_1_1__leaf_net565),
    .A1(net685),
    .A2(net714),
    .A3(net875),
    .S0(net776),
    .S1(net777),
    .X(net578));
 sky130_fd_sc_hd__mux4_1 c740 (.A0(clknet_1_1__leaf_net573),
    .A1(clknet_1_0__leaf_net578),
    .A2(net875),
    .A3(net774),
    .S0(net775),
    .S1(net777),
    .X(net579));
 sky130_fd_sc_hd__mux4_1 c741 (.A0(clknet_1_1__leaf_net578),
    .A1(net714),
    .A2(net875),
    .A3(net934),
    .S0(net776),
    .S1(net777),
    .X(net580));
 sky130_fd_sc_hd__mux4_1 c742 (.A0(clknet_1_1__leaf_net564),
    .A1(clknet_1_0__leaf_net578),
    .A2(clknet_1_0__leaf_net571),
    .A3(net875),
    .S0(net776),
    .S1(net777),
    .X(net581));
 sky130_fd_sc_hd__mux4_2 c743 (.A0(net685),
    .A1(net691),
    .A2(net714),
    .A3(net934),
    .S0(net776),
    .S1(net777),
    .X(net582));
 sky130_fd_sc_hd__mux4_1 c744 (.A0(net582),
    .A1(clknet_1_1__leaf_net571),
    .A2(net685),
    .A3(net691),
    .S0(net714),
    .S1(net777),
    .X(net583));
 sky130_fd_sc_hd__a41o_1 c745 (.A1(clknet_1_1__leaf_net565),
    .A2(net582),
    .A3(clknet_1_0__leaf_net675),
    .A4(net685),
    .B1(net691),
    .X(net584));
 sky130_fd_sc_hd__mux4_1 c746 (.A0(net582),
    .A1(clknet_1_0__leaf_net584),
    .A2(clknet_1_1__leaf_net573),
    .A3(clknet_1_0__leaf_net675),
    .S0(net685),
    .S1(net875),
    .X(net585));
 sky130_fd_sc_hd__mux4_1 c747 (.A0(clknet_1_1__leaf_net584),
    .A1(net582),
    .A2(clknet_1_0__leaf_net675),
    .A3(net691),
    .S0(net934),
    .S1(net775),
    .X(net586));
 sky130_fd_sc_hd__sdfbbn_2 c748 (.CLK_N(clknet_4_14_0_clk),
    .D(clknet_1_1__leaf_net566),
    .RESET_B(clknet_1_0__leaf_net877),
    .SCD(clknet_1_0__leaf_net878),
    .SCE(clknet_1_0__leaf_net880),
    .SET_B(clknet_1_1__leaf_net884),
    .Q(net588),
    .Q_N(net587));
 sky130_fd_sc_hd__sdfbbn_2 c749 (.CLK_N(clknet_4_14_0_clk),
    .D(net588),
    .RESET_B(clknet_1_1__leaf_net566),
    .SCD(clknet_1_0__leaf_net877),
    .SCE(clknet_1_0__leaf_net880),
    .SET_B(clknet_1_0__leaf_net878),
    .Q(net590),
    .Q_N(net589));
 sky130_fd_sc_hd__mux4_1 c750 (.A0(net588),
    .A1(net590),
    .A2(net879),
    .A3(clknet_1_1__leaf_net566),
    .S0(clknet_1_1__leaf_net880),
    .S1(clknet_1_1__leaf_net877),
    .X(net591));
 sky130_fd_sc_hd__mux4_2 c751 (.A0(net590),
    .A1(clknet_1_0__leaf_net878),
    .A2(net587),
    .A3(clknet_1_1__leaf_net880),
    .S0(net673),
    .S1(net881),
    .X(net592));
 sky130_fd_sc_hd__mux4_2 c752 (.A0(clknet_1_1__leaf_net592),
    .A1(net587),
    .A2(net589),
    .A3(clknet_1_1__leaf_net877),
    .S0(clknet_1_1__leaf_net878),
    .S1(net673),
    .X(net593));
 sky130_fd_sc_hd__a41o_1 c753 (.A1(clknet_1_0__leaf_net593),
    .A2(net590),
    .A3(net587),
    .A4(clknet_1_1__leaf_net592),
    .B1(net673),
    .X(net594));
 sky130_fd_sc_hd__mux4_2 c754 (.A0(clknet_1_0__leaf_net593),
    .A1(clknet_1_1__leaf_net594),
    .A2(clknet_1_1__leaf_net878),
    .A3(net587),
    .S0(net589),
    .S1(net673),
    .X(net595));
 sky130_fd_sc_hd__mux4_2 c755 (.A0(net590),
    .A1(clknet_1_1__leaf_net594),
    .A2(clknet_1_0__leaf_net595),
    .A3(net587),
    .S0(clknet_1_0__leaf_net592),
    .S1(net673),
    .X(net596));
 sky130_fd_sc_hd__mux4_2 c756 (.A0(clknet_1_1__leaf_net596),
    .A1(clknet_1_0__leaf_net595),
    .A2(clknet_1_1__leaf_net594),
    .A3(clknet_1_1__leaf_net880),
    .S0(net587),
    .S1(net589),
    .X(net597));
 sky130_fd_sc_hd__mux4_2 c757 (.A0(clknet_1_1__leaf_net594),
    .A1(clknet_1_1__leaf_net593),
    .A2(clknet_1_0__leaf_net597),
    .A3(net589),
    .S0(clknet_1_0__leaf_net596),
    .S1(clknet_1_0__leaf_net595),
    .X(net598));
 sky130_fd_sc_hd__mux4_2 c758 (.A0(clknet_1_1__leaf_net595),
    .A1(net940),
    .A2(net587),
    .A3(clknet_1_0__leaf_net597),
    .S0(clknet_1_0__leaf_net598),
    .S1(net589),
    .X(net599));
 sky130_fd_sc_hd__mux4_2 c759 (.A0(clknet_1_0__leaf_net599),
    .A1(net588),
    .A2(clknet_1_1__leaf_net595),
    .A3(clknet_1_0__leaf_net594),
    .S0(net590),
    .S1(clknet_1_1__leaf_net598),
    .X(net600));
 sky130_fd_sc_hd__mux4_2 c760 (.A0(clknet_1_1__leaf_net598),
    .A1(clknet_1_0__leaf_net599),
    .A2(clknet_1_1__leaf_net595),
    .A3(net590),
    .S0(net588),
    .S1(clknet_1_0__leaf_net594),
    .X(net888));
 sky130_fd_sc_hd__mux4_2 c761 (.A0(clknet_1_0__leaf_net600),
    .A1(net588),
    .A2(clknet_1_1__leaf_net593),
    .A3(clknet_1_1__leaf_net595),
    .S0(clknet_1_1__leaf_net888),
    .S1(clknet_1_0__leaf_net594),
    .X(net601));
 sky130_fd_sc_hd__mux4_1 c762 (.A0(clknet_1_0__leaf_net601),
    .A1(clknet_1_1__leaf_net599),
    .A2(net589),
    .A3(clknet_1_0__leaf_net595),
    .S0(clknet_1_0__leaf_net600),
    .S1(clknet_1_1__leaf_net594),
    .X(net602));
 sky130_fd_sc_hd__mux4_2 c763 (.A0(clknet_1_0__leaf_net601),
    .A1(clknet_1_1__leaf_net594),
    .A2(clknet_1_1__leaf_net595),
    .A3(clknet_1_1__leaf_net600),
    .S0(clknet_1_1__leaf_net888),
    .S1(net672),
    .X(net603));
 sky130_fd_sc_hd__mux4_2 c764 (.A0(clknet_1_1__leaf_net597),
    .A1(clknet_1_0__leaf_net888),
    .A2(clknet_1_1__leaf_net595),
    .A3(net588),
    .S0(net672),
    .S1(clknet_1_1__leaf_net707),
    .X(net604));
 sky130_fd_sc_hd__mux4_2 c765 (.A0(clknet_1_1__leaf_net599),
    .A1(clknet_1_1__leaf_net604),
    .A2(clknet_1_1__leaf_net601),
    .A3(net590),
    .S0(net672),
    .S1(clknet_1_1__leaf_net707),
    .X(net605));
 sky130_fd_sc_hd__mux4_1 c766 (.A0(clknet_1_0__leaf_net596),
    .A1(clknet_1_0__leaf_net598),
    .A2(net588),
    .A3(clknet_1_0__leaf_net594),
    .S0(clknet_1_0__leaf_net604),
    .S1(clknet_1_0__leaf_net707),
    .X(net606));
 sky130_fd_sc_hd__mux4_1 c767 (.A0(clknet_1_1__leaf_net604),
    .A1(clknet_1_0__leaf_net599),
    .A2(clknet_1_0__leaf_net594),
    .A3(clknet_1_0__leaf_net888),
    .S0(net667),
    .S1(net704),
    .X(net607));
 sky130_fd_sc_hd__mux4_1 c768 (.A0(clknet_1_0__leaf_net604),
    .A1(clknet_1_0__leaf_net592),
    .A2(net667),
    .A3(net672),
    .S1(clknet_1_1__leaf_net884),
    .X(net707));
 sky130_fd_sc_hd__mux4_1 c769 (.A0(clknet_1_1__leaf_net604),
    .A1(net667),
    .A2(net672),
    .A3(clknet_1_0__leaf_net707),
    .S0(net875),
    .S1(clknet_1_1__leaf_net764),
    .X(net609));
 sky130_fd_sc_hd__xnor2_1 merge790 (.A(net552),
    .B(net557),
    .Y(net610));
 sky130_fd_sc_hd__xnor2_1 merge791 (.A(net538),
    .B(net537),
    .Y(net611));
 sky130_fd_sc_hd__dfrbp_2 merge792 (.CLK(clknet_4_4_0_clk),
    .D(net265),
    .Q(net268),
    .Q_N(net612));
 sky130_fd_sc_hd__xnor2_1 merge793 (.A(net585),
    .B(net579),
    .Y(net614));
 sky130_fd_sc_hd__xnor2_1 merge794 (.A(net420),
    .B(net424),
    .Y(net615));
 sky130_fd_sc_hd__xnor2_1 merge795 (.A(net140),
    .B(net141),
    .Y(net616));
 sky130_fd_sc_hd__xnor2_1 merge796 (.A(net377),
    .B(net378),
    .Y(net617));
 sky130_fd_sc_hd__dfrbp_2 merge797 (.CLK(clknet_4_0_0_clk),
    .RESET_B(net80),
    .Q(net619),
    .Q_N(net618));
 sky130_fd_sc_hd__xnor2_1 merge798 (.A(net74),
    .B(net61),
    .Y(net620));
 sky130_fd_sc_hd__xnor2_1 merge799 (.A(net603),
    .B(net605),
    .Y(net621));
 sky130_fd_sc_hd__xnor2_1 merge800 (.A(net466),
    .B(net459),
    .Y(net622));
 sky130_fd_sc_hd__xnor2_1 merge801 (.A(net328),
    .B(net330),
    .Y(net623));
 sky130_fd_sc_hd__xnor2_1 merge802 (.A(net401),
    .B(net391),
    .Y(net624));
 sky130_fd_sc_hd__xnor2_1 merge803 (.A(net111),
    .B(net119),
    .Y(net625));
 sky130_fd_sc_hd__dfrtn_1 merge804 (.CLK_N(clknet_4_10_0_clk),
    .RESET_B(net144),
    .Q(net146));
 sky130_fd_sc_hd__dfrtp_1 merge805 (.CLK(clknet_4_5_0_clk),
    .D(net494),
    .Q(net497));
 sky130_fd_sc_hd__xnor2_1 merge806 (.A(net308),
    .B(net310),
    .Y(net627));
 sky130_fd_sc_hd__dfrtp_4 merge807 (.CLK(clknet_4_11_0_clk),
    .D(net480),
    .Q(net628));
 sky130_fd_sc_hd__xnor2_1 merge808 (.A(net213),
    .B(net214),
    .Y(net629));
 sky130_fd_sc_hd__xnor2_1 merge809 (.A(net29),
    .B(net30),
    .Y(net630));
 sky130_fd_sc_hd__xnor2_1 merge810 (.A(net192),
    .B(net190),
    .Y(net631));
 sky130_fd_sc_hd__dfrtp_1 merge811 (.CLK(clknet_4_8_0_clk),
    .D(net338),
    .Q(net339));
 sky130_fd_sc_hd__xnor2_1 merge812 (.A(net261),
    .B(net260),
    .Y(net633));
 sky130_fd_sc_hd__xnor2_1 merge813 (.A(net167),
    .B(net157),
    .Y(net634));
 sky130_fd_sc_hd__xnor2_1 merge814 (.A(net630),
    .B(net27),
    .Y(net635));
 sky130_fd_sc_hd__dfsbp_1 merge815 (.CLK(clknet_4_8_0_clk),
    .D(net121),
    .SET_B(net28),
    .Q(net637),
    .Q_N(net636));
 sky130_fd_sc_hd__xnor2_1 merge816 (.A(net465),
    .B(net586),
    .Y(net638));
 sky130_fd_sc_hd__dfsbp_1 merge817 (.CLK(clknet_4_2_0_clk),
    .D(net110),
    .SET_B(net112),
    .Q(net640),
    .Q_N(net639));
 sky130_fd_sc_hd__xnor2_1 merge818 (.A(net633),
    .B(net617),
    .Y(net641));
 sky130_fd_sc_hd__dfstp_2 merge819 (.CLK(clknet_4_0_0_clk),
    .D(net64),
    .SET_B(net75),
    .Q(net642));
 sky130_fd_sc_hd__dfstp_2 merge820 (.CLK(clknet_4_1_0_clk),
    .D(net76),
    .SET_B(net70),
    .Q(net643));
 sky130_fd_sc_hd__xnor2_1 merge821 (.A(net215),
    .B(net216),
    .Y(net644));
 sky130_fd_sc_hd__dfstp_1 merge822 (.CLK(clknet_4_2_0_clk),
    .D(net625),
    .Q(net120));
 sky130_fd_sc_hd__xnor2_1 merge823 (.A(net611),
    .B(net398),
    .Y(net646));
 sky130_fd_sc_hd__dlrbn_1 merge824 (.D(net168),
    .GATE_N(clknet_4_4_0_clk),
    .RESET_B(net161),
    .Q(net648),
    .Q_N(net647));
 sky130_fd_sc_hd__dlrbn_1 merge825 (.D(net255),
    .GATE_N(clknet_4_3_0_clk),
    .RESET_B(net203),
    .Q(net650),
    .Q_N(net649));
 sky130_fd_sc_hd__xnor2_1 merge826 (.A(net332),
    .B(net321),
    .Y(net651));
 sky130_fd_sc_hd__xnor2_1 merge827 (.A(net460),
    .B(net461),
    .Y(net652));
 sky130_fd_sc_hd__dlrbp_1 merge828 (.D(net250),
    .GATE(clknet_4_9_0_clk),
    .Q(net654),
    .Q_N(net653));
 sky130_fd_sc_hd__xnor2_1 merge829 (.A(net561),
    .B(net558),
    .Y(net655));
 sky130_fd_sc_hd__xnor2_1 merge830 (.A(net311),
    .B(net326),
    .Y(net656));
 sky130_fd_sc_hd__xnor2_1 merge831 (.A(net372),
    .B(net467),
    .Y(net657));
 sky130_fd_sc_hd__xnor2_1 merge832 (.A(net400),
    .B(net399),
    .Y(net658));
 sky130_fd_sc_hd__xnor2_1 merge833 (.A(net470),
    .B(net623),
    .Y(net659));
 sky130_fd_sc_hd__dlrbp_1 merge834 (.D(net258),
    .GATE(clknet_4_8_0_clk),
    .RESET_B(net26),
    .Q(net661),
    .Q_N(net660));
 sky130_fd_sc_hd__dlrtn_1 merge835 (.D(net415),
    .GATE_N(clknet_4_6_0_clk),
    .RESET_B(net307),
    .Q(net662));
 sky130_fd_sc_hd__xnor2_1 merge836 (.A(net335),
    .B(net333),
    .Y(net663));
 sky130_fd_sc_hd__xnor2_1 merge837 (.A(net331),
    .B(net447),
    .Y(net664));
 sky130_fd_sc_hd__xnor2_1 merge838 (.A(net651),
    .B(net324),
    .Y(net665));
 sky130_fd_sc_hd__xnor2_1 merge839 (.A(net458),
    .B(net374),
    .Y(net666));
 sky130_fd_sc_hd__dlrtn_2 merge840 (.D(net606),
    .GATE_N(clknet_4_14_0_clk),
    .RESET_B(net375),
    .Q(net667));
 sky130_fd_sc_hd__dlrtn_1 merge841 (.D(net624),
    .GATE_N(clknet_4_6_0_clk),
    .RESET_B(net320),
    .Q(net668));
 sky130_fd_sc_hd__dlrtp_2 merge842 (.D(net305),
    .GATE(clknet_4_1_0_clk),
    .RESET_B(net634),
    .Q(net669));
 sky130_fd_sc_hd__dlrtp_2 merge843 (.D(net202),
    .GATE(clknet_4_3_0_clk),
    .RESET_B(net641),
    .Q(net670));
 sky130_fd_sc_hd__dlrtp_2 merge844 (.D(net657),
    .GATE(clknet_4_10_0_clk),
    .RESET_B(net245),
    .Q(net671));
 sky130_fd_sc_hd__edfxbp_1 merge845 (.CLK(clknet_4_15_0_clk),
    .D(net591),
    .DE(net602),
    .Q(net673),
    .Q_N(net672));
 sky130_fd_sc_hd__edfxtp_1 merge846 (.CLK(clknet_4_4_0_clk),
    .D(net153),
    .Q(net154));
 sky130_fd_sc_hd__sdlclkp_1 merge847 (.CLK(clknet_4_13_0_clk),
    .GATE(net551),
    .SCE(net583),
    .GCLK(net675));
 sky130_fd_sc_hd__sdlclkp_2 merge848 (.CLK(clknet_4_8_0_clk),
    .GATE(net253),
    .SCE(net113),
    .GCLK(net676));
 sky130_fd_sc_hd__sdlclkp_4 merge849 (.CLK(clknet_4_13_0_clk),
    .GATE(net658),
    .SCE(net536),
    .GCLK(net677));
 sky130_fd_sc_hd__xnor2_1 merge850 (.A(net469),
    .B(net614),
    .Y(net678));
 sky130_fd_sc_hd__dfrbp_2 merge851 (.CLK(clknet_4_1_0_clk),
    .D(net631),
    .RESET_B(net663),
    .Q(net680),
    .Q_N(net679));
 sky130_fd_sc_hd__dfrbp_2 merge852 (.CLK(clknet_4_2_0_clk),
    .D(net114),
    .RESET_B(net616),
    .Q(net682),
    .Q_N(net681));
 sky130_fd_sc_hd__dfrtn_1 merge853 (.CLK_N(clknet_4_1_0_clk),
    .D(net163),
    .RESET_B(net211),
    .Q(net683));
 sky130_fd_sc_hd__dfrtp_2 merge854 (.CLK(clknet_4_12_0_clk),
    .D(net615),
    .RESET_B(net622),
    .Q(net684));
 sky130_fd_sc_hd__dfrtp_4 merge855 (.CLK(clknet_4_12_0_clk),
    .D(net317),
    .RESET_B(net638),
    .Q(net881));
 sky130_fd_sc_hd__dfrtp_2 merge856 (.CLK(clknet_4_15_0_clk),
    .D(net575),
    .RESET_B(net581),
    .Q(net685));
 sky130_fd_sc_hd__dfsbp_1 merge857 (.CLK(clknet_4_3_0_clk),
    .D(net659),
    .SET_B(net629),
    .Q(net687),
    .Q_N(net686));
 sky130_fd_sc_hd__dfsbp_2 merge858 (.CLK(clknet_4_13_0_clk),
    .D(net387),
    .SET_B(net425),
    .Q(net689),
    .Q_N(net688));
 sky130_fd_sc_hd__dfstp_2 merge859 (.CLK(clknet_4_13_0_clk),
    .D(net300),
    .SET_B(net534),
    .Q(net690));
 sky130_fd_sc_hd__dfstp_2 merge860 (.CLK(clknet_4_15_0_clk),
    .D(net655),
    .SET_B(net580),
    .Q(net691));
 sky130_fd_sc_hd__dfstp_4 merge861 (.CLK(clknet_4_10_0_clk),
    .D(net373),
    .SET_B(net635),
    .Q(net692));
 sky130_fd_sc_hd__dlrbn_1 merge862 (.D(net165),
    .GATE_N(clknet_4_4_0_clk),
    .RESET_B(net58),
    .Q(net694),
    .Q_N(net693));
 sky130_fd_sc_hd__dlrbn_1 merge863 (.D(net198),
    .GATE_N(clknet_4_3_0_clk),
    .RESET_B(net644),
    .Q(net696),
    .Q_N(net695));
 sky130_fd_sc_hd__dlrbp_1 merge864 (.D(net530),
    .GATE(clknet_4_13_0_clk),
    .RESET_B(net539),
    .Q(net698),
    .Q_N(net697));
 sky130_fd_sc_hd__dlrbp_1 merge865 (.D(net656),
    .GATE(clknet_4_6_0_clk),
    .RESET_B(net627),
    .Q(net700),
    .Q_N(net699));
 sky130_fd_sc_hd__dlrtn_4 merge866 (.D(net201),
    .GATE_N(clknet_4_3_0_clk),
    .RESET_B(net664),
    .Q(net701));
 sky130_fd_sc_hd__dlrtn_4 merge867 (.D(net409),
    .GATE_N(clknet_4_13_0_clk),
    .RESET_B(net553),
    .Q(net702));
 sky130_fd_sc_hd__dlrtn_2 merge868 (.D(net528),
    .GATE_N(clknet_4_13_0_clk),
    .RESET_B(net646),
    .Q(net703));
 sky130_fd_sc_hd__dlrtp_2 merge869 (.D(net393),
    .GATE(clknet_4_13_0_clk),
    .RESET_B(net548),
    .Q(net704));
 sky130_fd_sc_hd__dlrtp_2 merge870 (.D(net652),
    .GATE(clknet_4_14_0_clk),
    .RESET_B(net463),
    .Q(net705));
 sky130_fd_sc_hd__dlrtp_4 merge871 (.D(net620),
    .GATE(clknet_4_1_0_clk),
    .RESET_B(net210),
    .Q(net706));
 sky130_fd_sc_hd__edfxbp_1 merge872 (.CLK(clknet_4_15_0_clk),
    .D(net621),
    .Q(net707),
    .Q_N(net876));
 sky130_fd_sc_hd__edfxtp_1 merge873 (.CLK(clknet_4_15_0_clk),
    .D(net563),
    .DE(net610),
    .Q(net708));
 sky130_fd_sc_hd__sdlclkp_1 merge874 (.CLK(clknet_4_1_0_clk),
    .GATE(net176),
    .SCE(net155),
    .GCLK(net709));
 sky130_fd_sc_hd__sdlclkp_2 merge875 (.CLK(clknet_4_4_0_clk),
    .GATE(net162),
    .SCE(net169),
    .GCLK(net710));
 sky130_fd_sc_hd__sdlclkp_4 merge876 (.CLK(clknet_4_2_0_clk),
    .GATE(net252),
    .SCE(net107),
    .GCLK(net711));
 sky130_fd_sc_hd__dfrbp_2 merge877 (.CLK(clknet_4_5_0_clk),
    .D(net296),
    .RESET_B(net408),
    .Q(net713),
    .Q_N(net712));
 sky130_fd_sc_hd__dfrbp_1 merge878 (.CLK(clknet_4_15_0_clk),
    .D(net576),
    .RESET_B(net609),
    .Q(net714),
    .Q_N(net874));
 sky130_fd_sc_hd__dfrtn_1 merge879 (.CLK_N(clknet_4_4_0_clk),
    .D(net59),
    .Q(net62));
 sky130_fd_sc_hd__dfrtp_4 merge880 (.CLK(clknet_4_15_0_clk),
    .D(net607),
    .RESET_B(net577),
    .Q(net875));
 sky130_fd_sc_hd__dfrtp_1 merge881 (.CLK(clknet_4_12_0_clk),
    .D(net318),
    .RESET_B(net678),
    .Q(net716));
 sky130_fd_sc_hd__dfrtp_2 merge882 (.CLK(clknet_4_1_0_clk),
    .D(net150),
    .RESET_B(net666),
    .Q(net717));
 sky130_fd_sc_hd__dfsbp_2 merge883 (.CLK(clknet_4_3_0_clk),
    .D(net665),
    .SET_B(net156),
    .Q(net719),
    .Q_N(net718));
 sky130_fd_sc_hd__dfsbp_2 merge884 (.CLK(clknet_4_11_0_clk),
    .D(net485),
    .SET_B(net464),
    .Q(net721),
    .Q_N(net720));
 sky130_fd_sc_hd__dfstp_4 merge885 (.CLK(clknet_4_14_0_clk),
    .D(net547),
    .SET_B(net262),
    .Q(net896));
 sky130_fd_sc_hd__dfxbp_1 s886 (.CLK(clknet_4_0_0_clk),
    .D(net63),
    .Q(net723),
    .Q_N(net722));
 sky130_fd_sc_hd__dfxbp_1 s887 (.CLK(clknet_4_0_0_clk),
    .D(net68),
    .Q(net725),
    .Q_N(net724));
 sky130_fd_sc_hd__dfxtp_1 s888 (.CLK(clknet_4_0_0_clk),
    .D(net79),
    .Q(net726));
 sky130_fd_sc_hd__dfxtp_1 s889 (.CLK(clknet_4_0_0_clk),
    .D(net82),
    .Q(net727));
 sky130_fd_sc_hd__dfxtp_1 s890 (.CLK(clknet_4_0_0_clk),
    .D(net109),
    .Q(net728));
 sky130_fd_sc_hd__dlclkp_1 s891 (.CLK(clknet_4_2_0_clk),
    .GATE(net115),
    .GCLK(net889));
 sky130_fd_sc_hd__dlclkp_2 s892 (.CLK(clknet_4_2_0_clk),
    .GATE(net118),
    .GCLK(net729));
 sky130_fd_sc_hd__dlclkp_4 s893 (.CLK(clknet_4_10_0_clk),
    .GATE(net145),
    .GCLK(net891));
 sky130_fd_sc_hd__dlxbn_1 s894 (.D(net158),
    .GATE_N(clknet_4_4_0_clk),
    .Q(net731),
    .Q_N(net730));
 sky130_fd_sc_hd__dlxbn_1 s895 (.D(net195),
    .GATE_N(clknet_4_1_0_clk),
    .Q(net733),
    .Q_N(net732));
 sky130_fd_sc_hd__dlxbp_1 s896 (.D(net199),
    .GATE(clknet_4_3_0_clk),
    .Q(net735),
    .Q_N(net734));
 sky130_fd_sc_hd__dlxtn_1 s897 (.D(net200),
    .GATE_N(clknet_4_3_0_clk),
    .Q(net736));
 sky130_fd_sc_hd__dlxtn_1 s898 (.D(net206),
    .GATE_N(clknet_4_2_0_clk),
    .Q(net737));
 sky130_fd_sc_hd__dlxtn_1 s899 (.D(net251),
    .GATE_N(clknet_4_9_0_clk),
    .Q(net897));
 sky130_fd_sc_hd__dlxtp_1 s900 (.D(net257),
    .GATE(clknet_4_9_0_clk),
    .Q(net892));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s901 (.D(net295),
    .SLEEP_B(clknet_4_5_0_clk),
    .Q(net738));
 sky130_fd_sc_hd__dfxbp_1 s902 (.CLK(clknet_4_6_0_clk),
    .D(net297),
    .Q(net740),
    .Q_N(net739));
 sky130_fd_sc_hd__dfxbp_1 s903 (.CLK(clknet_4_4_0_clk),
    .D(net298),
    .Q(net742),
    .Q_N(net741));
 sky130_fd_sc_hd__dfxtp_1 s904 (.CLK(clknet_4_12_0_clk),
    .D(net319),
    .Q(net743));
 sky130_fd_sc_hd__dfxtp_1 s905 (.CLK(clknet_4_3_0_clk),
    .D(net322),
    .Q(net744));
 sky130_fd_sc_hd__dfxtp_2 s906 (.CLK(clknet_4_12_0_clk),
    .D(net323),
    .Q(net745));
 sky130_fd_sc_hd__dlclkp_1 s907 (.CLK(clknet_4_3_0_clk),
    .GATE(net325),
    .GCLK(net746));
 sky130_fd_sc_hd__dlclkp_2 s908 (.CLK(clknet_4_9_0_clk),
    .GATE(net329),
    .GCLK(net747));
 sky130_fd_sc_hd__dlclkp_4 s909 (.CLK(clknet_4_11_0_clk),
    .GATE(net371),
    .GCLK(net884));
 sky130_fd_sc_hd__dlxbn_1 s910 (.D(net379),
    .GATE_N(clknet_4_11_0_clk),
    .Q(net886),
    .Q_N(net885));
 sky130_fd_sc_hd__dlxbn_1 s911 (.D(net390),
    .GATE_N(clknet_4_7_0_clk),
    .Q(net749),
    .Q_N(net748));
 sky130_fd_sc_hd__dlxbp_1 s912 (.D(net392),
    .GATE(clknet_4_7_0_clk),
    .Q(net751),
    .Q_N(net750));
 sky130_fd_sc_hd__dlxtn_2 s913 (.D(net394),
    .GATE_N(clknet_4_7_0_clk),
    .Q(net752));
 sky130_fd_sc_hd__dlxtn_1 s914 (.D(net395),
    .GATE_N(clknet_4_7_0_clk),
    .Q(net753));
 sky130_fd_sc_hd__dlxtn_1 s915 (.D(net403),
    .GATE_N(clknet_4_7_0_clk),
    .Q(net754));
 sky130_fd_sc_hd__dlxtp_1 s916 (.D(net412),
    .GATE(clknet_4_7_0_clk),
    .Q(net755));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s917 (.D(net413),
    .SLEEP_B(clknet_4_6_0_clk),
    .Q(net756));
 sky130_fd_sc_hd__dfxbp_1 s918 (.CLK(clknet_4_7_0_clk),
    .D(net416),
    .Q(net758),
    .Q_N(net757));
 sky130_fd_sc_hd__dfxbp_1 s919 (.CLK(clknet_4_7_0_clk),
    .D(net421),
    .Q(net760),
    .Q_N(net759));
 sky130_fd_sc_hd__dfxtp_1 s920 (.CLK(clknet_4_12_0_clk),
    .D(net422),
    .Q(net761));
 sky130_fd_sc_hd__dfxtp_2 s921 (.CLK(clknet_4_11_0_clk),
    .D(net456),
    .Q(net762));
 sky130_fd_sc_hd__dfxtp_1 s922 (.CLK(clknet_4_11_0_clk),
    .D(net457),
    .Q(net763));
 sky130_fd_sc_hd__dlclkp_1 s923 (.CLK(clknet_4_9_0_clk),
    .GATE(net472),
    .GCLK(net764));
 sky130_fd_sc_hd__dlclkp_2 s924 (.CLK(clknet_4_11_0_clk),
    .GATE(net482),
    .GCLK(net765));
 sky130_fd_sc_hd__dlclkp_4 s925 (.CLK(clknet_4_13_0_clk),
    .GATE(net529),
    .GCLK(net766));
 sky130_fd_sc_hd__dlxbn_1 s926 (.D(net533),
    .GATE_N(clknet_4_13_0_clk),
    .Q(net768),
    .Q_N(net767));
 sky130_fd_sc_hd__dlxbn_1 s927 (.D(net542),
    .GATE_N(clknet_4_12_0_clk),
    .Q(net770),
    .Q_N(net769));
 sky130_fd_sc_hd__dlxbp_1 s928 (.D(net549),
    .GATE(clknet_4_13_0_clk),
    .Q(net772),
    .Q_N(net771));
 sky130_fd_sc_hd__dlxtn_1 s929 (.D(net554),
    .GATE_N(clknet_4_13_0_clk),
    .Q(net773));
 sky130_fd_sc_hd__dlxtn_2 s930 (.D(net569),
    .GATE_N(clknet_4_14_0_clk),
    .Q(net774));
 sky130_fd_sc_hd__dlxtn_2 s931 (.D(net570),
    .GATE_N(clknet_4_14_0_clk),
    .Q(net775));
 sky130_fd_sc_hd__dlxtp_1 s932 (.D(net572),
    .GATE(clknet_4_14_0_clk),
    .Q(net776));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s933 (.D(net574),
    .SLEEP_B(clknet_4_14_0_clk),
    .Q(net777));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Right_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Right_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Right_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Right_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Right_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Right_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Right_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Right_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Right_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Right_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Right_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Right_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Right_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Right_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Right_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Right_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Right_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Right_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Right_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Right_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Right_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_161 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_162 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_163 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_164 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_165 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_166 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_167 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_168 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_169 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_170 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_171 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_172 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_173 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_174 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_175 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_176 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_177 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_178 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_179 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_180 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_181 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_182 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Left_183 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Left_184 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Left_185 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Left_186 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Left_187 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Left_188 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Left_189 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Left_190 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Left_191 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Left_192 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Left_193 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Left_194 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Left_195 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Left_196 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Left_197 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Left_198 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Left_199 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Left_200 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Left_201 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Left_202 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Left_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1347 ();
 sky130_fd_sc_hd__buf_1 input1 (.A(in0),
    .X(net84));
 sky130_fd_sc_hd__buf_1 input2 (.A(in1),
    .X(net254));
 sky130_fd_sc_hd__buf_1 input3 (.A(in10),
    .X(net481));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(in11),
    .X(net608));
 sky130_fd_sc_hd__buf_1 input5 (.A(in12),
    .X(net778));
 sky130_fd_sc_hd__buf_1 input6 (.A(in13),
    .X(net779));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(in14),
    .X(net780));
 sky130_fd_sc_hd__buf_1 input8 (.A(in15),
    .X(net781));
 sky130_fd_sc_hd__buf_1 input9 (.A(in16),
    .X(net782));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(in17),
    .X(net783));
 sky130_fd_sc_hd__buf_1 input11 (.A(in18),
    .X(net784));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(in19),
    .X(net785));
 sky130_fd_sc_hd__buf_1 input13 (.A(in2),
    .X(net786));
 sky130_fd_sc_hd__buf_1 input14 (.A(in20),
    .X(net787));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(in21),
    .X(net788));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(in22),
    .X(net789));
 sky130_fd_sc_hd__buf_1 input17 (.A(in23),
    .X(net790));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(in24),
    .X(net791));
 sky130_fd_sc_hd__clkbuf_1 input19 (.A(in25),
    .X(net792));
 sky130_fd_sc_hd__clkbuf_1 input20 (.A(in26),
    .X(net793));
 sky130_fd_sc_hd__buf_1 input21 (.A(in27),
    .X(net794));
 sky130_fd_sc_hd__buf_1 input22 (.A(in28),
    .X(net795));
 sky130_fd_sc_hd__clkbuf_1 input23 (.A(in29),
    .X(net796));
 sky130_fd_sc_hd__clkbuf_1 input24 (.A(in3),
    .X(net797));
 sky130_fd_sc_hd__clkbuf_1 input25 (.A(in30),
    .X(net798));
 sky130_fd_sc_hd__clkbuf_1 input26 (.A(in31),
    .X(net799));
 sky130_fd_sc_hd__buf_1 input27 (.A(in32),
    .X(net800));
 sky130_fd_sc_hd__clkbuf_1 input28 (.A(in33),
    .X(net801));
 sky130_fd_sc_hd__clkbuf_1 input29 (.A(in34),
    .X(net802));
 sky130_fd_sc_hd__buf_1 input30 (.A(in35),
    .X(net803));
 sky130_fd_sc_hd__buf_1 input31 (.A(in36),
    .X(net804));
 sky130_fd_sc_hd__buf_1 input32 (.A(in37),
    .X(net805));
 sky130_fd_sc_hd__buf_1 input33 (.A(in38),
    .X(net806));
 sky130_fd_sc_hd__buf_1 input34 (.A(in39),
    .X(net807));
 sky130_fd_sc_hd__clkbuf_1 input35 (.A(in4),
    .X(net808));
 sky130_fd_sc_hd__buf_1 input36 (.A(in40),
    .X(net809));
 sky130_fd_sc_hd__clkbuf_1 input37 (.A(in41),
    .X(net810));
 sky130_fd_sc_hd__clkbuf_1 input38 (.A(in42),
    .X(net811));
 sky130_fd_sc_hd__clkbuf_1 input39 (.A(in43),
    .X(net812));
 sky130_fd_sc_hd__buf_1 input40 (.A(in44),
    .X(net813));
 sky130_fd_sc_hd__buf_1 input41 (.A(in45),
    .X(net814));
 sky130_fd_sc_hd__buf_1 input42 (.A(in46),
    .X(net815));
 sky130_fd_sc_hd__dlymetal6s2s_1 input43 (.A(in47),
    .X(net816));
 sky130_fd_sc_hd__clkbuf_1 input44 (.A(in48),
    .X(net817));
 sky130_fd_sc_hd__clkbuf_1 input45 (.A(in49),
    .X(net818));
 sky130_fd_sc_hd__buf_1 input46 (.A(in5),
    .X(net819));
 sky130_fd_sc_hd__buf_1 input47 (.A(in50),
    .X(net820));
 sky130_fd_sc_hd__clkbuf_1 input48 (.A(in51),
    .X(net821));
 sky130_fd_sc_hd__clkbuf_1 input49 (.A(in52),
    .X(net822));
 sky130_fd_sc_hd__clkbuf_1 input50 (.A(in53),
    .X(net823));
 sky130_fd_sc_hd__clkbuf_1 input51 (.A(in54),
    .X(net824));
 sky130_fd_sc_hd__buf_1 input52 (.A(in55),
    .X(net825));
 sky130_fd_sc_hd__buf_1 input53 (.A(in56),
    .X(net826));
 sky130_fd_sc_hd__buf_1 input54 (.A(in57),
    .X(net827));
 sky130_fd_sc_hd__clkbuf_1 input55 (.A(in58),
    .X(net828));
 sky130_fd_sc_hd__clkbuf_1 input56 (.A(in59),
    .X(net829));
 sky130_fd_sc_hd__buf_1 input57 (.A(in6),
    .X(net830));
 sky130_fd_sc_hd__buf_1 input58 (.A(in60),
    .X(net831));
 sky130_fd_sc_hd__buf_1 input59 (.A(in61),
    .X(net832));
 sky130_fd_sc_hd__buf_1 input60 (.A(in62),
    .X(net833));
 sky130_fd_sc_hd__buf_1 input61 (.A(in63),
    .X(net834));
 sky130_fd_sc_hd__buf_1 input62 (.A(in64),
    .X(net835));
 sky130_fd_sc_hd__clkbuf_1 input63 (.A(in65),
    .X(net836));
 sky130_fd_sc_hd__buf_1 input64 (.A(in66),
    .X(net837));
 sky130_fd_sc_hd__clkbuf_1 input65 (.A(in67),
    .X(net838));
 sky130_fd_sc_hd__buf_1 input66 (.A(in68),
    .X(net839));
 sky130_fd_sc_hd__clkbuf_1 input67 (.A(in69),
    .X(net840));
 sky130_fd_sc_hd__clkbuf_1 input68 (.A(in7),
    .X(net841));
 sky130_fd_sc_hd__buf_1 input69 (.A(in70),
    .X(net842));
 sky130_fd_sc_hd__buf_1 input70 (.A(in71),
    .X(net843));
 sky130_fd_sc_hd__clkbuf_1 input71 (.A(in72),
    .X(net844));
 sky130_fd_sc_hd__buf_1 input72 (.A(in73),
    .X(net845));
 sky130_fd_sc_hd__buf_1 input73 (.A(in74),
    .X(net846));
 sky130_fd_sc_hd__buf_1 input74 (.A(in75),
    .X(net847));
 sky130_fd_sc_hd__clkbuf_1 input75 (.A(in76),
    .X(net848));
 sky130_fd_sc_hd__clkbuf_1 input76 (.A(in77),
    .X(net849));
 sky130_fd_sc_hd__clkbuf_1 input77 (.A(in78),
    .X(net850));
 sky130_fd_sc_hd__clkbuf_1 input78 (.A(in79),
    .X(net851));
 sky130_fd_sc_hd__buf_1 input79 (.A(in8),
    .X(net852));
 sky130_fd_sc_hd__clkbuf_1 input80 (.A(in80),
    .X(net853));
 sky130_fd_sc_hd__buf_1 input81 (.A(in81),
    .X(net854));
 sky130_fd_sc_hd__buf_1 input82 (.A(in82),
    .X(net855));
 sky130_fd_sc_hd__clkbuf_1 input83 (.A(in83),
    .X(net856));
 sky130_fd_sc_hd__clkbuf_1 input84 (.A(in84),
    .X(net857));
 sky130_fd_sc_hd__buf_1 input85 (.A(in85),
    .X(net858));
 sky130_fd_sc_hd__clkbuf_1 input86 (.A(in86),
    .X(net859));
 sky130_fd_sc_hd__clkbuf_1 input87 (.A(in87),
    .X(net860));
 sky130_fd_sc_hd__buf_1 input88 (.A(in88),
    .X(net861));
 sky130_fd_sc_hd__buf_1 input89 (.A(in89),
    .X(net862));
 sky130_fd_sc_hd__buf_1 input90 (.A(in9),
    .X(net863));
 sky130_fd_sc_hd__clkbuf_1 input91 (.A(in90),
    .X(net864));
 sky130_fd_sc_hd__clkbuf_2 input92 (.A(in91),
    .X(net865));
 sky130_fd_sc_hd__clkbuf_2 input93 (.A(in92),
    .X(net866));
 sky130_fd_sc_hd__dlymetal6s2s_1 input94 (.A(in93),
    .X(net867));
 sky130_fd_sc_hd__buf_1 input95 (.A(in94),
    .X(net868));
 sky130_fd_sc_hd__clkbuf_1 input96 (.A(in95),
    .X(net869));
 sky130_fd_sc_hd__buf_1 input97 (.A(in96),
    .X(net870));
 sky130_fd_sc_hd__buf_1 input98 (.A(in97),
    .X(net871));
 sky130_fd_sc_hd__clkbuf_1 input99 (.A(in98),
    .X(net872));
 sky130_fd_sc_hd__buf_1 input100 (.A(in99),
    .X(net873));
 sky130_fd_sc_hd__buf_2 output101 (.A(net874),
    .X(out0));
 sky130_fd_sc_hd__buf_2 output102 (.A(net875),
    .X(out15));
 sky130_fd_sc_hd__buf_2 output103 (.A(net876),
    .X(out19));
 sky130_fd_sc_hd__clkbuf_1 output104 (.A(clknet_1_1__leaf_net877),
    .X(out20));
 sky130_fd_sc_hd__clkbuf_1 output105 (.A(clknet_1_1__leaf_net878),
    .X(out22));
 sky130_fd_sc_hd__buf_2 output106 (.A(net879),
    .X(out26));
 sky130_fd_sc_hd__clkbuf_1 output107 (.A(clknet_1_1__leaf_net880),
    .X(out33));
 sky130_fd_sc_hd__buf_2 output108 (.A(net881),
    .X(out4));
 sky130_fd_sc_hd__buf_2 output109 (.A(net882),
    .X(out40));
 sky130_fd_sc_hd__clkbuf_1 output110 (.A(clknet_1_1__leaf_net883),
    .X(out42));
 sky130_fd_sc_hd__clkbuf_1 output111 (.A(clknet_1_0__leaf_net884),
    .X(out47));
 sky130_fd_sc_hd__buf_2 output112 (.A(net885),
    .X(out50));
 sky130_fd_sc_hd__buf_2 output113 (.A(net886),
    .X(out55));
 sky130_fd_sc_hd__clkbuf_1 output114 (.A(clknet_1_1__leaf_net887),
    .X(out58));
 sky130_fd_sc_hd__clkbuf_1 output115 (.A(clknet_1_1__leaf_net888),
    .X(out6));
 sky130_fd_sc_hd__clkbuf_1 output116 (.A(clknet_1_0__leaf_net889),
    .X(out67));
 sky130_fd_sc_hd__clkbuf_1 output117 (.A(clknet_1_1__leaf_net890),
    .X(out68));
 sky130_fd_sc_hd__clkbuf_1 output118 (.A(clknet_1_1__leaf_net891),
    .X(out70));
 sky130_fd_sc_hd__buf_2 output119 (.A(net892),
    .X(out71));
 sky130_fd_sc_hd__buf_2 output120 (.A(net893),
    .X(out72));
 sky130_fd_sc_hd__clkbuf_1 output121 (.A(clknet_1_1__leaf_net894),
    .X(out76));
 sky130_fd_sc_hd__clkbuf_1 output122 (.A(clknet_1_1__leaf_net895),
    .X(out79));
 sky130_fd_sc_hd__buf_2 output123 (.A(net896),
    .X(out81));
 sky130_fd_sc_hd__buf_2 output124 (.A(net897),
    .X(out82));
 sky130_fd_sc_hd__clkbuf_1 output125 (.A(clknet_1_1__leaf_net898),
    .X(out86));
 sky130_fd_sc_hd__buf_2 output126 (.A(net899),
    .X(out87));
 sky130_fd_sc_hd__buf_2 output127 (.A(net900),
    .X(out90));
 sky130_fd_sc_hd__clkbuf_1 output128 (.A(clknet_1_1__leaf_net901),
    .X(out94));
 sky130_fd_sc_hd__clkbuf_2 fanout129 (.A(net196),
    .X(net902));
 sky130_fd_sc_hd__clkbuf_2 fanout130 (.A(net312),
    .X(net903));
 sky130_fd_sc_hd__buf_2 fanout131 (.A(net388),
    .X(net904));
 sky130_fd_sc_hd__buf_2 fanout132 (.A(net383),
    .X(net905));
 sky130_fd_sc_hd__buf_2 fanout133 (.A(net304),
    .X(net906));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout134 (.A(net304),
    .X(net907));
 sky130_fd_sc_hd__buf_2 fanout135 (.A(net73),
    .X(net908));
 sky130_fd_sc_hd__buf_2 fanout136 (.A(net148),
    .X(net909));
 sky130_fd_sc_hd__buf_2 fanout137 (.A(net54),
    .X(net910));
 sky130_fd_sc_hd__buf_2 fanout138 (.A(net147),
    .X(net911));
 sky130_fd_sc_hd__buf_2 fanout139 (.A(net380),
    .X(net912));
 sky130_fd_sc_hd__buf_2 fanout140 (.A(net20),
    .X(net913));
 sky130_fd_sc_hd__buf_2 fanout141 (.A(net11),
    .X(net914));
 sky130_fd_sc_hd__buf_2 fanout142 (.A(net432),
    .X(net915));
 sky130_fd_sc_hd__clkbuf_4 fanout143 (.A(net10),
    .X(net916));
 sky130_fd_sc_hd__buf_2 fanout144 (.A(net35),
    .X(net917));
 sky130_fd_sc_hd__clkbuf_2 fanout145 (.A(net269),
    .X(net918));
 sky130_fd_sc_hd__buf_2 fanout146 (.A(net32),
    .X(net919));
 sky130_fd_sc_hd__buf_2 fanout147 (.A(net763),
    .X(net920));
 sky130_fd_sc_hd__clkbuf_4 fanout148 (.A(net761),
    .X(net921));
 sky130_fd_sc_hd__clkbuf_4 fanout149 (.A(net754),
    .X(net922));
 sky130_fd_sc_hd__clkbuf_4 fanout150 (.A(net753),
    .X(net923));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout151 (.A(net753),
    .X(net924));
 sky130_fd_sc_hd__clkbuf_4 fanout152 (.A(net743),
    .X(net925));
 sky130_fd_sc_hd__clkbuf_2 fanout153 (.A(net743),
    .X(net926));
 sky130_fd_sc_hd__clkbuf_4 fanout154 (.A(net897),
    .X(net927));
 sky130_fd_sc_hd__clkbuf_4 fanout155 (.A(net737),
    .X(net928));
 sky130_fd_sc_hd__clkbuf_4 fanout156 (.A(net736),
    .X(net929));
 sky130_fd_sc_hd__clkbuf_4 fanout157 (.A(net727),
    .X(net930));
 sky130_fd_sc_hd__clkbuf_2 fanout158 (.A(net727),
    .X(net931));
 sky130_fd_sc_hd__clkbuf_4 fanout159 (.A(net726),
    .X(net932));
 sky130_fd_sc_hd__buf_4 fanout160 (.A(net717),
    .X(net933));
 sky130_fd_sc_hd__clkbuf_4 fanout161 (.A(net716),
    .X(net934));
 sky130_fd_sc_hd__buf_2 max_cap162 (.A(net101),
    .X(net935));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net766 (.A(net766),
    .X(clknet_0_net766));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net766 (.A(clknet_0_net766),
    .X(clknet_1_0__leaf_net766));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net766 (.A(clknet_0_net766),
    .X(clknet_1_1__leaf_net766));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net535 (.A(net535),
    .X(clknet_0_net535));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net535 (.A(clknet_0_net535),
    .X(clknet_1_0__leaf_net535));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net535 (.A(clknet_0_net535),
    .X(clknet_1_1__leaf_net535));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net677 (.A(net677),
    .X(clknet_0_net677));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net677 (.A(clknet_0_net677),
    .X(clknet_1_0__leaf_net677));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net677 (.A(clknet_0_net677),
    .X(clknet_1_1__leaf_net677));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net402 (.A(net402),
    .X(clknet_0_net402));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net402 (.A(clknet_0_net402),
    .X(clknet_1_0__leaf_net402));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net402 (.A(clknet_0_net402),
    .X(clknet_1_1__leaf_net402));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net501 (.A(net501),
    .X(clknet_0_net501));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net501 (.A(clknet_0_net501),
    .X(clknet_1_0__leaf_net501));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net501 (.A(clknet_0_net501),
    .X(clknet_1_1__leaf_net501));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net512 (.A(net512),
    .X(clknet_0_net512));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net512 (.A(clknet_0_net512),
    .X(clknet_1_0__leaf_net512));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net512 (.A(clknet_0_net512),
    .X(clknet_1_1__leaf_net512));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net517 (.A(net517),
    .X(clknet_0_net517));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net517 (.A(clknet_0_net517),
    .X(clknet_1_0__leaf_net517));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net517 (.A(clknet_0_net517),
    .X(clknet_1_1__leaf_net517));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net522 (.A(net522),
    .X(clknet_0_net522));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net522 (.A(clknet_0_net522),
    .X(clknet_1_0__leaf_net522));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net522 (.A(clknet_0_net522),
    .X(clknet_1_1__leaf_net522));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net526 (.A(net526),
    .X(clknet_0_net526));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net526 (.A(clknet_0_net526),
    .X(clknet_1_0__leaf_net526));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net526 (.A(clknet_0_net526),
    .X(clknet_1_1__leaf_net526));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net532 (.A(net532),
    .X(clknet_0_net532));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net532 (.A(clknet_0_net532),
    .X(clknet_1_0__leaf_net532));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net532 (.A(clknet_0_net532),
    .X(clknet_1_1__leaf_net532));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net527 (.A(net527),
    .X(clknet_0_net527));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net527 (.A(clknet_0_net527),
    .X(clknet_1_0__leaf_net527));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net527 (.A(clknet_0_net527),
    .X(clknet_1_1__leaf_net527));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net525 (.A(net525),
    .X(clknet_0_net525));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net525 (.A(clknet_0_net525),
    .X(clknet_1_0__leaf_net525));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net525 (.A(clknet_0_net525),
    .X(clknet_1_1__leaf_net525));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net565 (.A(net565),
    .X(clknet_0_net565));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net565 (.A(clknet_0_net565),
    .X(clknet_1_0__leaf_net565));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net565 (.A(clknet_0_net565),
    .X(clknet_1_1__leaf_net565));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net584 (.A(net584),
    .X(clknet_0_net584));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net584 (.A(clknet_0_net584),
    .X(clknet_1_0__leaf_net584));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net584 (.A(clknet_0_net584),
    .X(clknet_1_1__leaf_net584));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net578 (.A(net578),
    .X(clknet_0_net578));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net578 (.A(clknet_0_net578),
    .X(clknet_1_0__leaf_net578));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net578 (.A(clknet_0_net578),
    .X(clknet_1_1__leaf_net578));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net573 (.A(net573),
    .X(clknet_0_net573));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net573 (.A(clknet_0_net573),
    .X(clknet_1_0__leaf_net573));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net573 (.A(clknet_0_net573),
    .X(clknet_1_1__leaf_net573));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net571 (.A(net571),
    .X(clknet_0_net571));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net571 (.A(clknet_0_net571),
    .X(clknet_1_0__leaf_net571));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net571 (.A(clknet_0_net571),
    .X(clknet_1_1__leaf_net571));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net675 (.A(net675),
    .X(clknet_0_net675));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net675 (.A(clknet_0_net675),
    .X(clknet_1_0__leaf_net675));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net675 (.A(clknet_0_net675),
    .X(clknet_1_1__leaf_net675));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net556 (.A(net556),
    .X(clknet_0_net556));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net556 (.A(clknet_0_net556),
    .X(clknet_1_0__leaf_net556));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net556 (.A(clknet_0_net556),
    .X(clknet_1_1__leaf_net556));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net559 (.A(net559),
    .X(clknet_0_net559));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net559 (.A(clknet_0_net559),
    .X(clknet_1_0__leaf_net559));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net559 (.A(clknet_0_net559),
    .X(clknet_1_1__leaf_net559));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net562 (.A(net562),
    .X(clknet_0_net562));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net562 (.A(clknet_0_net562),
    .X(clknet_1_0__leaf_net562));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net562 (.A(clknet_0_net562),
    .X(clknet_1_1__leaf_net562));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net564 (.A(net564),
    .X(clknet_0_net564));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net564 (.A(clknet_0_net564),
    .X(clknet_1_0__leaf_net564));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net564 (.A(clknet_0_net564),
    .X(clknet_1_1__leaf_net564));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net566 (.A(net566),
    .X(clknet_0_net566));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net566 (.A(clknet_0_net566),
    .X(clknet_1_0__leaf_net566));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net566 (.A(clknet_0_net566),
    .X(clknet_1_1__leaf_net566));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net560 (.A(net560),
    .X(clknet_0_net560));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net560 (.A(clknet_0_net560),
    .X(clknet_1_0__leaf_net560));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net560 (.A(clknet_0_net560),
    .X(clknet_1_1__leaf_net560));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net555 (.A(net555),
    .X(clknet_0_net555));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net555 (.A(clknet_0_net555),
    .X(clknet_1_0__leaf_net555));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net555 (.A(clknet_0_net555),
    .X(clknet_1_1__leaf_net555));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net541 (.A(net541),
    .X(clknet_0_net541));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net541 (.A(clknet_0_net541),
    .X(clknet_1_0__leaf_net541));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net541 (.A(clknet_0_net541),
    .X(clknet_1_1__leaf_net541));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net540 (.A(net540),
    .X(clknet_0_net540));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net540 (.A(clknet_0_net540),
    .X(clknet_1_0__leaf_net540));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net540 (.A(clknet_0_net540),
    .X(clknet_1_1__leaf_net540));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net550 (.A(net550),
    .X(clknet_0_net550));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net550 (.A(clknet_0_net550),
    .X(clknet_1_0__leaf_net550));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net550 (.A(clknet_0_net550),
    .X(clknet_1_1__leaf_net550));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net531 (.A(net531),
    .X(clknet_0_net531));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net531 (.A(clknet_0_net531),
    .X(clknet_1_0__leaf_net531));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net531 (.A(clknet_0_net531),
    .X(clknet_1_1__leaf_net531));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net524 (.A(net524),
    .X(clknet_0_net524));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net524 (.A(clknet_0_net524),
    .X(clknet_1_0__leaf_net524));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net524 (.A(clknet_0_net524),
    .X(clknet_1_1__leaf_net524));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net523 (.A(net523),
    .X(clknet_0_net523));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net523 (.A(clknet_0_net523),
    .X(clknet_1_0__leaf_net523));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net523 (.A(clknet_0_net523),
    .X(clknet_1_1__leaf_net523));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net515 (.A(net515),
    .X(clknet_0_net515));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net515 (.A(clknet_0_net515),
    .X(clknet_1_0__leaf_net515));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net515 (.A(clknet_0_net515),
    .X(clknet_1_1__leaf_net515));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net514 (.A(net514),
    .X(clknet_0_net514));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net514 (.A(clknet_0_net514),
    .X(clknet_1_0__leaf_net514));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net514 (.A(clknet_0_net514),
    .X(clknet_1_1__leaf_net514));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net513 (.A(net513),
    .X(clknet_0_net513));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net513 (.A(clknet_0_net513),
    .X(clknet_1_0__leaf_net513));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net513 (.A(clknet_0_net513),
    .X(clknet_1_1__leaf_net513));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net510 (.A(net510),
    .X(clknet_0_net510));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net510 (.A(clknet_0_net510),
    .X(clknet_1_0__leaf_net510));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net510 (.A(clknet_0_net510),
    .X(clknet_1_1__leaf_net510));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net509 (.A(net509),
    .X(clknet_0_net509));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net509 (.A(clknet_0_net509),
    .X(clknet_1_0__leaf_net509));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net509 (.A(clknet_0_net509),
    .X(clknet_1_1__leaf_net509));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net511 (.A(net511),
    .X(clknet_0_net511));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net511 (.A(clknet_0_net511),
    .X(clknet_1_0__leaf_net511));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net511 (.A(clknet_0_net511),
    .X(clknet_1_1__leaf_net511));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net508 (.A(net508),
    .X(clknet_0_net508));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net508 (.A(clknet_0_net508),
    .X(clknet_1_0__leaf_net508));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net508 (.A(clknet_0_net508),
    .X(clknet_1_1__leaf_net508));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net521 (.A(net521),
    .X(clknet_0_net521));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net521 (.A(clknet_0_net521),
    .X(clknet_1_0__leaf_net521));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net521 (.A(clknet_0_net521),
    .X(clknet_1_1__leaf_net521));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net518 (.A(net518),
    .X(clknet_0_net518));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net518 (.A(clknet_0_net518),
    .X(clknet_1_0__leaf_net518));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net518 (.A(clknet_0_net518),
    .X(clknet_1_1__leaf_net518));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net520 (.A(net520),
    .X(clknet_0_net520));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net520 (.A(clknet_0_net520),
    .X(clknet_1_0__leaf_net520));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net520 (.A(clknet_0_net520),
    .X(clknet_1_1__leaf_net520));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net519 (.A(net519),
    .X(clknet_0_net519));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net519 (.A(clknet_0_net519),
    .X(clknet_1_0__leaf_net519));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net519 (.A(clknet_0_net519),
    .X(clknet_1_1__leaf_net519));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net507 (.A(net507),
    .X(clknet_0_net507));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net507 (.A(clknet_0_net507),
    .X(clknet_1_0__leaf_net507));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net507 (.A(clknet_0_net507),
    .X(clknet_1_1__leaf_net507));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net506 (.A(net506),
    .X(clknet_0_net506));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net506 (.A(clknet_0_net506),
    .X(clknet_1_0__leaf_net506));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net506 (.A(clknet_0_net506),
    .X(clknet_1_1__leaf_net506));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net505 (.A(net505),
    .X(clknet_0_net505));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net505 (.A(clknet_0_net505),
    .X(clknet_1_0__leaf_net505));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net505 (.A(clknet_0_net505),
    .X(clknet_1_1__leaf_net505));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net504 (.A(net504),
    .X(clknet_0_net504));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net504 (.A(clknet_0_net504),
    .X(clknet_1_0__leaf_net504));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net504 (.A(clknet_0_net504),
    .X(clknet_1_1__leaf_net504));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net503 (.A(net503),
    .X(clknet_0_net503));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net503 (.A(clknet_0_net503),
    .X(clknet_1_0__leaf_net503));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net503 (.A(clknet_0_net503),
    .X(clknet_1_1__leaf_net503));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net502 (.A(net502),
    .X(clknet_0_net502));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net502 (.A(clknet_0_net502),
    .X(clknet_1_0__leaf_net502));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net502 (.A(clknet_0_net502),
    .X(clknet_1_1__leaf_net502));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net765 (.A(net765),
    .X(clknet_0_net765));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net765 (.A(clknet_0_net765),
    .X(clknet_1_0__leaf_net765));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net765 (.A(clknet_0_net765),
    .X(clknet_1_1__leaf_net765));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net878 (.A(net878),
    .X(clknet_0_net878));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net878 (.A(clknet_0_net878),
    .X(clknet_1_0__leaf_net878));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net878 (.A(clknet_0_net878),
    .X(clknet_1_1__leaf_net878));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net595 (.A(net595),
    .X(clknet_0_net595));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net595 (.A(clknet_0_net595),
    .X(clknet_1_0__leaf_net595));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net595 (.A(clknet_0_net595),
    .X(clknet_1_1__leaf_net595));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net604 (.A(net604),
    .X(clknet_0_net604));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net604 (.A(clknet_0_net604),
    .X(clknet_1_0__leaf_net604));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net604 (.A(clknet_0_net604),
    .X(clknet_1_1__leaf_net604));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net707 (.A(net707),
    .X(clknet_0_net707));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net707 (.A(clknet_0_net707),
    .X(clknet_1_0__leaf_net707));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net707 (.A(clknet_0_net707),
    .X(clknet_1_1__leaf_net707));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net601 (.A(net601),
    .X(clknet_0_net601));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net601 (.A(clknet_0_net601),
    .X(clknet_1_0__leaf_net601));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net601 (.A(clknet_0_net601),
    .X(clknet_1_1__leaf_net601));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net888 (.A(net888),
    .X(clknet_0_net888));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net888 (.A(clknet_0_net888),
    .X(clknet_1_0__leaf_net888));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net888 (.A(clknet_0_net888),
    .X(clknet_1_1__leaf_net888));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net600 (.A(net600),
    .X(clknet_0_net600));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net600 (.A(clknet_0_net600),
    .X(clknet_1_0__leaf_net600));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net600 (.A(clknet_0_net600),
    .X(clknet_1_1__leaf_net600));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net599 (.A(net599),
    .X(clknet_0_net599));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net599 (.A(clknet_0_net599),
    .X(clknet_1_0__leaf_net599));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net599 (.A(clknet_0_net599),
    .X(clknet_1_1__leaf_net599));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net598 (.A(net598),
    .X(clknet_0_net598));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net598 (.A(clknet_0_net598),
    .X(clknet_1_0__leaf_net598));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net598 (.A(clknet_0_net598),
    .X(clknet_1_1__leaf_net598));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net597 (.A(net597),
    .X(clknet_0_net597));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net597 (.A(clknet_0_net597),
    .X(clknet_1_0__leaf_net597));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net597 (.A(net939),
    .X(clknet_1_1__leaf_net597));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net596 (.A(net596),
    .X(clknet_0_net596));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net596 (.A(clknet_0_net596),
    .X(clknet_1_0__leaf_net596));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net596 (.A(clknet_0_net596),
    .X(clknet_1_1__leaf_net596));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net593 (.A(net593),
    .X(clknet_0_net593));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net593 (.A(clknet_0_net593),
    .X(clknet_1_0__leaf_net593));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net593 (.A(clknet_0_net593),
    .X(clknet_1_1__leaf_net593));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net594 (.A(net594),
    .X(clknet_0_net594));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net594 (.A(clknet_0_net594),
    .X(clknet_1_0__leaf_net594));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net594 (.A(clknet_0_net594),
    .X(clknet_1_1__leaf_net594));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net592 (.A(net592),
    .X(clknet_0_net592));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net592 (.A(clknet_0_net592),
    .X(clknet_1_0__leaf_net592));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net592 (.A(clknet_0_net592),
    .X(clknet_1_1__leaf_net592));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net488 (.A(net488),
    .X(clknet_0_net488));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net488 (.A(clknet_0_net488),
    .X(clknet_1_0__leaf_net488));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net488 (.A(clknet_0_net488),
    .X(clknet_1_1__leaf_net488));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net491 (.A(net491),
    .X(clknet_0_net491));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net491 (.A(clknet_0_net491),
    .X(clknet_1_0__leaf_net491));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net491 (.A(clknet_0_net491),
    .X(clknet_1_1__leaf_net491));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net492 (.A(net492),
    .X(clknet_0_net492));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net492 (.A(clknet_0_net492),
    .X(clknet_1_0__leaf_net492));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net492 (.A(clknet_0_net492),
    .X(clknet_1_1__leaf_net492));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net490 (.A(net490),
    .X(clknet_0_net490));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net490 (.A(clknet_0_net490),
    .X(clknet_1_0__leaf_net490));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net490 (.A(clknet_0_net490),
    .X(clknet_1_1__leaf_net490));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net489 (.A(net489),
    .X(clknet_0_net489));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net489 (.A(clknet_0_net489),
    .X(clknet_1_0__leaf_net489));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net489 (.A(clknet_0_net489),
    .X(clknet_1_1__leaf_net489));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net877 (.A(net877),
    .X(clknet_0_net877));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net877 (.A(clknet_0_net877),
    .X(clknet_1_0__leaf_net877));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net877 (.A(clknet_0_net877),
    .X(clknet_1_1__leaf_net877));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net486 (.A(net486),
    .X(clknet_0_net486));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net486 (.A(clknet_0_net486),
    .X(clknet_1_0__leaf_net486));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net486 (.A(clknet_0_net486),
    .X(clknet_1_1__leaf_net486));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net487 (.A(net487),
    .X(clknet_0_net487));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net487 (.A(clknet_0_net487),
    .X(clknet_1_0__leaf_net487));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net487 (.A(clknet_0_net487),
    .X(clknet_1_1__leaf_net487));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net880 (.A(net880),
    .X(clknet_0_net880));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net880 (.A(clknet_0_net880),
    .X(clknet_1_0__leaf_net880));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net880 (.A(clknet_0_net880),
    .X(clknet_1_1__leaf_net880));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net484 (.A(net484),
    .X(clknet_0_net484));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net484 (.A(clknet_0_net484),
    .X(clknet_1_0__leaf_net484));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net484 (.A(clknet_0_net484),
    .X(clknet_1_1__leaf_net484));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net483 (.A(net483),
    .X(clknet_0_net483));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net483 (.A(clknet_0_net483),
    .X(clknet_1_0__leaf_net483));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net483 (.A(clknet_0_net483),
    .X(clknet_1_1__leaf_net483));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net764 (.A(net764),
    .X(clknet_0_net764));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net764 (.A(clknet_0_net764),
    .X(clknet_1_0__leaf_net764));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net764 (.A(clknet_0_net764),
    .X(clknet_1_1__leaf_net764));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net884 (.A(net884),
    .X(clknet_0_net884));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net884 (.A(clknet_0_net884),
    .X(clknet_1_0__leaf_net884));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net884 (.A(clknet_0_net884),
    .X(clknet_1_1__leaf_net884));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net473 (.A(net473),
    .X(clknet_0_net473));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net473 (.A(clknet_0_net473),
    .X(clknet_1_0__leaf_net473));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net473 (.A(clknet_0_net473),
    .X(clknet_1_1__leaf_net473));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net628 (.A(net628),
    .X(clknet_0_net628));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net628 (.A(clknet_0_net628),
    .X(clknet_1_0__leaf_net628));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net628 (.A(clknet_0_net628),
    .X(clknet_1_1__leaf_net628));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net747 (.A(net747),
    .X(clknet_0_net747));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net747 (.A(clknet_0_net747),
    .X(clknet_1_0__leaf_net747));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net747 (.A(clknet_0_net747),
    .X(clknet_1_1__leaf_net747));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net746 (.A(net746),
    .X(clknet_0_net746));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net746 (.A(clknet_0_net746),
    .X(clknet_1_0__leaf_net746));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net746 (.A(clknet_0_net746),
    .X(clknet_1_1__leaf_net746));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net327 (.A(net327),
    .X(clknet_0_net327));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net327 (.A(clknet_0_net327),
    .X(clknet_1_0__leaf_net327));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net327 (.A(clknet_0_net327),
    .X(clknet_1_1__leaf_net327));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net891 (.A(net891),
    .X(clknet_0_net891));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net891 (.A(clknet_0_net891),
    .X(clknet_1_0__leaf_net891));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net891 (.A(clknet_0_net891),
    .X(clknet_1_1__leaf_net891));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net729 (.A(net729),
    .X(clknet_0_net729));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net729 (.A(clknet_0_net729),
    .X(clknet_1_0__leaf_net729));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net729 (.A(clknet_0_net729),
    .X(clknet_1_1__leaf_net729));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net219 (.A(net219),
    .X(clknet_0_net219));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net219 (.A(clknet_0_net219),
    .X(clknet_1_0__leaf_net219));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net219 (.A(clknet_0_net219),
    .X(clknet_1_1__leaf_net219));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net451 (.A(net451),
    .X(clknet_0_net451));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net451 (.A(clknet_0_net451),
    .X(clknet_1_0__leaf_net451));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net451 (.A(clknet_0_net451),
    .X(clknet_1_1__leaf_net451));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net453 (.A(net453),
    .X(clknet_0_net453));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net453 (.A(clknet_0_net453),
    .X(clknet_1_0__leaf_net453));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net453 (.A(clknet_0_net453),
    .X(clknet_1_1__leaf_net453));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net452 (.A(net452),
    .X(clknet_0_net452));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net452 (.A(clknet_0_net452),
    .X(clknet_1_0__leaf_net452));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net452 (.A(clknet_0_net452),
    .X(clknet_1_1__leaf_net452));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net468 (.A(net468),
    .X(clknet_0_net468));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net468 (.A(clknet_0_net468),
    .X(clknet_1_0__leaf_net468));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net468 (.A(clknet_0_net468),
    .X(clknet_1_1__leaf_net468));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net462 (.A(net462),
    .X(clknet_0_net462));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net462 (.A(clknet_0_net462),
    .X(clknet_1_0__leaf_net462));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net462 (.A(clknet_0_net462),
    .X(clknet_1_1__leaf_net462));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net247 (.A(net247),
    .X(clknet_0_net247));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net247 (.A(clknet_0_net247),
    .X(clknet_1_0__leaf_net247));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net247 (.A(clknet_0_net247),
    .X(clknet_1_1__leaf_net247));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net256 (.A(net256),
    .X(clknet_0_net256));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net256 (.A(clknet_0_net256),
    .X(clknet_1_0__leaf_net256));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net256 (.A(clknet_0_net256),
    .X(clknet_1_1__leaf_net256));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net711 (.A(net711),
    .X(clknet_0_net711));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net711 (.A(clknet_0_net711),
    .X(clknet_1_0__leaf_net711));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net711 (.A(clknet_0_net711),
    .X(clknet_1_1__leaf_net711));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net259 (.A(net259),
    .X(clknet_0_net259));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net259 (.A(clknet_0_net259),
    .X(clknet_1_0__leaf_net259));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net259 (.A(clknet_0_net259),
    .X(clknet_1_1__leaf_net259));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net654 (.A(net654),
    .X(clknet_0_net654));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net654 (.A(clknet_0_net654),
    .X(clknet_1_0__leaf_net654));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net654 (.A(clknet_0_net654),
    .X(clknet_1_1__leaf_net654));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net676 (.A(net676),
    .X(clknet_0_net676));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net676 (.A(clknet_0_net676),
    .X(clknet_1_0__leaf_net676));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net676 (.A(clknet_0_net676),
    .X(clknet_1_1__leaf_net676));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net117 (.A(net117),
    .X(clknet_0_net117));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net117 (.A(clknet_0_net117),
    .X(clknet_1_0__leaf_net117));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net117 (.A(clknet_0_net117),
    .X(clknet_1_1__leaf_net117));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net116 (.A(net116),
    .X(clknet_0_net116));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net116 (.A(clknet_0_net116),
    .X(clknet_1_0__leaf_net116));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net116 (.A(clknet_0_net116),
    .X(clknet_1_1__leaf_net116));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net889 (.A(net889),
    .X(clknet_0_net889));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net889 (.A(clknet_0_net889),
    .X(clknet_1_0__leaf_net889));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net889 (.A(clknet_0_net889),
    .X(clknet_1_1__leaf_net889));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net344 (.A(net344),
    .X(clknet_0_net344));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net344 (.A(clknet_0_net344),
    .X(clknet_1_0__leaf_net344));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net344 (.A(clknet_0_net344),
    .X(clknet_1_1__leaf_net344));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net356 (.A(net356),
    .X(clknet_0_net356));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net356 (.A(clknet_0_net356),
    .X(clknet_1_0__leaf_net356));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net356 (.A(clknet_0_net356),
    .X(clknet_1_1__leaf_net356));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net360 (.A(net360),
    .X(clknet_0_net360));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net360 (.A(clknet_0_net360),
    .X(clknet_1_0__leaf_net360));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net360 (.A(clknet_0_net360),
    .X(clknet_1_1__leaf_net360));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net370 (.A(net370),
    .X(clknet_0_net370));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net370 (.A(clknet_0_net370),
    .X(clknet_1_0__leaf_net370));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net370 (.A(clknet_0_net370),
    .X(clknet_1_1__leaf_net370));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net369 (.A(net369),
    .X(clknet_0_net369));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net369 (.A(clknet_0_net369),
    .X(clknet_1_0__leaf_net369));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net369 (.A(clknet_0_net369),
    .X(clknet_1_1__leaf_net369));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net376 (.A(net376),
    .X(clknet_0_net376));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net376 (.A(clknet_0_net376),
    .X(clknet_1_0__leaf_net376));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net376 (.A(clknet_0_net376),
    .X(clknet_1_1__leaf_net376));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net367 (.A(net367),
    .X(clknet_0_net367));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net367 (.A(clknet_0_net367),
    .X(clknet_1_0__leaf_net367));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net367 (.A(clknet_0_net367),
    .X(clknet_1_1__leaf_net367));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net366 (.A(net366),
    .X(clknet_0_net366));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net366 (.A(clknet_0_net366),
    .X(clknet_1_0__leaf_net366));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net366 (.A(clknet_0_net366),
    .X(clknet_1_1__leaf_net366));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net365 (.A(net365),
    .X(clknet_0_net365));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net365 (.A(clknet_0_net365),
    .X(clknet_1_0__leaf_net365));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net365 (.A(clknet_0_net365),
    .X(clknet_1_1__leaf_net365));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net364 (.A(net364),
    .X(clknet_0_net364));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net364 (.A(clknet_0_net364),
    .X(clknet_1_0__leaf_net364));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net364 (.A(clknet_0_net364),
    .X(clknet_1_1__leaf_net364));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net363 (.A(net363),
    .X(clknet_0_net363));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net363 (.A(clknet_0_net363),
    .X(clknet_1_0__leaf_net363));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net363 (.A(clknet_0_net363),
    .X(clknet_1_1__leaf_net363));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net362 (.A(net362),
    .X(clknet_0_net362));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net362 (.A(clknet_0_net362),
    .X(clknet_1_0__leaf_net362));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net362 (.A(clknet_0_net362),
    .X(clknet_1_1__leaf_net362));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net361 (.A(net361),
    .X(clknet_0_net361));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net361 (.A(clknet_0_net361),
    .X(clknet_1_0__leaf_net361));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net361 (.A(clknet_0_net361),
    .X(clknet_1_1__leaf_net361));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net883 (.A(net883),
    .X(clknet_0_net883));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net883 (.A(clknet_0_net883),
    .X(clknet_1_0__leaf_net883));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net883 (.A(clknet_0_net883),
    .X(clknet_1_1__leaf_net883));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net354 (.A(net354),
    .X(clknet_0_net354));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net354 (.A(clknet_0_net354),
    .X(clknet_1_0__leaf_net354));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net354 (.A(clknet_0_net354),
    .X(clknet_1_1__leaf_net354));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net357 (.A(net357),
    .X(clknet_0_net357));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net357 (.A(clknet_0_net357),
    .X(clknet_1_0__leaf_net357));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net357 (.A(clknet_0_net357),
    .X(clknet_1_1__leaf_net357));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net355 (.A(net355),
    .X(clknet_0_net355));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net355 (.A(clknet_0_net355),
    .X(clknet_1_0__leaf_net355));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net355 (.A(clknet_0_net355),
    .X(clknet_1_1__leaf_net355));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net351 (.A(net351),
    .X(clknet_0_net351));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net351 (.A(clknet_0_net351),
    .X(clknet_1_0__leaf_net351));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net351 (.A(clknet_0_net351),
    .X(clknet_1_1__leaf_net351));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net353 (.A(net353),
    .X(clknet_0_net353));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net353 (.A(clknet_0_net353),
    .X(clknet_1_0__leaf_net353));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net353 (.A(clknet_0_net353),
    .X(clknet_1_1__leaf_net353));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net352 (.A(net352),
    .X(clknet_0_net352));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net352 (.A(clknet_0_net352),
    .X(clknet_1_0__leaf_net352));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net352 (.A(clknet_0_net352),
    .X(clknet_1_1__leaf_net352));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net346 (.A(net346),
    .X(clknet_0_net346));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net346 (.A(clknet_0_net346),
    .X(clknet_1_0__leaf_net346));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net346 (.A(clknet_0_net346),
    .X(clknet_1_1__leaf_net346));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net887 (.A(net887),
    .X(clknet_0_net887));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net887 (.A(clknet_0_net887),
    .X(clknet_1_0__leaf_net887));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net887 (.A(clknet_0_net887),
    .X(clknet_1_1__leaf_net887));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net350 (.A(net350),
    .X(clknet_0_net350));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net350 (.A(clknet_0_net350),
    .X(clknet_1_0__leaf_net350));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net350 (.A(clknet_0_net350),
    .X(clknet_1_1__leaf_net350));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net349 (.A(net349),
    .X(clknet_0_net349));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net349 (.A(clknet_0_net349),
    .X(clknet_1_0__leaf_net349));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net349 (.A(clknet_0_net349),
    .X(clknet_1_1__leaf_net349));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net348 (.A(net348),
    .X(clknet_0_net348));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net348 (.A(clknet_0_net348),
    .X(clknet_1_0__leaf_net348));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net348 (.A(clknet_0_net348),
    .X(clknet_1_1__leaf_net348));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net347 (.A(net347),
    .X(clknet_0_net347));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net347 (.A(clknet_0_net347),
    .X(clknet_1_0__leaf_net347));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net347 (.A(clknet_0_net347),
    .X(clknet_1_1__leaf_net347));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net345 (.A(net345),
    .X(clknet_0_net345));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net345 (.A(clknet_0_net345),
    .X(clknet_1_0__leaf_net345));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net345 (.A(clknet_0_net345),
    .X(clknet_1_1__leaf_net345));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net220 (.A(net220),
    .X(clknet_0_net220));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net220 (.A(clknet_0_net220),
    .X(clknet_1_0__leaf_net220));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net220 (.A(clknet_0_net220),
    .X(clknet_1_1__leaf_net220));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net233 (.A(net233),
    .X(clknet_0_net233));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net233 (.A(clknet_0_net233),
    .X(clknet_1_0__leaf_net233));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net233 (.A(clknet_0_net233),
    .X(clknet_1_1__leaf_net233));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net243 (.A(net243),
    .X(clknet_0_net243));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net243 (.A(clknet_0_net243),
    .X(clknet_1_0__leaf_net243));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net243 (.A(clknet_0_net243),
    .X(clknet_1_1__leaf_net243));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net248 (.A(net248),
    .X(clknet_0_net248));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net248 (.A(clknet_0_net248),
    .X(clknet_1_0__leaf_net248));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net248 (.A(clknet_0_net248),
    .X(clknet_1_1__leaf_net248));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net246 (.A(net246),
    .X(clknet_0_net246));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net246 (.A(clknet_0_net246),
    .X(clknet_1_0__leaf_net246));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net246 (.A(clknet_0_net246),
    .X(clknet_1_1__leaf_net246));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net249 (.A(net249),
    .X(clknet_0_net249));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net249 (.A(clknet_0_net249),
    .X(clknet_1_0__leaf_net249));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net249 (.A(clknet_0_net249),
    .X(clknet_1_1__leaf_net249));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net244 (.A(net244),
    .X(clknet_0_net244));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net244 (.A(clknet_0_net244),
    .X(clknet_1_0__leaf_net244));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net244 (.A(clknet_0_net244),
    .X(clknet_1_1__leaf_net244));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net236 (.A(net236),
    .X(clknet_0_net236));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net236 (.A(clknet_0_net236),
    .X(clknet_1_0__leaf_net236));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net236 (.A(clknet_0_net236),
    .X(clknet_1_1__leaf_net236));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net238 (.A(net238),
    .X(clknet_0_net238));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net238 (.A(clknet_0_net238),
    .X(clknet_1_0__leaf_net238));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net238 (.A(clknet_0_net238),
    .X(clknet_1_1__leaf_net238));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net234 (.A(net234),
    .X(clknet_0_net234));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net234 (.A(clknet_0_net234),
    .X(clknet_1_0__leaf_net234));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net234 (.A(clknet_0_net234),
    .X(clknet_1_1__leaf_net234));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net235 (.A(net235),
    .X(clknet_0_net235));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net235 (.A(clknet_0_net235),
    .X(clknet_1_0__leaf_net235));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net235 (.A(clknet_0_net235),
    .X(clknet_1_1__leaf_net235));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net231 (.A(net231),
    .X(clknet_0_net231));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net231 (.A(clknet_0_net231),
    .X(clknet_1_0__leaf_net231));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net231 (.A(clknet_0_net231),
    .X(clknet_1_1__leaf_net231));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net232 (.A(net232),
    .X(clknet_0_net232));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net232 (.A(clknet_0_net232),
    .X(clknet_1_0__leaf_net232));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net232 (.A(clknet_0_net232),
    .X(clknet_1_1__leaf_net232));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net230 (.A(net230),
    .X(clknet_0_net230));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net230 (.A(clknet_0_net230),
    .X(clknet_1_0__leaf_net230));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net230 (.A(clknet_0_net230),
    .X(clknet_1_1__leaf_net230));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net229 (.A(net229),
    .X(clknet_0_net229));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net229 (.A(clknet_0_net229),
    .X(clknet_1_0__leaf_net229));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net229 (.A(clknet_0_net229),
    .X(clknet_1_1__leaf_net229));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net228 (.A(net228),
    .X(clknet_0_net228));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net228 (.A(clknet_0_net228),
    .X(clknet_1_0__leaf_net228));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net228 (.A(clknet_0_net228),
    .X(clknet_1_1__leaf_net228));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net227 (.A(net227),
    .X(clknet_0_net227));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net227 (.A(clknet_0_net227),
    .X(clknet_1_0__leaf_net227));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net227 (.A(clknet_0_net227),
    .X(clknet_1_1__leaf_net227));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net226 (.A(net226),
    .X(clknet_0_net226));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net226 (.A(clknet_0_net226),
    .X(clknet_1_0__leaf_net226));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net226 (.A(clknet_0_net226),
    .X(clknet_1_1__leaf_net226));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net225 (.A(net225),
    .X(clknet_0_net225));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net225 (.A(clknet_0_net225),
    .X(clknet_1_0__leaf_net225));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net225 (.A(clknet_0_net225),
    .X(clknet_1_1__leaf_net225));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net224 (.A(net224),
    .X(clknet_0_net224));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net224 (.A(clknet_0_net224),
    .X(clknet_1_0__leaf_net224));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net224 (.A(clknet_0_net224),
    .X(clknet_1_1__leaf_net224));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net223 (.A(net223),
    .X(clknet_0_net223));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net223 (.A(clknet_0_net223),
    .X(clknet_1_0__leaf_net223));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net223 (.A(clknet_0_net223),
    .X(clknet_1_1__leaf_net223));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net222 (.A(net222),
    .X(clknet_0_net222));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net222 (.A(clknet_0_net222),
    .X(clknet_1_0__leaf_net222));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net222 (.A(clknet_0_net222),
    .X(clknet_1_1__leaf_net222));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net221 (.A(net221),
    .X(clknet_0_net221));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net221 (.A(clknet_0_net221),
    .X(clknet_1_0__leaf_net221));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net221 (.A(clknet_0_net221),
    .X(clknet_1_1__leaf_net221));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net218 (.A(net218),
    .X(clknet_0_net218));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net218 (.A(clknet_0_net218),
    .X(clknet_1_0__leaf_net218));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net218 (.A(clknet_0_net218),
    .X(clknet_1_1__leaf_net218));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net217 (.A(net217),
    .X(clknet_0_net217));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net217 (.A(clknet_0_net217),
    .X(clknet_1_0__leaf_net217));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net217 (.A(clknet_0_net217),
    .X(clknet_1_1__leaf_net217));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net127 (.A(net127),
    .X(clknet_0_net127));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net127 (.A(clknet_0_net127),
    .X(clknet_1_0__leaf_net127));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net127 (.A(clknet_0_net127),
    .X(clknet_1_1__leaf_net127));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net137 (.A(net137),
    .X(clknet_0_net137));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net137 (.A(clknet_0_net137),
    .X(clknet_1_0__leaf_net137));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net137 (.A(clknet_0_net137),
    .X(clknet_1_1__leaf_net137));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net142 (.A(net142),
    .X(clknet_0_net142));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net142 (.A(clknet_0_net142),
    .X(clknet_1_0__leaf_net142));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net142 (.A(clknet_0_net142),
    .X(clknet_1_1__leaf_net142));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net138 (.A(net138),
    .X(clknet_0_net138));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net138 (.A(clknet_0_net138),
    .X(clknet_1_0__leaf_net138));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net138 (.A(clknet_0_net138),
    .X(clknet_1_1__leaf_net138));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net139 (.A(net139),
    .X(clknet_0_net139));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net139 (.A(clknet_0_net139),
    .X(clknet_1_0__leaf_net139));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net139 (.A(clknet_0_net139),
    .X(clknet_1_1__leaf_net139));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net135 (.A(net135),
    .X(clknet_0_net135));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net135 (.A(clknet_0_net135),
    .X(clknet_1_0__leaf_net135));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net135 (.A(clknet_0_net135),
    .X(clknet_1_1__leaf_net135));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net133 (.A(net133),
    .X(clknet_0_net133));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net133 (.A(clknet_0_net133),
    .X(clknet_1_0__leaf_net133));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net133 (.A(clknet_0_net133),
    .X(clknet_1_1__leaf_net133));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net136 (.A(net136),
    .X(clknet_0_net136));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net136 (.A(clknet_0_net136),
    .X(clknet_1_0__leaf_net136));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net136 (.A(clknet_0_net136),
    .X(clknet_1_1__leaf_net136));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net134 (.A(net134),
    .X(clknet_0_net134));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net134 (.A(clknet_0_net134),
    .X(clknet_1_0__leaf_net134));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net134 (.A(clknet_0_net134),
    .X(clknet_1_1__leaf_net134));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net129 (.A(net129),
    .X(clknet_0_net129));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net129 (.A(clknet_0_net129),
    .X(clknet_1_0__leaf_net129));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net129 (.A(clknet_0_net129),
    .X(clknet_1_1__leaf_net129));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net132 (.A(net132),
    .X(clknet_0_net132));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net132 (.A(clknet_0_net132),
    .X(clknet_1_0__leaf_net132));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net132 (.A(clknet_0_net132),
    .X(clknet_1_1__leaf_net132));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net894 (.A(net894),
    .X(clknet_0_net894));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net894 (.A(clknet_0_net894),
    .X(clknet_1_0__leaf_net894));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net894 (.A(clknet_0_net894),
    .X(clknet_1_1__leaf_net894));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net901 (.A(net901),
    .X(clknet_0_net901));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net901 (.A(clknet_0_net901),
    .X(clknet_1_0__leaf_net901));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net901 (.A(clknet_0_net901),
    .X(clknet_1_1__leaf_net901));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net898 (.A(net898),
    .X(clknet_0_net898));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net898 (.A(clknet_0_net898),
    .X(clknet_1_0__leaf_net898));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net898 (.A(clknet_0_net898),
    .X(clknet_1_1__leaf_net898));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net895 (.A(net895),
    .X(clknet_0_net895));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net895 (.A(clknet_0_net895),
    .X(clknet_1_0__leaf_net895));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net895 (.A(clknet_0_net895),
    .X(clknet_1_1__leaf_net895));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net131 (.A(net131),
    .X(clknet_0_net131));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net131 (.A(clknet_0_net131),
    .X(clknet_1_0__leaf_net131));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net131 (.A(clknet_0_net131),
    .X(clknet_1_1__leaf_net131));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net130 (.A(net130),
    .X(clknet_0_net130));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net130 (.A(clknet_0_net130),
    .X(clknet_1_0__leaf_net130));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net130 (.A(clknet_0_net130),
    .X(clknet_1_1__leaf_net130));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net128 (.A(net128),
    .X(clknet_0_net128));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net128 (.A(clknet_0_net128),
    .X(clknet_1_0__leaf_net128));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net128 (.A(clknet_0_net128),
    .X(clknet_1_1__leaf_net128));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net890 (.A(net890),
    .X(clknet_0_net890));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net890 (.A(clknet_0_net890),
    .X(clknet_1_0__leaf_net890));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net890 (.A(clknet_0_net890),
    .X(clknet_1_1__leaf_net890));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net125 (.A(net125),
    .X(clknet_0_net125));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net125 (.A(clknet_0_net125),
    .X(clknet_1_0__leaf_net125));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net125 (.A(clknet_0_net125),
    .X(clknet_1_1__leaf_net125));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net126 (.A(net126),
    .X(clknet_0_net126));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net126 (.A(clknet_0_net126),
    .X(clknet_1_0__leaf_net126));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net126 (.A(clknet_0_net126),
    .X(clknet_1_1__leaf_net126));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net124 (.A(net124),
    .X(clknet_0_net124));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net124 (.A(clknet_0_net124),
    .X(clknet_1_0__leaf_net124));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net124 (.A(clknet_0_net124),
    .X(clknet_1_1__leaf_net124));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net123 (.A(net123),
    .X(clknet_0_net123));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net123 (.A(clknet_0_net123),
    .X(clknet_1_0__leaf_net123));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net123 (.A(clknet_0_net123),
    .X(clknet_1_1__leaf_net123));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net122 (.A(net122),
    .X(clknet_0_net122));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net122 (.A(clknet_0_net122),
    .X(clknet_1_0__leaf_net122));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net122 (.A(clknet_0_net122),
    .X(clknet_1_1__leaf_net122));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net108 (.A(net108),
    .X(clknet_0_net108));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net108 (.A(clknet_0_net108),
    .X(clknet_1_0__leaf_net108));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net108 (.A(clknet_0_net108),
    .X(clknet_1_1__leaf_net108));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net710 (.A(net710),
    .X(clknet_0_net710));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net710 (.A(clknet_0_net710),
    .X(clknet_1_0__leaf_net710));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net710 (.A(clknet_0_net710),
    .X(clknet_1_1__leaf_net710));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net207 (.A(net207),
    .X(clknet_0_net207));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net207 (.A(clknet_0_net207),
    .X(clknet_1_0__leaf_net207));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net207 (.A(clknet_0_net207),
    .X(clknet_1_1__leaf_net207));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net209 (.A(net209),
    .X(clknet_0_net209));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net209 (.A(clknet_0_net209),
    .X(clknet_1_0__leaf_net209));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net209 (.A(clknet_0_net209),
    .X(clknet_1_1__leaf_net209));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net208 (.A(net208),
    .X(clknet_0_net208));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net208 (.A(clknet_0_net208),
    .X(clknet_1_0__leaf_net208));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net208 (.A(clknet_0_net208),
    .X(clknet_1_1__leaf_net208));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net212 (.A(net212),
    .X(clknet_0_net212));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net212 (.A(clknet_0_net212),
    .X(clknet_1_0__leaf_net212));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net212 (.A(clknet_0_net212),
    .X(clknet_1_1__leaf_net212));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net166 (.A(net166),
    .X(clknet_0_net166));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net166 (.A(clknet_0_net166),
    .X(clknet_1_0__leaf_net166));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net166 (.A(clknet_0_net166),
    .X(clknet_1_1__leaf_net166));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net164 (.A(net164),
    .X(clknet_0_net164));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net164 (.A(clknet_0_net164),
    .X(clknet_1_0__leaf_net164));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net164 (.A(clknet_0_net164),
    .X(clknet_1_1__leaf_net164));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net709 (.A(net709),
    .X(clknet_0_net709));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net709 (.A(clknet_0_net709),
    .X(clknet_1_0__leaf_net709));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net709 (.A(clknet_0_net709),
    .X(clknet_1_1__leaf_net709));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net181 (.A(net181),
    .X(clknet_0_net181));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net181 (.A(clknet_0_net181),
    .X(clknet_1_0__leaf_net181));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net181 (.A(clknet_0_net181),
    .X(clknet_1_1__leaf_net181));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net189 (.A(net189),
    .X(clknet_0_net189));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net189 (.A(clknet_0_net189),
    .X(clknet_1_0__leaf_net189));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net189 (.A(clknet_0_net189),
    .X(clknet_1_1__leaf_net189));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net194 (.A(net194),
    .X(clknet_0_net194));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net194 (.A(clknet_0_net194),
    .X(clknet_1_0__leaf_net194));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net194 (.A(clknet_0_net194),
    .X(clknet_1_1__leaf_net194));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net191 (.A(net191),
    .X(clknet_0_net191));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net191 (.A(clknet_0_net191),
    .X(clknet_1_0__leaf_net191));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net191 (.A(clknet_0_net191),
    .X(clknet_1_1__leaf_net191));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net193 (.A(net193),
    .X(clknet_0_net193));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net193 (.A(clknet_0_net193),
    .X(clknet_1_0__leaf_net193));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net193 (.A(clknet_0_net193),
    .X(clknet_1_1__leaf_net193));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net292 (.A(net292),
    .X(clknet_0_net292));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net292 (.A(clknet_0_net292),
    .X(clknet_1_0__leaf_net292));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net292 (.A(clknet_0_net292),
    .X(clknet_1_1__leaf_net292));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net197 (.A(net197),
    .X(clknet_0_net197));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net197 (.A(clknet_0_net197),
    .X(clknet_1_0__leaf_net197));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net197 (.A(clknet_0_net197),
    .X(clknet_1_1__leaf_net197));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net188 (.A(net188),
    .X(clknet_0_net188));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net188 (.A(clknet_0_net188),
    .X(clknet_1_0__leaf_net188));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net188 (.A(clknet_0_net188),
    .X(clknet_1_1__leaf_net188));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net187 (.A(net187),
    .X(clknet_0_net187));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net187 (.A(clknet_0_net187),
    .X(clknet_1_0__leaf_net187));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net187 (.A(clknet_0_net187),
    .X(clknet_1_1__leaf_net187));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net186 (.A(net186),
    .X(clknet_0_net186));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net186 (.A(clknet_0_net186),
    .X(clknet_1_0__leaf_net186));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net186 (.A(clknet_0_net186),
    .X(clknet_1_1__leaf_net186));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net185 (.A(net185),
    .X(clknet_0_net185));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net185 (.A(clknet_0_net185),
    .X(clknet_1_0__leaf_net185));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net185 (.A(clknet_0_net185),
    .X(clknet_1_1__leaf_net185));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net184 (.A(net184),
    .X(clknet_0_net184));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net184 (.A(clknet_0_net184),
    .X(clknet_1_0__leaf_net184));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net184 (.A(clknet_0_net184),
    .X(clknet_1_1__leaf_net184));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net183 (.A(net183),
    .X(clknet_0_net183));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net183 (.A(clknet_0_net183),
    .X(clknet_1_0__leaf_net183));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net183 (.A(clknet_0_net183),
    .X(clknet_1_1__leaf_net183));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net182 (.A(net182),
    .X(clknet_0_net182));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net182 (.A(clknet_0_net182),
    .X(clknet_1_0__leaf_net182));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net182 (.A(clknet_0_net182),
    .X(clknet_1_1__leaf_net182));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net180 (.A(net180),
    .X(clknet_0_net180));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net180 (.A(clknet_0_net180),
    .X(clknet_1_0__leaf_net180));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net180 (.A(clknet_0_net180),
    .X(clknet_1_1__leaf_net180));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net179 (.A(net179),
    .X(clknet_0_net179));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net179 (.A(clknet_0_net179),
    .X(clknet_1_0__leaf_net179));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net179 (.A(clknet_0_net179),
    .X(clknet_1_1__leaf_net179));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net178 (.A(net178),
    .X(clknet_0_net178));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net178 (.A(clknet_0_net178),
    .X(clknet_1_0__leaf_net178));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net178 (.A(clknet_0_net178),
    .X(clknet_1_1__leaf_net178));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net177 (.A(net177),
    .X(clknet_0_net177));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net177 (.A(clknet_0_net177),
    .X(clknet_1_0__leaf_net177));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net177 (.A(clknet_0_net177),
    .X(clknet_1_1__leaf_net177));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net160 (.A(net160),
    .X(clknet_0_net160));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net160 (.A(clknet_0_net160),
    .X(clknet_1_0__leaf_net160));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net160 (.A(clknet_0_net160),
    .X(clknet_1_1__leaf_net160));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net159 (.A(net159),
    .X(clknet_0_net159));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net159 (.A(clknet_0_net159),
    .X(clknet_1_0__leaf_net159));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net159 (.A(clknet_0_net159),
    .X(clknet_1_1__leaf_net159));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer1 (.A(net444),
    .X(net936));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer2 (.A(net410),
    .X(net937));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer3 (.A(net410),
    .X(net938));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer4 (.A(clknet_0_net597),
    .X(net939));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer5 (.A(clknet_1_1__leaf_net594),
    .X(net940));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(net932),
    .X(net941));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(net693),
    .X(net942));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(net643),
    .X(net943));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(net288),
    .X(net944));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(net706),
    .X(net945));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(net723),
    .X(net946));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(net749),
    .X(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_A (.DIODE(clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(in0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(in1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(in10));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(in11));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(in12));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(in13));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(in14));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(in15));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(in16));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(in17));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(in18));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(in19));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(in2));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(in20));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(in21));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(in22));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(in23));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(in24));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(in25));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(in26));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(in27));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_A (.DIODE(in28));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_A (.DIODE(in29));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_A (.DIODE(in3));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_A (.DIODE(in30));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_A (.DIODE(in31));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_A (.DIODE(in32));
 sky130_fd_sc_hd__diode_2 ANTENNA_input28_A (.DIODE(in33));
 sky130_fd_sc_hd__diode_2 ANTENNA_input29_A (.DIODE(in34));
 sky130_fd_sc_hd__diode_2 ANTENNA_input30_A (.DIODE(in35));
 sky130_fd_sc_hd__diode_2 ANTENNA_input31_A (.DIODE(in36));
 sky130_fd_sc_hd__diode_2 ANTENNA_input32_A (.DIODE(in37));
 sky130_fd_sc_hd__diode_2 ANTENNA_input33_A (.DIODE(in38));
 sky130_fd_sc_hd__diode_2 ANTENNA_input34_A (.DIODE(in39));
 sky130_fd_sc_hd__diode_2 ANTENNA_input35_A (.DIODE(in4));
 sky130_fd_sc_hd__diode_2 ANTENNA_input36_A (.DIODE(in40));
 sky130_fd_sc_hd__diode_2 ANTENNA_input37_A (.DIODE(in41));
 sky130_fd_sc_hd__diode_2 ANTENNA_input38_A (.DIODE(in42));
 sky130_fd_sc_hd__diode_2 ANTENNA_input39_A (.DIODE(in43));
 sky130_fd_sc_hd__diode_2 ANTENNA_input40_A (.DIODE(in44));
 sky130_fd_sc_hd__diode_2 ANTENNA_input41_A (.DIODE(in45));
 sky130_fd_sc_hd__diode_2 ANTENNA_input42_A (.DIODE(in46));
 sky130_fd_sc_hd__diode_2 ANTENNA_input43_A (.DIODE(in47));
 sky130_fd_sc_hd__diode_2 ANTENNA_input44_A (.DIODE(in48));
 sky130_fd_sc_hd__diode_2 ANTENNA_input45_A (.DIODE(in49));
 sky130_fd_sc_hd__diode_2 ANTENNA_input46_A (.DIODE(in5));
 sky130_fd_sc_hd__diode_2 ANTENNA_input47_A (.DIODE(in50));
 sky130_fd_sc_hd__diode_2 ANTENNA_input48_A (.DIODE(in51));
 sky130_fd_sc_hd__diode_2 ANTENNA_input49_A (.DIODE(in52));
 sky130_fd_sc_hd__diode_2 ANTENNA_input50_A (.DIODE(in53));
 sky130_fd_sc_hd__diode_2 ANTENNA_input51_A (.DIODE(in54));
 sky130_fd_sc_hd__diode_2 ANTENNA_input52_A (.DIODE(in55));
 sky130_fd_sc_hd__diode_2 ANTENNA_input53_A (.DIODE(in56));
 sky130_fd_sc_hd__diode_2 ANTENNA_input54_A (.DIODE(in57));
 sky130_fd_sc_hd__diode_2 ANTENNA_input55_A (.DIODE(in58));
 sky130_fd_sc_hd__diode_2 ANTENNA_input56_A (.DIODE(in59));
 sky130_fd_sc_hd__diode_2 ANTENNA_input57_A (.DIODE(in6));
 sky130_fd_sc_hd__diode_2 ANTENNA_input58_A (.DIODE(in60));
 sky130_fd_sc_hd__diode_2 ANTENNA_input59_A (.DIODE(in61));
 sky130_fd_sc_hd__diode_2 ANTENNA_input60_A (.DIODE(in62));
 sky130_fd_sc_hd__diode_2 ANTENNA_input61_A (.DIODE(in63));
 sky130_fd_sc_hd__diode_2 ANTENNA_input62_A (.DIODE(in64));
 sky130_fd_sc_hd__diode_2 ANTENNA_input63_A (.DIODE(in65));
 sky130_fd_sc_hd__diode_2 ANTENNA_input64_A (.DIODE(in66));
 sky130_fd_sc_hd__diode_2 ANTENNA_input65_A (.DIODE(in67));
 sky130_fd_sc_hd__diode_2 ANTENNA_input66_A (.DIODE(in68));
 sky130_fd_sc_hd__diode_2 ANTENNA_input67_A (.DIODE(in69));
 sky130_fd_sc_hd__diode_2 ANTENNA_input68_A (.DIODE(in7));
 sky130_fd_sc_hd__diode_2 ANTENNA_input69_A (.DIODE(in70));
 sky130_fd_sc_hd__diode_2 ANTENNA_input70_A (.DIODE(in71));
 sky130_fd_sc_hd__diode_2 ANTENNA_input71_A (.DIODE(in72));
 sky130_fd_sc_hd__diode_2 ANTENNA_input72_A (.DIODE(in73));
 sky130_fd_sc_hd__diode_2 ANTENNA_input73_A (.DIODE(in74));
 sky130_fd_sc_hd__diode_2 ANTENNA_input74_A (.DIODE(in75));
 sky130_fd_sc_hd__diode_2 ANTENNA_input75_A (.DIODE(in76));
 sky130_fd_sc_hd__diode_2 ANTENNA_input76_A (.DIODE(in77));
 sky130_fd_sc_hd__diode_2 ANTENNA_input77_A (.DIODE(in78));
 sky130_fd_sc_hd__diode_2 ANTENNA_input78_A (.DIODE(in79));
 sky130_fd_sc_hd__diode_2 ANTENNA_input79_A (.DIODE(in8));
 sky130_fd_sc_hd__diode_2 ANTENNA_input80_A (.DIODE(in80));
 sky130_fd_sc_hd__diode_2 ANTENNA_input81_A (.DIODE(in81));
 sky130_fd_sc_hd__diode_2 ANTENNA_input82_A (.DIODE(in82));
 sky130_fd_sc_hd__diode_2 ANTENNA_input83_A (.DIODE(in83));
 sky130_fd_sc_hd__diode_2 ANTENNA_input84_A (.DIODE(in84));
 sky130_fd_sc_hd__diode_2 ANTENNA_input85_A (.DIODE(in85));
 sky130_fd_sc_hd__diode_2 ANTENNA_input86_A (.DIODE(in86));
 sky130_fd_sc_hd__diode_2 ANTENNA_input87_A (.DIODE(in87));
 sky130_fd_sc_hd__diode_2 ANTENNA_input88_A (.DIODE(in88));
 sky130_fd_sc_hd__diode_2 ANTENNA_input89_A (.DIODE(in89));
 sky130_fd_sc_hd__diode_2 ANTENNA_input90_A (.DIODE(in9));
 sky130_fd_sc_hd__diode_2 ANTENNA_input91_A (.DIODE(in90));
 sky130_fd_sc_hd__diode_2 ANTENNA_input92_A (.DIODE(in91));
 sky130_fd_sc_hd__diode_2 ANTENNA_input93_A (.DIODE(in92));
 sky130_fd_sc_hd__diode_2 ANTENNA_input94_A (.DIODE(in93));
 sky130_fd_sc_hd__diode_2 ANTENNA_input95_A (.DIODE(in94));
 sky130_fd_sc_hd__diode_2 ANTENNA_input96_A (.DIODE(in95));
 sky130_fd_sc_hd__diode_2 ANTENNA_input97_A (.DIODE(in96));
 sky130_fd_sc_hd__diode_2 ANTENNA_input98_A (.DIODE(in97));
 sky130_fd_sc_hd__diode_2 ANTENNA_input99_A (.DIODE(in98));
 sky130_fd_sc_hd__diode_2 ANTENNA_input100_A (.DIODE(in99));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout143_A (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA_c120_S1 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA_c110_X (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_A0 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_A2 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA_c221_A2 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_A1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_A0 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA_c206_A2 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA_c205_A1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA_c203_A3 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_Q (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA_c125_A3 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_c122_A3 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_c121_S1 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_c120_S0 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_c118_A0 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_c117_A0 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_c116_A3 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_c115_A3 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_c114_X (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge804_RESET_B (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_c261_X (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge804_Q (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_c263_X (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout138_A (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_c273_A2 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_c279_A3 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_c272_A1 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_c264_X (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_c119_A0 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_c118_A1 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_c117_A1 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_c116_S1 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_c115_X (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_c131_A2 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c130_A2 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c124_S0 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c123_S1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c122_A0 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c121_S0 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c120_A2 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c119_A2 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c118_A2 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c117_A3 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c116_X (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c131_A1 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_c125_A0 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_c122_S1 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_c118_A3 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_c117_X (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_B1 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_SCD (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_SCE (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_A3 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_A3 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_S1 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_A2 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_Q_N (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_A3 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA_c321_A0 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_A3 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA_c295_S0 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_A2 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_A3 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_A1 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_A1 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_Q (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA_c127_A3 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_c126_S0 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_c124_S1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_c123_A3 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_c122_A2 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_c121_A0 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_c120_A3 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_c119_A1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_c118_X (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_c128_A3 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c127_S0 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c126_A0 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c125_S0 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c123_A1 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c122_A1 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c121_A2 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c120_A1 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c119_X (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout140_A (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA_c261_S1 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA_c262_A0 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA_c120_X (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA_c129_A1 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_c128_A1 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_c127_A2 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_c125_S1 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_c124_A1 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_c123_A2 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_c121_X (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_A2 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_A2 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA_c532_B1 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA_c531_A4 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA_c530_A4 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA_c528_A3 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_A4 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_SET_B (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA_c398_Q_N (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA_c531_B1 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_c530_A3 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_c529_B1 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_c528_A2 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_SCD (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_A1 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_A1 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_SCE (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_A3 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_c416_S0 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_c415_X (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_A1 (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA_c663_A2 (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA_c662_A2 (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA_c661_RESET_B (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA_c660_A2 (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_A2 (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_RESET_B (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_A3 (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA_c541_A2 (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA_c537_A3 (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA_c533_Q_N (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout131_A (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_S1 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA_c546_A0 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA_c535_X (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA_c528_B1 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_A0 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_SCE (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_c267_B1 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_c266_B1 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_c265_A3 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_c264_B1 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_A2 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_X (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge843_RESET_B (.DIODE(net641));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge818_Y (.DIODE(net641));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge825_Q (.DIODE(net650));
 sky130_fd_sc_hd__diode_2 ANTENNA_c370_A0 (.DIODE(net650));
 sky130_fd_sc_hd__diode_2 ANTENNA_c369_A2 (.DIODE(net650));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_A2 (.DIODE(net650));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_A2 (.DIODE(net650));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge834_Q (.DIODE(net661));
 sky130_fd_sc_hd__diode_2 ANTENNA_c373_A3 (.DIODE(net661));
 sky130_fd_sc_hd__diode_2 ANTENNA_c372_A3 (.DIODE(net661));
 sky130_fd_sc_hd__diode_2 ANTENNA_c371_S0 (.DIODE(net661));
 sky130_fd_sc_hd__diode_2 ANTENNA_c370_A2 (.DIODE(net661));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge882_RESET_B (.DIODE(net666));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge839_Y (.DIODE(net666));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge840_Q (.DIODE(net667));
 sky130_fd_sc_hd__diode_2 ANTENNA_c769_A1 (.DIODE(net667));
 sky130_fd_sc_hd__diode_2 ANTENNA_c768_A2 (.DIODE(net667));
 sky130_fd_sc_hd__diode_2 ANTENNA_c767_S0 (.DIODE(net667));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_A2 (.DIODE(net667));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_A3 (.DIODE(net667));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_S0 (.DIODE(net667));
 sky130_fd_sc_hd__diode_2 ANTENNA_c502_A3 (.DIODE(net667));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge841_Q (.DIODE(net668));
 sky130_fd_sc_hd__diode_2 ANTENNA_c549_A1 (.DIODE(net668));
 sky130_fd_sc_hd__diode_2 ANTENNA_c543_A1 (.DIODE(net668));
 sky130_fd_sc_hd__diode_2 ANTENNA_c540_A3 (.DIODE(net668));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_A1 (.DIODE(net668));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_A2 (.DIODE(net668));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_A3 (.DIODE(net668));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge842_Q (.DIODE(net669));
 sky130_fd_sc_hd__diode_2 ANTENNA_c437_S0 (.DIODE(net669));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_S0 (.DIODE(net669));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_S0 (.DIODE(net669));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_A3 (.DIODE(net669));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_A3 (.DIODE(net669));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_A3 (.DIODE(net669));
 sky130_fd_sc_hd__diode_2 ANTENNA_c274_S0 (.DIODE(net669));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_A0 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_A2 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_A2 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_X (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge843_Q (.DIODE(net670));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_A3 (.DIODE(net670));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_S0 (.DIODE(net670));
 sky130_fd_sc_hd__diode_2 ANTENNA_c373_A4 (.DIODE(net670));
 sky130_fd_sc_hd__diode_2 ANTENNA_c372_S0 (.DIODE(net670));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_A1 (.DIODE(net670));
 sky130_fd_sc_hd__diode_2 ANTENNA_c323_S0 (.DIODE(net670));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_A3 (.DIODE(net670));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_A2 (.DIODE(net670));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge844_Q (.DIODE(net671));
 sky130_fd_sc_hd__diode_2 ANTENNA_c615_A2 (.DIODE(net671));
 sky130_fd_sc_hd__diode_2 ANTENNA_c613_A2 (.DIODE(net671));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_A3 (.DIODE(net671));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_S0 (.DIODE(net671));
 sky130_fd_sc_hd__diode_2 ANTENNA_c373_B1 (.DIODE(net671));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_S0 (.DIODE(net671));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_S1 (.DIODE(net671));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_S1 (.DIODE(net671));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_B1 (.DIODE(net671));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge851_Q_N (.DIODE(net679));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_A4 (.DIODE(net679));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_A3 (.DIODE(net679));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_A3 (.DIODE(net679));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_A1 (.DIODE(net679));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge852_Q_N (.DIODE(net681));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_SET_B (.DIODE(net681));
 sky130_fd_sc_hd__diode_2 ANTENNA_c263_S0 (.DIODE(net681));
 sky130_fd_sc_hd__diode_2 ANTENNA_c256_B1 (.DIODE(net681));
 sky130_fd_sc_hd__diode_2 ANTENNA_c241_B1 (.DIODE(net681));
 sky130_fd_sc_hd__diode_2 ANTENNA_c240_S1 (.DIODE(net681));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge853_Q (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_A2 (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_A2 (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_A2 (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_A2 (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_A4 (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA_c283_A3 (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_A3 (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_S0 (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge854_Q (.DIODE(net684));
 sky130_fd_sc_hd__diode_2 ANTENNA_c611_A2 (.DIODE(net684));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_A2 (.DIODE(net684));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_A3 (.DIODE(net684));
 sky130_fd_sc_hd__diode_2 ANTENNA_c571_A2 (.DIODE(net684));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_A1 (.DIODE(net684));
 sky130_fd_sc_hd__diode_2 ANTENNA_c566_A2 (.DIODE(net684));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge859_Q (.DIODE(net690));
 sky130_fd_sc_hd__diode_2 ANTENNA_c703_A4 (.DIODE(net690));
 sky130_fd_sc_hd__diode_2 ANTENNA_c701_S0 (.DIODE(net690));
 sky130_fd_sc_hd__diode_2 ANTENNA_c700_S0 (.DIODE(net690));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_A2 (.DIODE(net690));
 sky130_fd_sc_hd__diode_2 ANTENNA_c434_S0 (.DIODE(net690));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_S0 (.DIODE(net690));
 sky130_fd_sc_hd__diode_2 ANTENNA_c430_A3 (.DIODE(net690));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_A2 (.DIODE(net690));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge861_Q (.DIODE(net692));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_S0 (.DIODE(net692));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_S1 (.DIODE(net692));
 sky130_fd_sc_hd__diode_2 ANTENNA_c502_S0 (.DIODE(net692));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_S0 (.DIODE(net692));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_S1 (.DIODE(net692));
 sky130_fd_sc_hd__diode_2 ANTENNA_c258_B1 (.DIODE(net692));
 sky130_fd_sc_hd__diode_2 ANTENNA_c131_B1 (.DIODE(net692));
 sky130_fd_sc_hd__diode_2 ANTENNA_c130_S1 (.DIODE(net692));
 sky130_fd_sc_hd__diode_2 ANTENNA_c129_S1 (.DIODE(net692));
 sky130_fd_sc_hd__diode_2 ANTENNA_c128_S1 (.DIODE(net692));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge862_Q (.DIODE(net694));
 sky130_fd_sc_hd__diode_2 ANTENNA_c397_A4 (.DIODE(net694));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_RESET_B (.DIODE(net694));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_SCE (.DIODE(net694));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_B1 (.DIODE(net694));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_SCD (.DIODE(net694));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge866_Q (.DIODE(net701));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_B1 (.DIODE(net701));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_SET_B (.DIODE(net701));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_S1 (.DIODE(net701));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_A2 (.DIODE(net701));
 sky130_fd_sc_hd__diode_2 ANTENNA_c458_A3 (.DIODE(net701));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_A3 (.DIODE(net701));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_A3 (.DIODE(net701));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_A3 (.DIODE(net701));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_A2 (.DIODE(net701));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_S0 (.DIODE(net701));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge867_Q (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_S1 (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_A3 (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_A2 (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_A3 (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c566_A3 (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c561_A3 (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c557_S0 (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c555_A3 (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge869_Q (.DIODE(net704));
 sky130_fd_sc_hd__diode_2 ANTENNA_c767_S1 (.DIODE(net704));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_A3 (.DIODE(net704));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_A3 (.DIODE(net704));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_S0 (.DIODE(net704));
 sky130_fd_sc_hd__diode_2 ANTENNA_c546_A3 (.DIODE(net704));
 sky130_fd_sc_hd__diode_2 ANTENNA_c544_A2 (.DIODE(net704));
 sky130_fd_sc_hd__diode_2 ANTENNA_c542_A3 (.DIODE(net704));
 sky130_fd_sc_hd__diode_2 ANTENNA_c541_A3 (.DIODE(net704));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold10_A (.DIODE(net706));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge871_Q (.DIODE(net706));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_S0 (.DIODE(net706));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_S0 (.DIODE(net706));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_A3 (.DIODE(net706));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_S0 (.DIODE(net706));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_S1 (.DIODE(net706));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_SET_B (.DIODE(net706));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_S1 (.DIODE(net706));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_S0 (.DIODE(net706));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_S0 (.DIODE(net706));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout160_A (.DIODE(net717));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_A3 (.DIODE(net717));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge882_Q (.DIODE(net717));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge883_Q (.DIODE(net719));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_A2 (.DIODE(net719));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_S1 (.DIODE(net719));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_A4 (.DIODE(net719));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_A2 (.DIODE(net719));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_A3 (.DIODE(net719));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_S0 (.DIODE(net719));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout135_A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_SCE (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_c183_A3 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_A0 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_S0 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_X (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout155_A (.DIODE(net737));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_S1 (.DIODE(net737));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_B1 (.DIODE(net737));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_B1 (.DIODE(net737));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_SCE (.DIODE(net737));
 sky130_fd_sc_hd__diode_2 ANTENNA_s898_Q (.DIODE(net737));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_A2 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_A3 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_c321_A2 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_A1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_c311_S0 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_A3 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_A1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_A0 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_A1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_X (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_X (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_A0 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_A3 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_X (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_A3 (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_S0 (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_input33_X (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_RESET_B (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA_input40_X (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_A2 (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_A0 (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_input43_X (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_A0 (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_A3 (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_input60_X (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_c194_A3 (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_A3 (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_input81_X (.DIODE(net854));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_S0 (.DIODE(net854));
 sky130_fd_sc_hd__diode_2 ANTENNA_c102_A3 (.DIODE(net854));
 sky130_fd_sc_hd__diode_2 ANTENNA_output102_A (.DIODE(net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge880_Q (.DIODE(net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_c769_S0 (.DIODE(net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_c746_S1 (.DIODE(net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_c742_A3 (.DIODE(net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_A2 (.DIODE(net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_A2 (.DIODE(net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_c739_A3 (.DIODE(net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_output108_A (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge855_Q (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_S1 (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c610_A3 (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_A2 (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_S0 (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c446_A3 (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_A3 (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_A4 (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net891_A (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_s893_GCLK (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_output119_A (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_s900_Q (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_A3 (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_S1 (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_S1 (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_c372_S1 (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_c371_S1 (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_c370_S1 (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_c369_B1 (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net894_A (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c259_X (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net895_A (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_c256_X (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_output123_A (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge885_Q (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_A2 (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_A3 (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_S0 (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_S0 (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_S1 (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_S0 (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_SCE (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_A4 (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout154_A (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_output124_A (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_s899_Q (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net898_A (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c258_X (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net901_A (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_c260_X (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout133_X (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_A0 (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_c564_A3 (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_A2 (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_A2 (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_A1 (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_c434_A1 (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_A0 (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_D (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_A1 (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_A1 (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout135_X (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_A3 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_A2 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_S0 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_SCE (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_A4 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_RESET_B (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_A0 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_A3 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_A1 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c286_SCD (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout138_X (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_c267_A1 (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_c276_A1 (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_c275_A0 (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_c271_A2 (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_c265_A1 (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_c266_A2 (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_c270_A0 (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_c269_A2 (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_RESET_B (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_c274_A1 (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout140_X (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA_c260_B1 (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA_c259_A4 (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA_c258_A4 (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA_c257_SCD (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA_c256_A2 (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA_c130_A0 (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA_c126_A1 (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA_c123_S0 (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA_c122_S0 (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA_c121_A1 (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout141_X (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA_c131_A3 (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA_c124_A3 (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA_c119_S0 (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA_c117_A2 (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA_c116_A1 (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA_c115_A4 (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA_c114_A3 (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA_c113_A2 (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA_c112_A1 (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA_c118_S1 (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout143_X (.DIODE(net916));
 sky130_fd_sc_hd__diode_2 ANTENNA_c116_A0 (.DIODE(net916));
 sky130_fd_sc_hd__diode_2 ANTENNA_c115_A2 (.DIODE(net916));
 sky130_fd_sc_hd__diode_2 ANTENNA_c129_A0 (.DIODE(net916));
 sky130_fd_sc_hd__diode_2 ANTENNA_c119_S1 (.DIODE(net916));
 sky130_fd_sc_hd__diode_2 ANTENNA_c118_S0 (.DIODE(net916));
 sky130_fd_sc_hd__diode_2 ANTENNA_c117_S0 (.DIODE(net916));
 sky130_fd_sc_hd__diode_2 ANTENNA_c114_B1 (.DIODE(net916));
 sky130_fd_sc_hd__diode_2 ANTENNA_c113_A1 (.DIODE(net916));
 sky130_fd_sc_hd__diode_2 ANTENNA_c112_A2 (.DIODE(net916));
 sky130_fd_sc_hd__diode_2 ANTENNA_c111_A1 (.DIODE(net916));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout148_X (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_S1 (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_c571_B1 (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_S1 (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_B1 (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_B1 (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_B1 (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_B1 (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_B1 (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_S1 (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_B1 (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout150_X (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_A4 (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c660_B1 (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c664_SET_B (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c663_B1 (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c662_B1 (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c661_SET_B (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_SCE (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_SCE (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_S0 (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_S1 (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout152_X (.DIODE(net925));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_A3 (.DIODE(net925));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_S0 (.DIODE(net925));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_S0 (.DIODE(net925));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_A3 (.DIODE(net925));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_S1 (.DIODE(net925));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_S0 (.DIODE(net925));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_SET_B (.DIODE(net925));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_SCE (.DIODE(net925));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_B1 (.DIODE(net925));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_B1 (.DIODE(net925));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout154_X (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_RESET_B (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_S0 (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_S1 (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_S0 (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_B1 (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_SET_B (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_B1 (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c369_A4 (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c365_S1 (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_S1 (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout155_X (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_SET_B (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_B1 (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_S1 (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c321_S1 (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_S1 (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_S1 (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_S1 (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_B1 (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_S1 (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_S1 (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout157_X (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_S1 (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_c190_S1 (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_S1 (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_S1 (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_c184_S1 (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_c182_S1 (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_S0 (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_S0 (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_c203_S1 (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_S1 (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout160_X (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_S0 (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_A3 (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_S1 (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c502_S1 (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_S1 (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_S0 (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c273_S1 (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c270_S1 (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c269_B1 (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_SET_B (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout161_X (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c613_A3 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c743_A3 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_A3 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c747_S0 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_A2 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_A2 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_A3 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_A3 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c446_S0 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_S0 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap162_X (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_SCD (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_S0 (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c220_A2 (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_A4 (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_A1 (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_S0 (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_15_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_14_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_13_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_12_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_11_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_10_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_9_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_8_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_7_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_6_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_5_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_4_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_3_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_2_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_1_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_0_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_X (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_CLK_N (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge797_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge819_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s886_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s887_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s888_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s889_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s890_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_0_0_clk_X (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_CLK_N (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_CLK_N (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c286_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_CLK_N (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge820_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge842_GATE (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge851_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge853_CLK_N (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge871_GATE (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge874_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge882_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s895_GATE_N (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_1_0_clk_X (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge817_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge822_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge852_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge876_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s891_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s892_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s898_GATE_N (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_2_0_clk_X (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_CLK_N (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge825_GATE_N (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge843_GATE (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge857_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge863_GATE_N (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge866_GATE_N (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge883_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s896_GATE (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s897_GATE_N (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s905_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s907_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_3_0_clk_X (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_CLK_N (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_CLK_N (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c398_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_CLK_N (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge792_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge824_GATE_N (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge846_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge862_GATE_N (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge875_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge879_CLK_N (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s894_GATE_N (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s903_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_4_0_clk_X (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge835_GATE_N (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge841_GATE_N (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge865_GATE (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s902_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s917_SLEEP_B (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_6_0_clk_X (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_CLK_N (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s911_GATE_N (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s912_GATE (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s913_GATE_N (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s914_GATE_N (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s915_GATE_N (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s916_GATE (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s918_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s919_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_7_0_clk_X (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_CLK_N (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_CLK_N (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge811_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge815_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge834_GATE (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge848_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_8_0_clk_X (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c257_CLK_N (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_CLK_N (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge804_CLK_N (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge844_GATE (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge861_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s893_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_10_0_clk_X (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_CLK_N (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge854_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge855_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge881_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s904_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s906_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s920_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s927_GATE_N (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_12_0_clk_X (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_CLK_N (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge847_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge849_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge858_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge859_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge864_GATE (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge867_GATE_N (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge868_GATE_N (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge869_GATE (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s925_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s926_GATE_N (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s928_GATE (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s929_GATE_N (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_13_0_clk_X (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge845_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge856_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge860_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge872_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge873_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge878_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge880_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_15_0_clk_X (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net491_A (.DIODE(clknet_0_net491));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net491_A (.DIODE(clknet_0_net491));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net491_X (.DIODE(clknet_0_net491));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_S0 (.DIODE(clknet_1_1__leaf_net491));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net491_X (.DIODE(clknet_1_1__leaf_net491));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_A1 (.DIODE(clknet_1_1__leaf_net489));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_A2 (.DIODE(clknet_1_1__leaf_net489));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_A0 (.DIODE(clknet_1_1__leaf_net489));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net489_X (.DIODE(clknet_1_1__leaf_net489));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_SET_B (.DIODE(clknet_1_0__leaf_net764));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_SET_B (.DIODE(clknet_1_0__leaf_net764));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_SET_B (.DIODE(clknet_1_0__leaf_net764));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_S1 (.DIODE(clknet_1_0__leaf_net764));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net764_X (.DIODE(clknet_1_0__leaf_net764));
 sky130_fd_sc_hd__diode_2 ANTENNA_c263_S1 (.DIODE(clknet_1_0__leaf_net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net891_X (.DIODE(clknet_1_0__leaf_net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_output118_A (.DIODE(clknet_1_1__leaf_net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net891_X (.DIODE(clknet_1_1__leaf_net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net889_A (.DIODE(clknet_0_net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net889_A (.DIODE(clknet_0_net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net889_X (.DIODE(clknet_0_net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_S1 (.DIODE(clknet_1_0__leaf_net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c215_B1 (.DIODE(clknet_1_0__leaf_net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_A4 (.DIODE(clknet_1_0__leaf_net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_A3 (.DIODE(clknet_1_0__leaf_net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_B1 (.DIODE(clknet_1_0__leaf_net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_output116_A (.DIODE(clknet_1_0__leaf_net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net889_X (.DIODE(clknet_1_0__leaf_net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c220_B1 (.DIODE(clknet_1_1__leaf_net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c221_B1 (.DIODE(clknet_1_1__leaf_net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c222_B1 (.DIODE(clknet_1_1__leaf_net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_B1 (.DIODE(clknet_1_1__leaf_net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_S1 (.DIODE(clknet_1_1__leaf_net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_A4 (.DIODE(clknet_1_1__leaf_net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_SET_B (.DIODE(clknet_1_1__leaf_net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_SCE (.DIODE(clknet_1_1__leaf_net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_S1 (.DIODE(clknet_1_1__leaf_net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net889_X (.DIODE(clknet_1_1__leaf_net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net370_A (.DIODE(clknet_0_net370));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net370_A (.DIODE(clknet_0_net370));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net370_X (.DIODE(clknet_0_net370));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_A2 (.DIODE(clknet_1_1__leaf_net370));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_S0 (.DIODE(clknet_1_1__leaf_net370));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net370_X (.DIODE(clknet_1_1__leaf_net370));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net366_A (.DIODE(clknet_0_net366));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net366_A (.DIODE(clknet_0_net366));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net366_X (.DIODE(clknet_0_net366));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_A2 (.DIODE(clknet_1_1__leaf_net366));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_A2 (.DIODE(clknet_1_1__leaf_net366));
 sky130_fd_sc_hd__diode_2 ANTENNA_c496_A1 (.DIODE(clknet_1_1__leaf_net366));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_S0 (.DIODE(clknet_1_1__leaf_net366));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_A2 (.DIODE(clknet_1_1__leaf_net366));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net366_X (.DIODE(clknet_1_1__leaf_net366));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net364_A (.DIODE(clknet_0_net364));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net364_A (.DIODE(clknet_0_net364));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net364_X (.DIODE(clknet_0_net364));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net363_A (.DIODE(clknet_0_net363));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net363_A (.DIODE(clknet_0_net363));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net363_X (.DIODE(clknet_0_net363));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net883_A (.DIODE(clknet_0_net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net883_A (.DIODE(clknet_0_net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net883_X (.DIODE(clknet_0_net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_A1 (.DIODE(clknet_1_1__leaf_net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_A1 (.DIODE(clknet_1_1__leaf_net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_output110_A (.DIODE(clknet_1_1__leaf_net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net883_X (.DIODE(clknet_1_1__leaf_net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net354_A (.DIODE(clknet_0_net354));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net354_A (.DIODE(clknet_0_net354));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net354_X (.DIODE(clknet_0_net354));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_A2 (.DIODE(clknet_1_0__leaf_net354));
 sky130_fd_sc_hd__diode_2 ANTENNA_c482_S1 (.DIODE(clknet_1_0__leaf_net354));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net354_X (.DIODE(clknet_1_0__leaf_net354));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net353_A (.DIODE(clknet_0_net353));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net353_A (.DIODE(clknet_0_net353));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net353_X (.DIODE(clknet_0_net353));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_A1 (.DIODE(clknet_1_0__leaf_net353));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net353_X (.DIODE(clknet_1_0__leaf_net353));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net346_A (.DIODE(clknet_0_net346));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net346_A (.DIODE(clknet_0_net346));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net346_X (.DIODE(clknet_0_net346));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_A1 (.DIODE(clknet_1_1__leaf_net346));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_A1 (.DIODE(clknet_1_1__leaf_net346));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_A3 (.DIODE(clknet_1_1__leaf_net346));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net346_X (.DIODE(clknet_1_1__leaf_net346));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_A1 (.DIODE(clknet_1_0__leaf_net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_A3 (.DIODE(clknet_1_0__leaf_net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_SCD (.DIODE(clknet_1_0__leaf_net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_A3 (.DIODE(clknet_1_0__leaf_net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_A4 (.DIODE(clknet_1_0__leaf_net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_A4 (.DIODE(clknet_1_0__leaf_net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_SET_B (.DIODE(clknet_1_0__leaf_net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_A2 (.DIODE(clknet_1_0__leaf_net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net887_X (.DIODE(clknet_1_0__leaf_net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_S1 (.DIODE(clknet_1_1__leaf_net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_S0 (.DIODE(clknet_1_1__leaf_net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_A1 (.DIODE(clknet_1_1__leaf_net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_SCD (.DIODE(clknet_1_1__leaf_net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_A4 (.DIODE(clknet_1_1__leaf_net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_A3 (.DIODE(clknet_1_1__leaf_net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_S1 (.DIODE(clknet_1_1__leaf_net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_output114_A (.DIODE(clknet_1_1__leaf_net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net887_X (.DIODE(clknet_1_1__leaf_net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net348_A (.DIODE(clknet_0_net348));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net348_A (.DIODE(clknet_0_net348));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net348_X (.DIODE(clknet_0_net348));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_A0 (.DIODE(clknet_1_1__leaf_net348));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net348_X (.DIODE(clknet_1_1__leaf_net348));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net345_A (.DIODE(clknet_0_net345));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net345_A (.DIODE(clknet_0_net345));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net345_X (.DIODE(clknet_0_net345));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_S0 (.DIODE(clknet_1_1__leaf_net345));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_A2 (.DIODE(clknet_1_1__leaf_net345));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_A0 (.DIODE(clknet_1_1__leaf_net345));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net345_X (.DIODE(clknet_1_1__leaf_net345));
 sky130_fd_sc_hd__diode_2 ANTENNA_c232_A1 (.DIODE(clknet_1_0__leaf_net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_S1 (.DIODE(clknet_1_0__leaf_net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_c234_A0 (.DIODE(clknet_1_0__leaf_net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_c237_A2 (.DIODE(clknet_1_0__leaf_net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_c239_S1 (.DIODE(clknet_1_0__leaf_net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_D (.DIODE(clknet_1_0__leaf_net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_A4 (.DIODE(clknet_1_0__leaf_net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_B1 (.DIODE(clknet_1_0__leaf_net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_c366_A2 (.DIODE(clknet_1_0__leaf_net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_A1 (.DIODE(clknet_1_0__leaf_net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net132_X (.DIODE(clknet_1_0__leaf_net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_c256_A3 (.DIODE(clknet_1_1__leaf_net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_c257_SCE (.DIODE(clknet_1_1__leaf_net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_c258_A3 (.DIODE(clknet_1_1__leaf_net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_c259_B1 (.DIODE(clknet_1_1__leaf_net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_RESET_B (.DIODE(clknet_1_1__leaf_net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net132_X (.DIODE(clknet_1_1__leaf_net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_c260_A2 (.DIODE(clknet_1_0__leaf_net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c261_A2 (.DIODE(clknet_1_0__leaf_net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c262_S0 (.DIODE(clknet_1_0__leaf_net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c263_A2 (.DIODE(clknet_1_0__leaf_net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net894_X (.DIODE(clknet_1_0__leaf_net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_output121_A (.DIODE(clknet_1_1__leaf_net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net894_X (.DIODE(clknet_1_1__leaf_net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c261_A1 (.DIODE(clknet_1_0__leaf_net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_c262_A1 (.DIODE(clknet_1_0__leaf_net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net901_X (.DIODE(clknet_1_0__leaf_net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_c263_A0 (.DIODE(clknet_1_1__leaf_net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_output128_A (.DIODE(clknet_1_1__leaf_net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net901_X (.DIODE(clknet_1_1__leaf_net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net898_A (.DIODE(clknet_0_net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net898_A (.DIODE(clknet_0_net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net898_X (.DIODE(clknet_0_net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c259_A1 (.DIODE(clknet_1_0__leaf_net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c260_A3 (.DIODE(clknet_1_0__leaf_net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c261_A0 (.DIODE(clknet_1_0__leaf_net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net898_X (.DIODE(clknet_1_0__leaf_net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c262_A3 (.DIODE(clknet_1_1__leaf_net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c263_A1 (.DIODE(clknet_1_1__leaf_net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_output125_A (.DIODE(clknet_1_1__leaf_net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net898_X (.DIODE(clknet_1_1__leaf_net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c258_A1 (.DIODE(clknet_1_0__leaf_net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_c259_A3 (.DIODE(clknet_1_0__leaf_net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_c260_A4 (.DIODE(clknet_1_0__leaf_net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net895_X (.DIODE(clknet_1_0__leaf_net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_c257_RESET_B (.DIODE(clknet_1_1__leaf_net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_c261_S0 (.DIODE(clknet_1_1__leaf_net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_output122_A (.DIODE(clknet_1_1__leaf_net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net895_X (.DIODE(clknet_1_1__leaf_net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net890_A (.DIODE(clknet_0_net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net890_A (.DIODE(clknet_0_net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net890_X (.DIODE(clknet_0_net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c229_A3 (.DIODE(clknet_1_0__leaf_net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c231_S1 (.DIODE(clknet_1_0__leaf_net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_RESET_B (.DIODE(clknet_1_0__leaf_net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_A0 (.DIODE(clknet_1_0__leaf_net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net890_X (.DIODE(clknet_1_0__leaf_net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c256_A4 (.DIODE(clknet_1_1__leaf_net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c257_SET_B (.DIODE(clknet_1_1__leaf_net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_S0 (.DIODE(clknet_1_1__leaf_net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_output117_A (.DIODE(clknet_1_1__leaf_net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net890_X (.DIODE(clknet_1_1__leaf_net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_A1 (.DIODE(clknet_1_1__leaf_net184));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_S0 (.DIODE(clknet_1_1__leaf_net184));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_RESET_B (.DIODE(clknet_1_1__leaf_net184));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net184_X (.DIODE(clknet_1_1__leaf_net184));
 sky130_fd_sc_hd__clkbuf_2 split1 (.A(net949),
    .X(net948));
 sky130_fd_sc_hd__clkbuf_2 split2 (.A(net702),
    .X(net949));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_511 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_535 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_254 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_507 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_171 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_415 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_20 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_115 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_143 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_338 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_616 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_8 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_497 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_582 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_382 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_140 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_283 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_624 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_10 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_507 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_226 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_146 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_385 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_590 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_130 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_612 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_270 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_451 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_158 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_411 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_591 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_339 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_563 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_115 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_5 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_14 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_580 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_6 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_87 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_8 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_224 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_553 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_525 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_170 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_8 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_50 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_20 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_564 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_413 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_422 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_600 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_245 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_5 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_256 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_336 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_617 ();
endmodule
