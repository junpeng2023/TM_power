module netlist_1 (clk,
    in0,
    in1,
    in10,
    in11,
    in12,
    in13,
    in14,
    in15,
    in16,
    in17,
    in18,
    in19,
    in2,
    in20,
    in21,
    in22,
    in23,
    in24,
    in3,
    in4,
    in5,
    in6,
    in7,
    in8,
    in9,
    out0,
    out1,
    out10,
    out11,
    out12,
    out13,
    out14,
    out15,
    out16,
    out17,
    out18,
    out19,
    out2,
    out20,
    out21,
    out22,
    out23,
    out24,
    out3,
    out4,
    out5,
    out6,
    out7,
    out8,
    out9,
    rst);
 input clk;
 input in0;
 input in1;
 input in10;
 input in11;
 input in12;
 input in13;
 input in14;
 input in15;
 input in16;
 input in17;
 input in18;
 input in19;
 input in2;
 input in20;
 input in21;
 input in22;
 input in23;
 input in24;
 input in3;
 input in4;
 input in5;
 input in6;
 input in7;
 input in8;
 input in9;
 output out0;
 output out1;
 output out10;
 output out11;
 output out12;
 output out13;
 output out14;
 output out15;
 output out16;
 output out17;
 output out18;
 output out19;
 output out2;
 output out20;
 output out21;
 output out22;
 output out23;
 output out24;
 output out3;
 output out4;
 output out5;
 output out6;
 output out7;
 output out8;
 output out9;
 input rst;

 wire net0;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net629;
 wire net63;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net64;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net65;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net66;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net67;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net68;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net69;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net7;
 wire net70;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net71;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net72;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net73;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net74;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net75;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net76;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net77;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net78;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net79;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net8;
 wire net80;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net81;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net82;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net83;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net84;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net85;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net86;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net87;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net88;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net89;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net9;
 wire net90;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net91;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net92;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net93;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net94;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net95;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net96;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net97;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net98;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net99;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net556;
 wire net628;
 wire net759;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_0_net1020;
 wire clknet_1_0__leaf_net1020;
 wire clknet_1_1__leaf_net1020;
 wire clknet_0_net994;
 wire clknet_1_0__leaf_net994;
 wire clknet_1_1__leaf_net994;
 wire clknet_0_net558;
 wire clknet_1_0__leaf_net558;
 wire clknet_1_1__leaf_net558;
 wire clknet_0_net563;
 wire clknet_1_0__leaf_net563;
 wire clknet_1_1__leaf_net563;
 wire clknet_0_net993;
 wire clknet_1_0__leaf_net993;
 wire clknet_1_1__leaf_net993;
 wire clknet_0_net694;
 wire clknet_1_0__leaf_net694;
 wire clknet_1_1__leaf_net694;
 wire clknet_0_net949;
 wire clknet_1_0__leaf_net949;
 wire clknet_1_1__leaf_net949;
 wire clknet_0_net710;
 wire clknet_1_0__leaf_net710;
 wire clknet_1_1__leaf_net710;
 wire clknet_0_net717;
 wire clknet_1_0__leaf_net717;
 wire clknet_1_1__leaf_net717;
 wire clknet_0_net719;
 wire clknet_1_0__leaf_net719;
 wire clknet_1_1__leaf_net719;
 wire clknet_0_net712;
 wire clknet_1_0__leaf_net712;
 wire clknet_1_1__leaf_net712;
 wire clknet_0_net442;
 wire clknet_1_0__leaf_net442;
 wire clknet_1_1__leaf_net442;
 wire clknet_0_net447;
 wire clknet_1_0__leaf_net447;
 wire clknet_1_1__leaf_net447;
 wire clknet_0_net914;
 wire clknet_1_0__leaf_net914;
 wire clknet_1_1__leaf_net914;
 wire clknet_0_net985;
 wire clknet_1_0__leaf_net985;
 wire clknet_1_1__leaf_net985;
 wire clknet_0_net984;
 wire clknet_1_0__leaf_net984;
 wire clknet_1_1__leaf_net984;
 wire clknet_0_net498;
 wire clknet_1_0__leaf_net498;
 wire clknet_1_1__leaf_net498;
 wire clknet_0_net357;
 wire clknet_1_0__leaf_net357;
 wire clknet_1_1__leaf_net357;
 wire clknet_0_net197;
 wire clknet_1_0__leaf_net197;
 wire clknet_1_1__leaf_net197;
 wire clknet_0_net201;
 wire clknet_1_0__leaf_net201;
 wire clknet_1_1__leaf_net201;
 wire clknet_0_net85;
 wire clknet_1_0__leaf_net85;
 wire clknet_1_1__leaf_net85;
 wire clknet_0_net205;
 wire clknet_1_0__leaf_net205;
 wire clknet_1_1__leaf_net205;
 wire clknet_0_net208;
 wire clknet_1_0__leaf_net208;
 wire clknet_1_1__leaf_net208;
 wire clknet_0_net226;
 wire clknet_1_0__leaf_net226;
 wire clknet_1_1__leaf_net226;
 wire clknet_0_net210;
 wire clknet_1_0__leaf_net210;
 wire clknet_1_1__leaf_net210;
 wire clknet_0_net207;
 wire clknet_1_0__leaf_net207;
 wire clknet_1_1__leaf_net207;
 wire clknet_0_net213;
 wire clknet_1_0__leaf_net213;
 wire clknet_1_1__leaf_net213;
 wire clknet_0_net87;
 wire clknet_1_0__leaf_net87;
 wire clknet_1_1__leaf_net87;
 wire clknet_0_net91;
 wire clknet_1_0__leaf_net91;
 wire clknet_1_1__leaf_net91;
 wire clknet_0_net89;
 wire clknet_1_0__leaf_net89;
 wire clknet_1_1__leaf_net89;
 wire clknet_0_net88;
 wire clknet_1_0__leaf_net88;
 wire clknet_1_1__leaf_net88;
 wire clknet_0_net95;
 wire clknet_1_0__leaf_net95;
 wire clknet_1_1__leaf_net95;
 wire clknet_0_net79;
 wire clknet_1_0__leaf_net79;
 wire clknet_1_1__leaf_net79;
 wire clknet_0_net81;
 wire clknet_1_0__leaf_net81;
 wire clknet_1_1__leaf_net81;
 wire clknet_0_net951;
 wire clknet_1_0__leaf_net951;
 wire clknet_1_1__leaf_net951;
 wire clknet_0_net42;
 wire clknet_1_0__leaf_net42;
 wire clknet_1_1__leaf_net42;
 wire clknet_0_net29;
 wire clknet_1_0__leaf_net29;
 wire clknet_1_1__leaf_net29;
 wire clknet_0_net912;
 wire clknet_1_0__leaf_net912;
 wire clknet_1_1__leaf_net912;
 wire clknet_0_net26;
 wire clknet_1_0__leaf_net26;
 wire clknet_1_1__leaf_net26;
 wire clknet_0_net21;
 wire clknet_1_0__leaf_net21;
 wire clknet_1_1__leaf_net21;
 wire clknet_0_net24;
 wire clknet_1_0__leaf_net24;
 wire clknet_1_1__leaf_net24;
 wire clknet_0_net20;
 wire clknet_1_0__leaf_net20;
 wire clknet_1_1__leaf_net20;
 wire clknet_0_net25;
 wire clknet_1_0__leaf_net25;
 wire clknet_1_1__leaf_net25;
 wire clknet_0_net23;
 wire clknet_1_0__leaf_net23;
 wire clknet_1_1__leaf_net23;
 wire clknet_0_net34;
 wire clknet_1_0__leaf_net34;
 wire clknet_1_1__leaf_net34;
 wire clknet_0_net161;
 wire clknet_1_0__leaf_net161;
 wire clknet_1_1__leaf_net161;
 wire clknet_0_net163;
 wire clknet_1_0__leaf_net163;
 wire clknet_1_1__leaf_net163;
 wire clknet_0_net168;
 wire clknet_1_0__leaf_net168;
 wire clknet_1_1__leaf_net168;
 wire clknet_0_net162;
 wire clknet_1_0__leaf_net162;
 wire clknet_1_1__leaf_net162;
 wire clknet_0_net27;
 wire clknet_1_0__leaf_net27;
 wire clknet_1_1__leaf_net27;
 wire clknet_0_net22;
 wire clknet_1_0__leaf_net22;
 wire clknet_1_1__leaf_net22;
 wire clknet_0_net352;
 wire clknet_1_0__leaf_net352;
 wire clknet_1_1__leaf_net352;
 wire clknet_0_net353;
 wire clknet_1_0__leaf_net353;
 wire clknet_1_1__leaf_net353;
 wire clknet_0_net950;
 wire clknet_1_0__leaf_net950;
 wire clknet_1_1__leaf_net950;
 wire clknet_0_net764;
 wire clknet_1_0__leaf_net764;
 wire clknet_1_1__leaf_net764;
 wire clknet_0_net482;
 wire clknet_1_0__leaf_net482;
 wire clknet_1_1__leaf_net482;
 wire clknet_0_net479;
 wire clknet_1_0__leaf_net479;
 wire clknet_1_1__leaf_net479;
 wire clknet_0_net491;
 wire clknet_1_0__leaf_net491;
 wire clknet_1_1__leaf_net491;
 wire clknet_0_net496;
 wire clknet_1_0__leaf_net496;
 wire clknet_1_1__leaf_net496;
 wire clknet_0_net493;
 wire clknet_1_0__leaf_net493;
 wire clknet_1_1__leaf_net493;
 wire clknet_0_net747;
 wire clknet_1_0__leaf_net747;
 wire clknet_1_1__leaf_net747;
 wire clknet_0_net318;
 wire clknet_1_0__leaf_net318;
 wire clknet_1_1__leaf_net318;
 wire clknet_0_net325;
 wire clknet_1_0__leaf_net325;
 wire clknet_1_1__leaf_net325;
 wire clknet_0_net320;
 wire clknet_1_0__leaf_net320;
 wire clknet_1_1__leaf_net320;
 wire clknet_0_net321;
 wire clknet_1_0__leaf_net321;
 wire clknet_1_1__leaf_net321;
 wire clknet_0_net317;
 wire clknet_1_0__leaf_net317;
 wire clknet_1_1__leaf_net317;
 wire clknet_0_net324;
 wire clknet_1_0__leaf_net324;
 wire clknet_1_1__leaf_net324;
 wire clknet_0_net329;
 wire clknet_1_0__leaf_net329;
 wire clknet_1_1__leaf_net329;
 wire clknet_0_net326;
 wire clknet_1_0__leaf_net326;
 wire clknet_1_1__leaf_net326;
 wire clknet_0_net330;
 wire clknet_1_0__leaf_net330;
 wire clknet_1_1__leaf_net330;
 wire clknet_0_net328;
 wire clknet_1_0__leaf_net328;
 wire clknet_1_1__leaf_net328;
 wire clknet_0_net915;
 wire clknet_1_0__leaf_net915;
 wire clknet_1_1__leaf_net915;
 wire clknet_0_net160;
 wire clknet_1_0__leaf_net160;
 wire clknet_1_1__leaf_net160;
 wire clknet_0_net144;
 wire clknet_1_0__leaf_net144;
 wire clknet_1_1__leaf_net144;
 wire clknet_0_net147;
 wire clknet_1_0__leaf_net147;
 wire clknet_1_1__leaf_net147;
 wire clknet_0_net145;
 wire clknet_1_0__leaf_net145;
 wire clknet_1_1__leaf_net145;
 wire clknet_0_net272;
 wire clknet_1_0__leaf_net272;
 wire clknet_1_1__leaf_net272;
 wire clknet_0_net126;
 wire clknet_1_0__leaf_net126;
 wire clknet_1_1__leaf_net126;
 wire clknet_0_net129;
 wire clknet_1_0__leaf_net129;
 wire clknet_1_1__leaf_net129;
 wire clknet_0_net127;
 wire clknet_1_0__leaf_net127;
 wire clknet_1_1__leaf_net127;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;

 sky130_fd_sc_hd__a21bo_1 c100 (.A1(net76),
    .A2(net67),
    .B1_N(net71),
    .X(net77));
 sky130_fd_sc_hd__a21bo_1 c101 (.A1(net57),
    .A2(net76),
    .B1_N(net963),
    .X(net78));
 sky130_fd_sc_hd__xnor2_1 c102 (.A(net73),
    .B(clknet_1_0__leaf_net985),
    .Y(net79));
 sky130_fd_sc_hd__xnor2_1 c103 (.A(net75),
    .B(net69),
    .Y(net80));
 sky130_fd_sc_hd__a21bo_1 c104 (.A1(net80),
    .A2(net76),
    .B1_N(clknet_1_0__leaf_net79),
    .X(net81));
 sky130_fd_sc_hd__mux4_1 c105 (.A0(net74),
    .A1(clknet_1_0__leaf_net79),
    .A2(net80),
    .A3(clknet_1_0__leaf_net81),
    .S0(net66),
    .S1(net43),
    .X(net82));
 sky130_fd_sc_hd__a31o_1 c106 (.A1(clknet_1_1__leaf_net79),
    .A2(net80),
    .A3(net76),
    .B1(net67),
    .X(net83));
 sky130_fd_sc_hd__mux4_1 c107 (.A0(net72),
    .A1(net80),
    .A2(net43),
    .A3(net68),
    .S0(clknet_1_0__leaf_net985),
    .S1(net987),
    .X(net84));
 sky130_fd_sc_hd__buf_1 c108 (.A(clknet_1_1__leaf_net985),
    .X(net85));
 sky130_fd_sc_hd__clkbuf_1 c109 (.A(net1039),
    .X(net86));
 sky130_fd_sc_hd__buf_1 c110 (.A(clknet_1_0__leaf_net85),
    .X(net87));
 sky130_fd_sc_hd__xnor2_1 c111 (.A(clknet_1_0__leaf_net87),
    .B(net73),
    .Y(net88));
 sky130_fd_sc_hd__xnor2_1 c112 (.A(clknet_1_0__leaf_net88),
    .B(clknet_1_0__leaf_net87),
    .Y(net89));
 sky130_fd_sc_hd__clkbuf_1 c113 (.A(net910),
    .X(net90));
 sky130_fd_sc_hd__buf_1 c114 (.A(clknet_1_1__leaf_net87),
    .X(net91));
 sky130_fd_sc_hd__buf_1 c115 (.A(net73),
    .X(net92));
 sky130_fd_sc_hd__clkbuf_2 c116 (.A(net90),
    .X(net93));
 sky130_fd_sc_hd__a21bo_1 c117 (.A1(net90),
    .A2(clknet_1_0__leaf_net88),
    .B1_N(net92),
    .X(net94));
 sky130_fd_sc_hd__xnor2_1 c118 (.A(clknet_1_1__leaf_net88),
    .B(net93),
    .Y(net95));
 sky130_fd_sc_hd__xnor2_1 c119 (.A(net92),
    .B(net93),
    .Y(net96));
 sky130_fd_sc_hd__buf_1 c120 (.A(net910),
    .X(net97));
 sky130_fd_sc_hd__dfbbn_1 c121 (.CLK_N(clknet_4_0_0_clk),
    .D(clknet_1_0__leaf_net89),
    .RESET_B(clknet_1_0__leaf_net95),
    .SET_B(net93),
    .Q(net99),
    .Q_N(net98));
 sky130_fd_sc_hd__dfbbn_2 c122 (.CLK_N(clknet_4_0_0_clk),
    .D(net1051),
    .RESET_B(net97),
    .SET_B(clknet_1_1__leaf_net95),
    .Q(net101),
    .Q_N(net100));
 sky130_fd_sc_hd__dfbbp_1 c123 (.CLK(clknet_4_0_0_clk),
    .D(clknet_1_0__leaf_net95),
    .RESET_B(net99),
    .SET_B(net92),
    .Q(net103),
    .Q_N(net102));
 sky130_fd_sc_hd__sdfxbp_1 c124 (.CLK(clknet_4_0_0_clk),
    .D(clknet_1_0__leaf_net95),
    .SCD(net98),
    .SCE(net101),
    .Q(net105),
    .Q_N(net104));
 sky130_fd_sc_hd__sdfrbp_1 c125 (.CLK(clknet_4_0_0_clk),
    .D(clknet_1_0__leaf_net91),
    .RESET_B(net1036),
    .SCD(net100),
    .SCE(clknet_1_1__leaf_net95),
    .Q(net107),
    .Q_N(net106));
 sky130_fd_sc_hd__a21bo_1 c126 (.A1(net93),
    .A2(net96),
    .B1_N(net106),
    .X(net108));
 sky130_fd_sc_hd__sdfxbp_1 c127 (.CLK(clknet_4_0_0_clk),
    .D(net97),
    .SCD(net1052),
    .SCE(net108),
    .Q(net110),
    .Q_N(net109));
 sky130_fd_sc_hd__a21bo_1 c128 (.A1(net107),
    .A2(net108),
    .B1_N(net109),
    .X(net111));
 sky130_fd_sc_hd__sdfbbn_1 c129 (.CLK_N(clknet_4_0_0_clk),
    .D(net105),
    .RESET_B(net110),
    .SCD(net97),
    .SCE(clknet_1_1__leaf_net95),
    .SET_B(net93),
    .Q(net113),
    .Q_N(net112));
 sky130_fd_sc_hd__a21bo_1 c130 (.A1(net86),
    .A2(net113),
    .B1_N(net108),
    .X(net114));
 sky130_fd_sc_hd__a41o_1 c131 (.A1(net96),
    .A2(net110),
    .A3(net112),
    .A4(net104),
    .B1(clknet_1_1__leaf_net95),
    .X(net115));
 sky130_fd_sc_hd__clkbuf_4 c132 (.A(in18),
    .X(net116));
 sky130_fd_sc_hd__dlymetal6s2s_1 c133 (.A(net116),
    .X(net117));
 sky130_fd_sc_hd__a21bo_2 c134 (.A1(net117),
    .A2(net1002),
    .B1_N(net116),
    .X(net118));
 sky130_fd_sc_hd__xnor2_1 c135 (.A(net116),
    .B(net117),
    .Y(net119));
 sky130_fd_sc_hd__buf_1 c136 (.A(net907),
    .X(net120));
 sky130_fd_sc_hd__xnor2_1 c137 (.A(net116),
    .B(net120),
    .Y(net121));
 sky130_fd_sc_hd__xnor2_1 c138 (.A(net117),
    .B(net116),
    .Y(net122));
 sky130_fd_sc_hd__buf_1 c139 (.A(net907),
    .X(net123));
 sky130_fd_sc_hd__a21bo_1 c140 (.A1(net121),
    .A2(net123),
    .B1_N(net116),
    .X(net124));
 sky130_fd_sc_hd__buf_1 c141 (.A(clknet_1_1__leaf_net915),
    .X(net125));
 sky130_fd_sc_hd__buf_1 c142 (.A(clknet_1_1__leaf_net915),
    .X(net126));
 sky130_fd_sc_hd__a21bo_1 c143 (.A1(clknet_1_0__leaf_net126),
    .A2(net116),
    .B1_N(net121),
    .X(net127));
 sky130_fd_sc_hd__mux4_1 c144 (.A0(clknet_1_1__leaf_net127),
    .A1(net117),
    .A2(net122),
    .A3(clknet_1_1__leaf_net126),
    .S0(net116),
    .S1(net119),
    .X(net128));
 sky130_fd_sc_hd__a21bo_1 c145 (.A1(net1011),
    .A2(clknet_1_1__leaf_net126),
    .B1_N(net870),
    .X(net129));
 sky130_fd_sc_hd__a21bo_2 c146 (.A1(net120),
    .A2(net1005),
    .B1_N(net556),
    .X(net130));
 sky130_fd_sc_hd__buf_1 c147 (.A(net980),
    .X(net131));
 sky130_fd_sc_hd__buf_1 c148 (.A(net976),
    .X(net132));
 sky130_fd_sc_hd__mux4_1 c149 (.A0(clknet_1_0__leaf_net129),
    .A1(net131),
    .A2(net130),
    .A3(net123),
    .S0(net116),
    .S1(clknet_1_0__leaf_net126),
    .X(net133));
 sky130_fd_sc_hd__clkbuf_1 c150 (.A(net932),
    .X(net134));
 sky130_fd_sc_hd__a21bo_1 c151 (.A1(net996),
    .A2(net132),
    .B1_N(clknet_1_1__leaf_net126),
    .X(net135));
 sky130_fd_sc_hd__mux4_1 c152 (.A0(net133),
    .A1(net123),
    .A2(clknet_1_1__leaf_net129),
    .A3(clknet_1_0__leaf_net126),
    .S0(net130),
    .S1(net116),
    .X(net136));
 sky130_fd_sc_hd__a21bo_1 c153 (.A1(net135),
    .A2(net134),
    .B1_N(net136),
    .X(net137));
 sky130_fd_sc_hd__clkbuf_4 c154 (.A(net1006),
    .X(net138));
 sky130_fd_sc_hd__clkbuf_4 c155 (.A(net138),
    .X(net139));
 sky130_fd_sc_hd__xnor2_4 c156 (.A(net139),
    .B(net138),
    .Y(net140));
 sky130_fd_sc_hd__clkbuf_1 c157 (.A(net975),
    .X(net141));
 sky130_fd_sc_hd__xnor2_4 c158 (.A(net139),
    .B(net999),
    .Y(net142));
 sky130_fd_sc_hd__buf_1 c159 (.A(net975),
    .X(net143));
 sky130_fd_sc_hd__buf_1 c160 (.A(clknet_1_0__leaf_net915),
    .X(net144));
 sky130_fd_sc_hd__xnor2_1 c161 (.A(clknet_1_0__leaf_net144),
    .B(net138),
    .Y(net145));
 sky130_fd_sc_hd__buf_1 c162 (.A(net916),
    .X(net146));
 sky130_fd_sc_hd__a21bo_1 c163 (.A1(net143),
    .A2(clknet_1_1__leaf_net144),
    .B1_N(net146),
    .X(net147));
 sky130_fd_sc_hd__sdfbbp_1 c164 (.CLK(clknet_4_7_0_clk),
    .D(net146),
    .RESET_B(clknet_1_0__leaf_net147),
    .SCD(net139),
    .SCE(net142),
    .SET_B(net140),
    .Q(net149),
    .Q_N(net148));
 sky130_fd_sc_hd__buf_1 c165 (.A(clknet_1_0__leaf_net915),
    .X(net150));
 sky130_fd_sc_hd__a21bo_1 c166 (.A1(net149),
    .A2(net143),
    .B1_N(clknet_1_1__leaf_net145),
    .X(net151));
 sky130_fd_sc_hd__clkbuf_1 c167 (.A(net957),
    .X(net152));
 sky130_fd_sc_hd__buf_1 c168 (.A(net976),
    .X(net153));
 sky130_fd_sc_hd__mux4_1 c169 (.A0(clknet_1_0__leaf_net144),
    .A1(clknet_1_0__leaf_net147),
    .A2(net149),
    .A3(net138),
    .S0(net13),
    .S1(net139),
    .X(net154));
 sky130_fd_sc_hd__a31o_1 c170 (.A1(net153),
    .A2(net146),
    .A3(net148),
    .B1(net142),
    .X(net155));
 sky130_fd_sc_hd__a21bo_1 c171 (.A1(net141),
    .A2(net146),
    .B1_N(net938),
    .X(net156));
 sky130_fd_sc_hd__mux4_1 c172 (.A0(clknet_1_1__leaf_net147),
    .A1(net153),
    .A2(net138),
    .A3(net140),
    .S0(net142),
    .S1(net938),
    .X(net157));
 sky130_fd_sc_hd__a21bo_1 c173 (.A1(net150),
    .A2(net156),
    .B1_N(net153),
    .X(net158));
 sky130_fd_sc_hd__xnor2_1 c174 (.A(net156),
    .B(net907),
    .Y(net159));
 sky130_fd_sc_hd__a21bo_1 c175 (.A1(net158),
    .A2(net159),
    .B1_N(net146),
    .X(net160));
 sky130_fd_sc_hd__xnor2_1 c176 (.A(clknet_1_1__leaf_net42),
    .B(net948),
    .Y(net161));
 sky130_fd_sc_hd__xnor2_1 c177 (.A(clknet_1_1__leaf_net145),
    .B(clknet_1_1__leaf_net161),
    .Y(net162));
 sky130_fd_sc_hd__xnor2_1 c178 (.A(net1015),
    .B(clknet_1_0__leaf_net161),
    .Y(net163));
 sky130_fd_sc_hd__clkbuf_1 c179 (.A(net904),
    .X(net164));
 sky130_fd_sc_hd__clkbuf_2 c180 (.A(net904),
    .X(net165));
 sky130_fd_sc_hd__clkbuf_2 c181 (.A(net976),
    .X(net166));
 sky130_fd_sc_hd__xnor2_1 c182 (.A(net166),
    .B(net165),
    .Y(net167));
 sky130_fd_sc_hd__xnor2_1 c183 (.A(clknet_1_1__leaf_net163),
    .B(net166),
    .Y(net168));
 sky130_fd_sc_hd__xnor2_1 c184 (.A(net167),
    .B(clknet_1_1__leaf_net163),
    .Y(net169));
 sky130_fd_sc_hd__buf_1 c185 (.A(net942),
    .X(net170));
 sky130_fd_sc_hd__buf_1 c186 (.A(net947),
    .X(net171));
 sky130_fd_sc_hd__a21bo_1 c187 (.A1(clknet_1_0__leaf_net168),
    .A2(net166),
    .B1_N(net165),
    .X(net172));
 sky130_fd_sc_hd__mux4_1 c188 (.A0(clknet_1_0__leaf_net163),
    .A1(clknet_1_1__leaf_net168),
    .A2(net171),
    .A3(net165),
    .S0(net166),
    .S1(net904),
    .X(net173));
 sky130_fd_sc_hd__a41o_1 c189 (.A1(net171),
    .A2(net166),
    .A3(clknet_1_0__leaf_net163),
    .A4(clknet_1_0__leaf_net162),
    .B1(net904),
    .X(net174));
 sky130_fd_sc_hd__clkbuf_1 c190 (.A(net954),
    .X(net175));
 sky130_fd_sc_hd__a21bo_1 c191 (.A1(net166),
    .A2(net170),
    .B1_N(net171),
    .X(net176));
 sky130_fd_sc_hd__xnor2_1 c192 (.A(net170),
    .B(net171),
    .Y(net177));
 sky130_fd_sc_hd__xnor2_1 c193 (.A(net164),
    .B(net177),
    .Y(net178));
 sky130_fd_sc_hd__clkbuf_1 c194 (.A(net947),
    .X(net179));
 sky130_fd_sc_hd__xnor2_1 c195 (.A(net175),
    .B(net179),
    .Y(net180));
 sky130_fd_sc_hd__xnor2_1 c196 (.A(net177),
    .B(net180),
    .Y(net181));
 sky130_fd_sc_hd__xnor2_1 c197 (.A(clknet_1_0__leaf_net161),
    .B(net178),
    .Y(net182));
 sky130_fd_sc_hd__clkbuf_4 c198 (.A(net930),
    .X(net183));
 sky130_fd_sc_hd__buf_1 c199 (.A(net183),
    .X(net184));
 sky130_fd_sc_hd__clkbuf_1 c200 (.A(net930),
    .X(net185));
 sky130_fd_sc_hd__buf_2 c201 (.A(net183),
    .X(net186));
 sky130_fd_sc_hd__xnor2_4 c202 (.A(net186),
    .B(net183),
    .Y(net187));
 sky130_fd_sc_hd__xnor2_1 c203 (.A(net185),
    .B(net187),
    .Y(net188));
 sky130_fd_sc_hd__xnor2_1 c204 (.A(net43),
    .B(net187),
    .Y(net189));
 sky130_fd_sc_hd__xnor2_1 c205 (.A(net186),
    .B(net183),
    .Y(net190));
 sky130_fd_sc_hd__xnor2_1 c206 (.A(net184),
    .B(net183),
    .Y(net191));
 sky130_fd_sc_hd__buf_1 c207 (.A(net944),
    .X(net192));
 sky130_fd_sc_hd__xnor2_1 c208 (.A(net187),
    .B(net882),
    .Y(net193));
 sky130_fd_sc_hd__clkbuf_1 c209 (.A(net974),
    .X(net194));
 sky130_fd_sc_hd__xnor2_1 c210 (.A(net192),
    .B(net882),
    .Y(net195));
 sky130_fd_sc_hd__a31o_1 c211 (.A1(net187),
    .A2(net193),
    .A3(clknet_1_1__leaf_net42),
    .B1(net183),
    .X(net196));
 sky130_fd_sc_hd__buf_1 c212 (.A(clknet_1_1__leaf_net984),
    .X(net197));
 sky130_fd_sc_hd__a21bo_1 c213 (.A1(net193),
    .A2(clknet_1_0__leaf_net197),
    .B1_N(net979),
    .X(net198));
 sky130_fd_sc_hd__clkbuf_1 c214 (.A(net942),
    .X(net199));
 sky130_fd_sc_hd__a31o_1 c215 (.A1(net194),
    .A2(net186),
    .A3(clknet_1_0__leaf_net197),
    .B1(net183),
    .X(net200));
 sky130_fd_sc_hd__a21bo_1 c216 (.A1(net200),
    .A2(net199),
    .B1_N(clknet_1_1__leaf_net197),
    .X(net201));
 sky130_fd_sc_hd__a41o_1 c217 (.A1(net195),
    .A2(net192),
    .A3(clknet_1_1__leaf_net201),
    .A4(net199),
    .B1(net979),
    .X(net202));
 sky130_fd_sc_hd__clkbuf_1 c218 (.A(net974),
    .X(net203));
 sky130_fd_sc_hd__a41o_1 c219 (.A1(net203),
    .A2(net192),
    .A3(clknet_1_0__leaf_net201),
    .A4(net187),
    .B1(net956),
    .X(net204));
 sky130_fd_sc_hd__buf_1 c220 (.A(clknet_1_1__leaf_net85),
    .X(net205));
 sky130_fd_sc_hd__clkbuf_2 c221 (.A(net771),
    .X(net206));
 sky130_fd_sc_hd__xnor2_1 c222 (.A(net206),
    .B(clknet_1_0__leaf_net205),
    .Y(net207));
 sky130_fd_sc_hd__xnor2_1 c223 (.A(clknet_1_1__leaf_net205),
    .B(net206),
    .Y(net208));
 sky130_fd_sc_hd__buf_1 c224 (.A(clknet_1_1__leaf_net207),
    .X(net209));
 sky130_fd_sc_hd__xnor2_1 c225 (.A(clknet_1_0__leaf_net208),
    .B(net987),
    .Y(net210));
 sky130_fd_sc_hd__xnor2_1 c226 (.A(clknet_1_0__leaf_net205),
    .B(clknet_1_0__leaf_net207),
    .Y(net211));
 sky130_fd_sc_hd__a21bo_1 c227 (.A1(net206),
    .A2(clknet_1_0__leaf_net208),
    .B1_N(clknet_1_0__leaf_net210),
    .X(net212));
 sky130_fd_sc_hd__xnor2_1 c228 (.A(clknet_1_0__leaf_net207),
    .B(net206),
    .Y(net213));
 sky130_fd_sc_hd__buf_1 c229 (.A(net771),
    .X(net214));
 sky130_fd_sc_hd__clkbuf_1 c230 (.A(net778),
    .X(net215));
 sky130_fd_sc_hd__clkbuf_2 c231 (.A(net809),
    .X(net216));
 sky130_fd_sc_hd__xnor2_1 c232 (.A(net215),
    .B(net216),
    .Y(net217));
 sky130_fd_sc_hd__xnor2_1 c233 (.A(net206),
    .B(net214),
    .Y(net218));
 sky130_fd_sc_hd__xnor2_1 c234 (.A(net216),
    .B(net218),
    .Y(net219));
 sky130_fd_sc_hd__xnor2_1 c235 (.A(net217),
    .B(net216),
    .Y(net220));
 sky130_fd_sc_hd__a21bo_1 c236 (.A1(net214),
    .A2(net220),
    .B1_N(net879),
    .X(net221));
 sky130_fd_sc_hd__sdfxtp_1 c237 (.CLK(clknet_4_4_0_clk),
    .D(net218),
    .SCD(net221),
    .SCE(clknet_1_1__leaf_net208),
    .Q(net222));
 sky130_fd_sc_hd__a21bo_1 c238 (.A1(net220),
    .A2(net1042),
    .B1_N(net221),
    .X(net223));
 sky130_fd_sc_hd__a31o_1 c239 (.A1(net209),
    .A2(net222),
    .A3(net221),
    .B1(net220),
    .X(net224));
 sky130_fd_sc_hd__a21bo_1 c240 (.A1(net216),
    .A2(net221),
    .B1_N(net942),
    .X(net225));
 sky130_fd_sc_hd__a31o_1 c241 (.A1(clknet_1_1__leaf_net208),
    .A2(net222),
    .A3(net878),
    .B1(net901),
    .X(net226));
 sky130_fd_sc_hd__buf_4 c242 (.A(net959),
    .X(net227));
 sky130_fd_sc_hd__xnor2_4 c243 (.A(net227),
    .B(net100),
    .Y(net228));
 sky130_fd_sc_hd__xnor2_4 c244 (.A(net227),
    .B(net959),
    .Y(net229));
 sky130_fd_sc_hd__xnor2_1 c245 (.A(net228),
    .B(net229),
    .Y(net230));
 sky130_fd_sc_hd__xnor2_2 c246 (.A(net1068),
    .B(net228),
    .Y(net231));
 sky130_fd_sc_hd__clkbuf_4 c247 (.A(net909),
    .X(net232));
 sky130_fd_sc_hd__buf_1 c248 (.A(net909),
    .X(net233));
 sky130_fd_sc_hd__dlymetal6s2s_1 c249 (.A(net928),
    .X(net234));
 sky130_fd_sc_hd__xnor2_1 c25 (.A(net1008),
    .B(net1006),
    .Y(net0));
 sky130_fd_sc_hd__sdfxtp_1 c250 (.CLK(clknet_4_0_0_clk),
    .D(net230),
    .SCD(net232),
    .SCE(net234),
    .Q(net235));
 sky130_fd_sc_hd__xnor2_1 c251 (.A(net235),
    .B(net233),
    .Y(net236));
 sky130_fd_sc_hd__xnor2_1 c252 (.A(net236),
    .B(net233),
    .Y(net237));
 sky130_fd_sc_hd__a41o_1 c253 (.A1(net103),
    .A2(net1062),
    .A3(net234),
    .A4(net231),
    .B1(net227),
    .X(net238));
 sky130_fd_sc_hd__sdfrtn_1 c254 (.CLK_N(clknet_4_0_0_clk),
    .D(net237),
    .RESET_B(net1047),
    .SCD(net231),
    .SCE(net959),
    .Q(net239));
 sky130_fd_sc_hd__sdfrtp_1 c255 (.CLK(clknet_4_0_0_clk),
    .D(net237),
    .RESET_B(net231),
    .SCD(net232),
    .SCE(net234),
    .Q(net240));
 sky130_fd_sc_hd__a21bo_1 c256 (.A1(net234),
    .A2(net240),
    .B1_N(net236),
    .X(net241));
 sky130_fd_sc_hd__xnor2_1 c257 (.A(net239),
    .B(net227),
    .Y(net242));
 sky130_fd_sc_hd__xnor2_1 c258 (.A(net241),
    .B(net242),
    .Y(net243));
 sky130_fd_sc_hd__xnor2_2 c259 (.A(net101),
    .B(net227),
    .Y(net244));
 sky130_fd_sc_hd__xnor2_1 c26 (.A(net8),
    .B(net1009),
    .Y(net1));
 sky130_fd_sc_hd__a41o_1 c260 (.A1(net244),
    .A2(net232),
    .A3(net228),
    .A4(net229),
    .B1(net243),
    .X(net245));
 sky130_fd_sc_hd__mux4_1 c261 (.A0(net243),
    .A1(net244),
    .A2(net239),
    .A3(net228),
    .S0(net232),
    .S1(net888),
    .X(net246));
 sky130_fd_sc_hd__a41o_1 c262 (.A1(net240),
    .A2(net235),
    .A3(net244),
    .A4(net228),
    .B1(net1061),
    .X(net247));
 sky130_fd_sc_hd__sdfbbn_1 c263 (.CLK_N(clknet_4_2_0_clk),
    .D(net247),
    .RESET_B(net241),
    .SCD(net244),
    .SCE(net889),
    .SET_B(net988),
    .Q(net249),
    .Q_N(net248));
 sky130_fd_sc_hd__buf_1 c264 (.A(net870),
    .X(net250));
 sky130_fd_sc_hd__buf_2 c265 (.A(net250),
    .X(net251));
 sky130_fd_sc_hd__buf_1 c266 (.A(net251),
    .X(net252));
 sky130_fd_sc_hd__buf_2 c267 (.A(net906),
    .X(net253));
 sky130_fd_sc_hd__dlymetal6s2s_1 c268 (.A(net253),
    .X(net254));
 sky130_fd_sc_hd__xnor2_1 c269 (.A(net250),
    .B(net253),
    .Y(net255));
 sky130_fd_sc_hd__xnor2_2 c27 (.A(net759),
    .B(net1006),
    .Y(net2));
 sky130_fd_sc_hd__xnor2_1 c270 (.A(net255),
    .B(net253),
    .Y(net256));
 sky130_fd_sc_hd__clkbuf_1 c271 (.A(net906),
    .X(net257));
 sky130_fd_sc_hd__buf_1 c272 (.A(net257),
    .X(net258));
 sky130_fd_sc_hd__xnor2_1 c273 (.A(net258),
    .B(net251),
    .Y(net259));
 sky130_fd_sc_hd__a21bo_1 c274 (.A1(net253),
    .A2(net251),
    .B1_N(net1001),
    .X(net260));
 sky130_fd_sc_hd__clkbuf_1 c275 (.A(net926),
    .X(net261));
 sky130_fd_sc_hd__xnor2_1 c276 (.A(net251),
    .B(net253),
    .Y(net262));
 sky130_fd_sc_hd__clkbuf_1 c277 (.A(net1049),
    .X(net263));
 sky130_fd_sc_hd__buf_2 c278 (.A(net925),
    .X(net264));
 sky130_fd_sc_hd__buf_1 c279 (.A(clknet_1_0__leaf_net994),
    .X(net265));
 sky130_fd_sc_hd__a21bo_1 c28 (.A1(net1007),
    .A2(net8),
    .B1_N(net1000),
    .X(net3));
 sky130_fd_sc_hd__buf_1 c280 (.A(net925),
    .X(net266));
 sky130_fd_sc_hd__a21bo_1 c281 (.A1(net266),
    .A2(net255),
    .B1_N(net264),
    .X(net267));
 sky130_fd_sc_hd__mux4_1 c282 (.A0(net265),
    .A1(net267),
    .A2(net260),
    .A3(net266),
    .S0(net251),
    .S1(net253),
    .X(net268));
 sky130_fd_sc_hd__a21bo_1 c283 (.A1(net264),
    .A2(net251),
    .B1_N(net946),
    .X(net269));
 sky130_fd_sc_hd__a21bo_1 c284 (.A1(net269),
    .A2(net266),
    .B1_N(net258),
    .X(net270));
 sky130_fd_sc_hd__a21bo_1 c285 (.A1(net250),
    .A2(net262),
    .B1_N(net946),
    .X(net271));
 sky130_fd_sc_hd__xnor2_1 c286 (.A(net264),
    .B(clknet_1_0__leaf_net145),
    .Y(net272));
 sky130_fd_sc_hd__buf_2 c287 (.A(net933),
    .X(net273));
 sky130_fd_sc_hd__xnor2_1 c288 (.A(net273),
    .B(net264),
    .Y(net274));
 sky130_fd_sc_hd__buf_1 c289 (.A(net933),
    .X(net275));
 sky130_fd_sc_hd__xnor2_1 c29 (.A(net2),
    .B(net0),
    .Y(net4));
 sky130_fd_sc_hd__xnor2_2 c290 (.A(net275),
    .B(net273),
    .Y(net276));
 sky130_fd_sc_hd__xnor2_2 c291 (.A(net254),
    .B(net276),
    .Y(net277));
 sky130_fd_sc_hd__dlymetal6s2s_1 c292 (.A(net277),
    .X(net278));
 sky130_fd_sc_hd__clkbuf_2 c293 (.A(net943),
    .X(net279));
 sky130_fd_sc_hd__sdfxtp_1 c294 (.CLK(clknet_4_15_0_clk),
    .D(net273),
    .SCD(net278),
    .SCE(net279),
    .Q(net280));
 sky130_fd_sc_hd__xnor2_1 c295 (.A(net277),
    .B(net273),
    .Y(net281));
 sky130_fd_sc_hd__a21bo_1 c296 (.A1(net276),
    .A2(net277),
    .B1_N(net280),
    .X(net282));
 sky130_fd_sc_hd__xnor2_1 c297 (.A(net280),
    .B(net279),
    .Y(net283));
 sky130_fd_sc_hd__clkbuf_2 c298 (.A(net966),
    .X(net284));
 sky130_fd_sc_hd__clkbuf_1 c299 (.A(net926),
    .X(net285));
 sky130_fd_sc_hd__a21bo_1 c30 (.A1(net1014),
    .A2(net1004),
    .B1_N(net998),
    .X(net5));
 sky130_fd_sc_hd__buf_1 c300 (.A(net941),
    .X(net286));
 sky130_fd_sc_hd__a21bo_1 c301 (.A1(net286),
    .A2(net279),
    .B1_N(net284),
    .X(net287));
 sky130_fd_sc_hd__a41o_1 c302 (.A1(net279),
    .A2(net278),
    .A3(net264),
    .A4(net287),
    .B1(net277),
    .X(net288));
 sky130_fd_sc_hd__a21bo_1 c303 (.A1(net278),
    .A2(net287),
    .B1_N(net284),
    .X(net289));
 sky130_fd_sc_hd__a21bo_1 c304 (.A1(net287),
    .A2(net279),
    .B1_N(net286),
    .X(net290));
 sky130_fd_sc_hd__mux4_1 c305 (.A0(net290),
    .A1(net286),
    .A2(net278),
    .A3(net279),
    .S0(net284),
    .S1(net977),
    .X(net291));
 sky130_fd_sc_hd__a41o_1 c306 (.A1(net285),
    .A2(net280),
    .A3(net290),
    .A4(clknet_1_1__leaf_net272),
    .B1(net977),
    .X(net292));
 sky130_fd_sc_hd__sdfbbn_2 c307 (.CLK_N(clknet_4_12_0_clk),
    .D(net282),
    .RESET_B(net290),
    .SCD(net287),
    .SCE(net279),
    .SET_B(net906),
    .Q(net294),
    .Q_N(net293));
 sky130_fd_sc_hd__clkbuf_4 c308 (.A(net876),
    .X(net295));
 sky130_fd_sc_hd__xnor2_2 c309 (.A(net295),
    .B(net294),
    .Y(net296));
 sky130_fd_sc_hd__xnor2_1 c31 (.A(net5),
    .B(net2),
    .Y(net6));
 sky130_fd_sc_hd__xnor2_4 c310 (.A(net295),
    .B(net293),
    .Y(net297));
 sky130_fd_sc_hd__xnor2_4 c311 (.A(net297),
    .B(net295),
    .Y(net298));
 sky130_fd_sc_hd__buf_1 c312 (.A(net875),
    .X(net299));
 sky130_fd_sc_hd__xnor2_1 c313 (.A(net297),
    .B(net298),
    .Y(net300));
 sky130_fd_sc_hd__xnor2_1 c314 (.A(net296),
    .B(net299),
    .Y(net301));
 sky130_fd_sc_hd__xnor2_4 c315 (.A(net298),
    .B(net956),
    .Y(net302));
 sky130_fd_sc_hd__buf_1 c316 (.A(net916),
    .X(net303));
 sky130_fd_sc_hd__clkbuf_1 c317 (.A(net955),
    .X(net304));
 sky130_fd_sc_hd__buf_1 c318 (.A(net945),
    .X(net305));
 sky130_fd_sc_hd__xnor2_1 c319 (.A(net298),
    .B(net299),
    .Y(net306));
 sky130_fd_sc_hd__a31o_1 c32 (.A1(net4),
    .A2(net6),
    .A3(net3),
    .B1(net1006),
    .X(net7));
 sky130_fd_sc_hd__buf_1 c320 (.A(net966),
    .X(net307));
 sky130_fd_sc_hd__a21bo_1 c321 (.A1(net299),
    .A2(net303),
    .B1_N(net293),
    .X(net308));
 sky130_fd_sc_hd__a21bo_1 c322 (.A1(net308),
    .A2(net296),
    .B1_N(net295),
    .X(net309));
 sky130_fd_sc_hd__mux4_1 c323 (.A0(net303),
    .A1(net296),
    .A2(net308),
    .A3(net307),
    .S0(net302),
    .S1(net305),
    .X(net310));
 sky130_fd_sc_hd__a21bo_1 c324 (.A1(net298),
    .A2(net307),
    .B1_N(net876),
    .X(net311));
 sky130_fd_sc_hd__clkbuf_1 c325 (.A(net973),
    .X(net312));
 sky130_fd_sc_hd__buf_1 c326 (.A(net929),
    .X(net313));
 sky130_fd_sc_hd__mux4_1 c327 (.A0(net304),
    .A1(net309),
    .A2(net308),
    .A3(net313),
    .S0(net297),
    .S1(net302),
    .X(net314));
 sky130_fd_sc_hd__a31o_1 c328 (.A1(net312),
    .A2(net297),
    .A3(net313),
    .B1(net990),
    .X(net315));
 sky130_fd_sc_hd__a31o_1 c329 (.A1(net315),
    .A2(net313),
    .A3(net301),
    .B1(net990),
    .X(net316));
 sky130_fd_sc_hd__xnor2_2 c33 (.A(net1010),
    .B(net1003),
    .Y(net8));
 sky130_fd_sc_hd__buf_1 c330 (.A(clknet_1_1__leaf_net747),
    .X(net317));
 sky130_fd_sc_hd__buf_1 c331 (.A(clknet_1_0__leaf_net747),
    .X(net318));
 sky130_fd_sc_hd__buf_1 c332 (.A(clknet_1_0__leaf_net318),
    .X(net319));
 sky130_fd_sc_hd__xnor2_1 c333 (.A(net319),
    .B(clknet_1_0__leaf_net317),
    .Y(net320));
 sky130_fd_sc_hd__xnor2_1 c334 (.A(clknet_1_0__leaf_net320),
    .B(clknet_1_0__leaf_net317),
    .Y(net321));
 sky130_fd_sc_hd__clkbuf_2 c335 (.A(net908),
    .X(net322));
 sky130_fd_sc_hd__clkbuf_1 c336 (.A(net923),
    .X(net323));
 sky130_fd_sc_hd__xnor2_1 c337 (.A(clknet_1_0__leaf_net317),
    .B(net956),
    .Y(net324));
 sky130_fd_sc_hd__xnor2_1 c338 (.A(clknet_1_1__leaf_net320),
    .B(clknet_1_1__leaf_net318),
    .Y(net325));
 sky130_fd_sc_hd__buf_1 c339 (.A(clknet_1_0__leaf_net950),
    .X(net326));
 sky130_fd_sc_hd__sdfrbp_1 c34 (.CLK(clknet_4_4_0_clk),
    .D(net0),
    .RESET_B(net7),
    .SCD(net2),
    .SCE(net1006),
    .Q(net10),
    .Q_N(net9));
 sky130_fd_sc_hd__xnor2_1 c340 (.A(clknet_1_0__leaf_net324),
    .B(clknet_1_1__leaf_net326),
    .Y(net327));
 sky130_fd_sc_hd__xnor2_1 c341 (.A(net323),
    .B(clknet_1_0__leaf_net326),
    .Y(net328));
 sky130_fd_sc_hd__xnor2_1 c342 (.A(net191),
    .B(clknet_1_1__leaf_net324),
    .Y(net329));
 sky130_fd_sc_hd__a21bo_1 c343 (.A1(clknet_1_0__leaf_net328),
    .A2(clknet_1_0__leaf_net326),
    .B1_N(net322),
    .X(net330));
 sky130_fd_sc_hd__clkbuf_1 c344 (.A(net935),
    .X(net331));
 sky130_fd_sc_hd__xnor2_1 c345 (.A(net322),
    .B(clknet_1_1__leaf_net328),
    .Y(net332));
 sky130_fd_sc_hd__clkbuf_2 c346 (.A(net923),
    .X(net333));
 sky130_fd_sc_hd__clkbuf_1 c347 (.A(net856),
    .X(net334));
 sky130_fd_sc_hd__a31o_1 c348 (.A1(clknet_1_0__leaf_net318),
    .A2(net334),
    .A3(clknet_1_1__leaf_net330),
    .B1(net322),
    .X(net335));
 sky130_fd_sc_hd__a21bo_1 c349 (.A1(net331),
    .A2(net332),
    .B1_N(net333),
    .X(net336));
 sky130_fd_sc_hd__buf_1 c35 (.A(net930),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 c350 (.A(net945),
    .X(net337));
 sky130_fd_sc_hd__a31o_1 c351 (.A1(net335),
    .A2(net337),
    .A3(net333),
    .B1(clknet_1_1__leaf_net324),
    .X(net338));
 sky130_fd_sc_hd__clkbuf_2 c352 (.A(net948),
    .X(net339));
 sky130_fd_sc_hd__buf_2 c353 (.A(net339),
    .X(net340));
 sky130_fd_sc_hd__xnor2_1 c354 (.A(net340),
    .B(net339),
    .Y(net341));
 sky130_fd_sc_hd__buf_2 c355 (.A(net948),
    .X(net342));
 sky130_fd_sc_hd__xnor2_2 c356 (.A(net342),
    .B(net340),
    .Y(net343));
 sky130_fd_sc_hd__xnor2_1 c357 (.A(net340),
    .B(net342),
    .Y(net344));
 sky130_fd_sc_hd__xnor2_2 c358 (.A(net342),
    .B(net343),
    .Y(net345));
 sky130_fd_sc_hd__clkbuf_1 c359 (.A(net827),
    .X(net346));
 sky130_fd_sc_hd__a21bo_1 c36 (.A1(net10),
    .A2(net11),
    .B1_N(net0),
    .X(net12));
 sky130_fd_sc_hd__buf_1 c360 (.A(net967),
    .X(net347));
 sky130_fd_sc_hd__mux4_1 c361 (.A0(net333),
    .A1(net345),
    .A2(net343),
    .A3(net347),
    .S0(net340),
    .S1(net339),
    .X(net348));
 sky130_fd_sc_hd__a21bo_1 c362 (.A1(net347),
    .A2(net344),
    .B1_N(net333),
    .X(net349));
 sky130_fd_sc_hd__xnor2_1 c363 (.A(net341),
    .B(net342),
    .Y(net350));
 sky130_fd_sc_hd__a41o_1 c364 (.A1(net350),
    .A2(net344),
    .A3(net342),
    .A4(net346),
    .B1(net339),
    .X(net351));
 sky130_fd_sc_hd__buf_1 c365 (.A(clknet_1_1__leaf_net951),
    .X(net352));
 sky130_fd_sc_hd__xnor2_1 c366 (.A(net344),
    .B(clknet_1_0__leaf_net352),
    .Y(net353));
 sky130_fd_sc_hd__xnor2_1 c367 (.A(clknet_1_0__leaf_net352),
    .B(net983),
    .Y(net354));
 sky130_fd_sc_hd__a31o_1 c368 (.A1(net316),
    .A2(clknet_1_1__leaf_net352),
    .A3(clknet_1_1__leaf_net353),
    .B1(net345),
    .X(net355));
 sky130_fd_sc_hd__xnor2_1 c369 (.A(net983),
    .B(clknet_1_0__leaf_net984),
    .Y(net356));
 sky130_fd_sc_hd__a21bo_4 c37 (.A1(net1),
    .A2(net10),
    .B1_N(net1006),
    .X(net13));
 sky130_fd_sc_hd__xnor2_1 c370 (.A(net356),
    .B(net340),
    .Y(net357));
 sky130_fd_sc_hd__xnor2_1 c371 (.A(net354),
    .B(clknet_1_0__leaf_net357),
    .Y(net358));
 sky130_fd_sc_hd__buf_1 c372 (.A(clknet_1_0__leaf_net984),
    .X(net359));
 sky130_fd_sc_hd__dlymetal6s2s_1 c373 (.A(net778),
    .X(net360));
 sky130_fd_sc_hd__xnor2_1 c374 (.A(net228),
    .B(net989),
    .Y(net361));
 sky130_fd_sc_hd__clkbuf_4 c375 (.A(net229),
    .X(net362));
 sky130_fd_sc_hd__xnor2_1 c376 (.A(net339),
    .B(net232),
    .Y(net363));
 sky130_fd_sc_hd__clkbuf_1 c377 (.A(net761),
    .X(net364));
 sky130_fd_sc_hd__xnor2_4 c378 (.A(net232),
    .B(net229),
    .Y(net365));
 sky130_fd_sc_hd__buf_2 c379 (.A(net761),
    .X(net366));
 sky130_fd_sc_hd__a31o_1 c38 (.A1(net12),
    .A2(net6),
    .A3(net11),
    .B1(net13),
    .X(net14));
 sky130_fd_sc_hd__buf_1 c380 (.A(clknet_1_1__leaf_net950),
    .X(net367));
 sky130_fd_sc_hd__xnor2_1 c381 (.A(net363),
    .B(net229),
    .Y(net368));
 sky130_fd_sc_hd__clkbuf_1 c382 (.A(net980),
    .X(net369));
 sky130_fd_sc_hd__a21bo_1 c383 (.A1(net362),
    .A2(net361),
    .B1_N(net364),
    .X(net370));
 sky130_fd_sc_hd__buf_1 c384 (.A(net983),
    .X(net371));
 sky130_fd_sc_hd__a31o_1 c385 (.A1(net361),
    .A2(net365),
    .A3(net362),
    .B1(net366),
    .X(net372));
 sky130_fd_sc_hd__xnor2_4 c386 (.A(net366),
    .B(net945),
    .Y(net373));
 sky130_fd_sc_hd__xnor2_2 c387 (.A(net371),
    .B(net373),
    .Y(net374));
 sky130_fd_sc_hd__buf_1 c388 (.A(clknet_1_1__leaf_net985),
    .X(net375));
 sky130_fd_sc_hd__clkbuf_1 c389 (.A(net827),
    .X(net376));
 sky130_fd_sc_hd__buf_1 c39 (.A(net930),
    .X(net15));
 sky130_fd_sc_hd__xnor2_1 c390 (.A(net373),
    .B(net931),
    .Y(net377));
 sky130_fd_sc_hd__xnor2_2 c391 (.A(net373),
    .B(net374),
    .Y(net378));
 sky130_fd_sc_hd__a41o_1 c392 (.A1(net374),
    .A2(net377),
    .A3(net378),
    .A4(net362),
    .B1(net373),
    .X(net379));
 sky130_fd_sc_hd__buf_1 c393 (.A(net940),
    .X(net380));
 sky130_fd_sc_hd__dfbbn_2 c394 (.CLK_N(clknet_4_3_0_clk),
    .D(net364),
    .RESET_B(net380),
    .SET_B(net378),
    .Q(net382),
    .Q_N(net381));
 sky130_fd_sc_hd__mux4_1 c395 (.A0(net375),
    .A1(net380),
    .A2(net377),
    .A3(net382),
    .S0(net378),
    .S1(net362),
    .X(net383));
 sky130_fd_sc_hd__buf_2 c396 (.A(net264),
    .X(net384));
 sky130_fd_sc_hd__buf_1 c397 (.A(net384),
    .X(net385));
 sky130_fd_sc_hd__clkbuf_1 c398 (.A(net385),
    .X(net386));
 sky130_fd_sc_hd__buf_1 c399 (.A(net756),
    .X(net387));
 sky130_fd_sc_hd__a41o_1 c40 (.A1(net7),
    .A2(net628),
    .A3(net15),
    .A4(net12),
    .B1(net1044),
    .X(net16));
 sky130_fd_sc_hd__buf_1 c400 (.A(net756),
    .X(net388));
 sky130_fd_sc_hd__xnor2_1 c401 (.A(net385),
    .B(net388),
    .Y(net389));
 sky130_fd_sc_hd__buf_1 c402 (.A(net781),
    .X(net390));
 sky130_fd_sc_hd__xnor2_1 c403 (.A(net384),
    .B(net387),
    .Y(net391));
 sky130_fd_sc_hd__xnor2_2 c404 (.A(net387),
    .B(net384),
    .Y(net392));
 sky130_fd_sc_hd__clkbuf_1 c405 (.A(net392),
    .X(net393));
 sky130_fd_sc_hd__clkbuf_1 c406 (.A(net902),
    .X(net394));
 sky130_fd_sc_hd__clkbuf_1 c407 (.A(net937),
    .X(net395));
 sky130_fd_sc_hd__buf_1 c408 (.A(net1033),
    .X(net396));
 sky130_fd_sc_hd__xnor2_1 c409 (.A(net391),
    .B(net396),
    .Y(net397));
 sky130_fd_sc_hd__mux4_1 c41 (.A0(net15),
    .A1(net12),
    .A2(net9),
    .A3(net13),
    .S0(net1007),
    .S1(net929),
    .X(net17));
 sky130_fd_sc_hd__buf_1 c410 (.A(net937),
    .X(net398));
 sky130_fd_sc_hd__xnor2_1 c411 (.A(net390),
    .B(net398),
    .Y(net399));
 sky130_fd_sc_hd__clkbuf_1 c412 (.A(net936),
    .X(net400));
 sky130_fd_sc_hd__a21bo_1 c413 (.A1(net396),
    .A2(net399),
    .B1_N(net388),
    .X(net401));
 sky130_fd_sc_hd__clkbuf_1 c414 (.A(net936),
    .X(net402));
 sky130_fd_sc_hd__a21bo_1 c415 (.A1(net397),
    .A2(net400),
    .B1_N(net392),
    .X(net403));
 sky130_fd_sc_hd__a21bo_2 c416 (.A1(net388),
    .A2(net400),
    .B1_N(net871),
    .X(net404));
 sky130_fd_sc_hd__a21bo_1 c417 (.A1(net391),
    .A2(net401),
    .B1_N(net399),
    .X(net405));
 sky130_fd_sc_hd__clkbuf_2 c418 (.A(net294),
    .X(net406));
 sky130_fd_sc_hd__clkbuf_4 c419 (.A(net406),
    .X(net407));
 sky130_fd_sc_hd__a41o_1 c42 (.A1(net8),
    .A2(net13),
    .A3(net1006),
    .A4(net929),
    .B1(net1044),
    .X(net18));
 sky130_fd_sc_hd__xnor2_1 c420 (.A(net407),
    .B(net406),
    .Y(net408));
 sky130_fd_sc_hd__xnor2_1 c421 (.A(net404),
    .B(net407),
    .Y(net409));
 sky130_fd_sc_hd__xnor2_1 c422 (.A(net284),
    .B(net407),
    .Y(net410));
 sky130_fd_sc_hd__xnor2_1 c423 (.A(net402),
    .B(net406),
    .Y(net411));
 sky130_fd_sc_hd__clkbuf_2 c424 (.A(net773),
    .X(net412));
 sky130_fd_sc_hd__xnor2_1 c425 (.A(net1032),
    .B(net407),
    .Y(net413));
 sky130_fd_sc_hd__xnor2_4 c426 (.A(net412),
    .B(net1032),
    .Y(net414));
 sky130_fd_sc_hd__clkbuf_1 c427 (.A(net773),
    .X(net415));
 sky130_fd_sc_hd__buf_1 c428 (.A(net935),
    .X(net416));
 sky130_fd_sc_hd__a31o_1 c429 (.A1(net413),
    .A2(net407),
    .A3(net1032),
    .B1(net416),
    .X(net417));
 sky130_fd_sc_hd__a21bo_1 c43 (.A1(net3),
    .A2(net15),
    .B1_N(net954),
    .X(net19));
 sky130_fd_sc_hd__buf_1 c430 (.A(net981),
    .X(net418));
 sky130_fd_sc_hd__xnor2_1 c431 (.A(net407),
    .B(net960),
    .Y(net419));
 sky130_fd_sc_hd__xnor2_1 c432 (.A(net418),
    .B(net411),
    .Y(net420));
 sky130_fd_sc_hd__xnor2_1 c433 (.A(net416),
    .B(net1032),
    .Y(net421));
 sky130_fd_sc_hd__buf_1 c434 (.A(net1043),
    .X(net422));
 sky130_fd_sc_hd__a21bo_1 c435 (.A1(net422),
    .A2(net1032),
    .B1_N(net407),
    .X(net423));
 sky130_fd_sc_hd__clkbuf_4 c436 (.A(net908),
    .X(net424));
 sky130_fd_sc_hd__clkbuf_1 c437 (.A(net807),
    .X(net425));
 sky130_fd_sc_hd__mux4_1 c438 (.A0(net425),
    .A1(net1032),
    .A2(net423),
    .A3(net407),
    .S0(net424),
    .S1(net421),
    .X(net426));
 sky130_fd_sc_hd__mux4_1 c439 (.A0(net423),
    .A1(net414),
    .A2(net425),
    .A3(net420),
    .S0(net424),
    .S1(net960),
    .X(net427));
 sky130_fd_sc_hd__buf_1 c44 (.A(clknet_1_0__leaf_net42),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_2 c440 (.A(net991),
    .X(net428));
 sky130_fd_sc_hd__xnor2_1 c441 (.A(net428),
    .B(net990),
    .Y(net429));
 sky130_fd_sc_hd__clkbuf_2 c442 (.A(net428),
    .X(net430));
 sky130_fd_sc_hd__xnor2_1 c443 (.A(net428),
    .B(net429),
    .Y(net431));
 sky130_fd_sc_hd__clkbuf_2 c444 (.A(net934),
    .X(net432));
 sky130_fd_sc_hd__clkbuf_1 c445 (.A(net934),
    .X(net433));
 sky130_fd_sc_hd__xnor2_4 c446 (.A(net432),
    .B(net430),
    .Y(net434));
 sky130_fd_sc_hd__buf_1 c447 (.A(net1065),
    .X(net435));
 sky130_fd_sc_hd__clkbuf_2 c448 (.A(net922),
    .X(net436));
 sky130_fd_sc_hd__buf_1 c449 (.A(net871),
    .X(net437));
 sky130_fd_sc_hd__xnor2_1 c45 (.A(clknet_1_0__leaf_net20),
    .B(clknet_1_0__leaf_net42),
    .Y(net21));
 sky130_fd_sc_hd__a21bo_1 c450 (.A1(net437),
    .A2(net431),
    .B1_N(net428),
    .X(net438));
 sky130_fd_sc_hd__xnor2_1 c451 (.A(net429),
    .B(net437),
    .Y(net439));
 sky130_fd_sc_hd__clkbuf_2 c452 (.A(net958),
    .X(net440));
 sky130_fd_sc_hd__buf_1 c453 (.A(clknet_1_0__leaf_net949),
    .X(net441));
 sky130_fd_sc_hd__a21bo_1 c454 (.A1(net441),
    .A2(net440),
    .B1_N(net436),
    .X(net442));
 sky130_fd_sc_hd__xnor2_1 c455 (.A(clknet_1_1__leaf_net442),
    .B(net440),
    .Y(net443));
 sky130_fd_sc_hd__a21bo_1 c456 (.A1(net436),
    .A2(net440),
    .B1_N(clknet_1_0__leaf_net442),
    .X(net444));
 sky130_fd_sc_hd__dfbbn_1 c457 (.CLK_N(clknet_4_9_0_clk),
    .D(net430),
    .RESET_B(net431),
    .SET_B(clknet_1_0__leaf_net442),
    .Q(net446),
    .Q_N(net445));
 sky130_fd_sc_hd__a21bo_1 c458 (.A1(net444),
    .A2(clknet_1_1__leaf_net442),
    .B1_N(net446),
    .X(net447));
 sky130_fd_sc_hd__a21bo_1 c459 (.A1(net446),
    .A2(net436),
    .B1_N(net440),
    .X(net448));
 sky130_fd_sc_hd__buf_1 c46 (.A(clknet_1_0__leaf_net951),
    .X(net22));
 sky130_fd_sc_hd__a41o_1 c460 (.A1(clknet_1_1__leaf_net447),
    .A2(net448),
    .A3(clknet_1_1__leaf_net442),
    .A4(net436),
    .B1(net445),
    .X(net449));
 sky130_fd_sc_hd__mux4_1 c461 (.A0(net443),
    .A1(net431),
    .A2(clknet_1_0__leaf_net447),
    .A3(net434),
    .S0(net436),
    .S1(net957),
    .X(net450));
 sky130_fd_sc_hd__buf_2 c462 (.A(net856),
    .X(net451));
 sky130_fd_sc_hd__buf_1 c463 (.A(net451),
    .X(net452));
 sky130_fd_sc_hd__xnor2_1 c464 (.A(net452),
    .B(net451),
    .Y(net453));
 sky130_fd_sc_hd__clkbuf_2 c465 (.A(net760),
    .X(net454));
 sky130_fd_sc_hd__buf_4 c466 (.A(net760),
    .X(net455));
 sky130_fd_sc_hd__a21bo_1 c467 (.A1(net440),
    .A2(net455),
    .B1_N(net451),
    .X(net456));
 sky130_fd_sc_hd__clkbuf_1 c468 (.A(net922),
    .X(net457));
 sky130_fd_sc_hd__xnor2_1 c469 (.A(net455),
    .B(net451),
    .Y(net458));
 sky130_fd_sc_hd__xnor2_1 c47 (.A(net1013),
    .B(clknet_1_0__leaf_net20),
    .Y(net23));
 sky130_fd_sc_hd__xnor2_1 c470 (.A(net452),
    .B(net957),
    .Y(net459));
 sky130_fd_sc_hd__xnor2_4 c471 (.A(net455),
    .B(net454),
    .Y(net460));
 sky130_fd_sc_hd__xnor2_2 c472 (.A(net458),
    .B(net460),
    .Y(net461));
 sky130_fd_sc_hd__a41o_1 c473 (.A1(net456),
    .A2(net457),
    .A3(net461),
    .A4(net454),
    .B1(net451),
    .X(net462));
 sky130_fd_sc_hd__buf_1 c474 (.A(net917),
    .X(net463));
 sky130_fd_sc_hd__mux4_1 c475 (.A0(net452),
    .A1(net455),
    .A2(net461),
    .A3(net460),
    .S0(net333),
    .S1(net451),
    .X(net464));
 sky130_fd_sc_hd__buf_1 c476 (.A(net944),
    .X(net465));
 sky130_fd_sc_hd__xnor2_1 c477 (.A(net465),
    .B(net965),
    .Y(net466));
 sky130_fd_sc_hd__a41o_1 c478 (.A1(net457),
    .A2(net455),
    .A3(net463),
    .A4(net456),
    .B1(net460),
    .X(net467));
 sky130_fd_sc_hd__xnor2_1 c479 (.A(net463),
    .B(net455),
    .Y(net468));
 sky130_fd_sc_hd__xnor2_1 c48 (.A(clknet_1_1__leaf_net22),
    .B(clknet_1_1__leaf_net21),
    .Y(net24));
 sky130_fd_sc_hd__mux4_1 c480 (.A0(net468),
    .A1(net463),
    .A2(net461),
    .A3(net456),
    .S0(net460),
    .S1(net455),
    .X(net469));
 sky130_fd_sc_hd__xnor2_1 c481 (.A(net466),
    .B(net939),
    .Y(net470));
 sky130_fd_sc_hd__a21bo_1 c482 (.A1(net454),
    .A2(net470),
    .B1_N(net460),
    .X(net471));
 sky130_fd_sc_hd__a41o_1 c483 (.A1(net465),
    .A2(net470),
    .A3(net471),
    .A4(net467),
    .B1(net455),
    .X(net472));
 sky130_fd_sc_hd__buf_2 c484 (.A(net360),
    .X(net473));
 sky130_fd_sc_hd__buf_1 c485 (.A(net473),
    .X(net474));
 sky130_fd_sc_hd__xnor2_1 c486 (.A(net474),
    .B(net360),
    .Y(net475));
 sky130_fd_sc_hd__clkbuf_2 c487 (.A(net473),
    .X(net476));
 sky130_fd_sc_hd__xnor2_1 c488 (.A(net476),
    .B(net473),
    .Y(net477));
 sky130_fd_sc_hd__xnor2_2 c489 (.A(net473),
    .B(net476),
    .Y(net478));
 sky130_fd_sc_hd__xnor2_1 c49 (.A(clknet_1_0__leaf_net20),
    .B(clknet_1_0__leaf_net23),
    .Y(net25));
 sky130_fd_sc_hd__buf_1 c490 (.A(clknet_1_0__leaf_net764),
    .X(net479));
 sky130_fd_sc_hd__buf_1 c491 (.A(clknet_1_1__leaf_net764),
    .X(net480));
 sky130_fd_sc_hd__buf_4 c492 (.A(net966),
    .X(net481));
 sky130_fd_sc_hd__a21bo_1 c493 (.A1(net480),
    .A2(net481),
    .B1_N(net476),
    .X(net482));
 sky130_fd_sc_hd__dfbbp_1 c494 (.CLK(clknet_4_6_0_clk),
    .D(net475),
    .RESET_B(clknet_1_0__leaf_net479),
    .SET_B(net473),
    .Q(net484),
    .Q_N(net483));
 sky130_fd_sc_hd__a21bo_1 c495 (.A1(clknet_1_0__leaf_net482),
    .A2(net481),
    .B1_N(net474),
    .X(net485));
 sky130_fd_sc_hd__buf_1 c496 (.A(net967),
    .X(net486));
 sky130_fd_sc_hd__buf_1 c497 (.A(net966),
    .X(net487));
 sky130_fd_sc_hd__buf_1 c498 (.A(net917),
    .X(net488));
 sky130_fd_sc_hd__clkbuf_1 c499 (.A(net923),
    .X(net489));
 sky130_fd_sc_hd__xnor2_1 c50 (.A(clknet_1_0__leaf_net42),
    .B(clknet_1_0__leaf_net20),
    .Y(net26));
 sky130_fd_sc_hd__a31o_1 c500 (.A1(net489),
    .A2(net484),
    .A3(net360),
    .B1(net488),
    .X(net490));
 sky130_fd_sc_hd__a21bo_1 c501 (.A1(clknet_1_1__leaf_net479),
    .A2(net487),
    .B1_N(net490),
    .X(net491));
 sky130_fd_sc_hd__a21bo_1 c502 (.A1(net467),
    .A2(net487),
    .B1_N(clknet_1_1__leaf_net482),
    .X(net492));
 sky130_fd_sc_hd__a31o_1 c503 (.A1(clknet_1_0__leaf_net491),
    .A2(net486),
    .A3(net481),
    .B1(net943),
    .X(net493));
 sky130_fd_sc_hd__a31o_1 c504 (.A1(net490),
    .A2(clknet_1_0__leaf_net493),
    .A3(net488),
    .B1(net473),
    .X(net494));
 sky130_fd_sc_hd__a21bo_1 c505 (.A1(net487),
    .A2(clknet_1_1__leaf_net493),
    .B1_N(net490),
    .X(net495));
 sky130_fd_sc_hd__xnor2_1 c506 (.A(clknet_1_1__leaf_net491),
    .B(net481),
    .Y(net496));
 sky130_fd_sc_hd__xnor2_2 c507 (.A(net481),
    .B(net381),
    .Y(net497));
 sky130_fd_sc_hd__xnor2_1 c508 (.A(net481),
    .B(clknet_1_1__leaf_net984),
    .Y(net498));
 sky130_fd_sc_hd__clkbuf_1 c509 (.A(net751),
    .X(net499));
 sky130_fd_sc_hd__buf_1 c51 (.A(clknet_1_0__leaf_net951),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_4 c510 (.A(net751),
    .X(net500));
 sky130_fd_sc_hd__xnor2_4 c511 (.A(net382),
    .B(net500),
    .Y(net501));
 sky130_fd_sc_hd__a21bo_1 c512 (.A1(net376),
    .A2(clknet_1_0__leaf_net498),
    .B1_N(net501),
    .X(net502));
 sky130_fd_sc_hd__a21bo_1 c513 (.A1(clknet_1_1__leaf_net498),
    .A2(net382),
    .B1_N(net942),
    .X(net503));
 sky130_fd_sc_hd__xnor2_1 c514 (.A(net501),
    .B(net481),
    .Y(net1026));
 sky130_fd_sc_hd__xnor2_4 c515 (.A(net500),
    .B(net501),
    .Y(net504));
 sky130_fd_sc_hd__a21bo_1 c516 (.A1(net504),
    .A2(clknet_1_0__leaf_net496),
    .B1_N(net501),
    .X(net505));
 sky130_fd_sc_hd__xnor2_1 c517 (.A(net502),
    .B(net499),
    .Y(net506));
 sky130_fd_sc_hd__sdfxbp_1 c518 (.CLK(clknet_4_12_0_clk),
    .D(clknet_1_1__leaf_net498),
    .SCD(net500),
    .SCE(clknet_1_1__leaf_net496),
    .Q(net508),
    .Q_N(net507));
 sky130_fd_sc_hd__xnor2_4 c519 (.A(net497),
    .B(net504),
    .Y(net509));
 sky130_fd_sc_hd__a31o_1 c52 (.A1(clknet_1_0__leaf_net24),
    .A2(clknet_1_0__leaf_net22),
    .A3(clknet_1_0__leaf_net27),
    .B1(clknet_1_1__leaf_net20),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_2 c520 (.A(net973),
    .X(net510));
 sky130_fd_sc_hd__a21bo_1 c521 (.A1(net509),
    .A2(net508),
    .B1_N(net510),
    .X(net511));
 sky130_fd_sc_hd__a21bo_1 c522 (.A1(net503),
    .A2(net507),
    .B1_N(net509),
    .X(net512));
 sky130_fd_sc_hd__a21bo_1 c523 (.A1(net500),
    .A2(net509),
    .B1_N(net965),
    .X(net513));
 sky130_fd_sc_hd__a21bo_1 c524 (.A1(net506),
    .A2(net510),
    .B1_N(net504),
    .X(net514));
 sky130_fd_sc_hd__a31o_1 c525 (.A1(net501),
    .A2(net509),
    .A3(net481),
    .B1(net1071),
    .X(net515));
 sky130_fd_sc_hd__clkbuf_1 c526 (.A(net944),
    .X(net516));
 sky130_fd_sc_hd__a21bo_1 c527 (.A1(net508),
    .A2(net516),
    .B1_N(net510),
    .X(net517));
 sky130_fd_sc_hd__buf_4 c528 (.A(net753),
    .X(net518));
 sky130_fd_sc_hd__buf_2 c529 (.A(net518),
    .X(net519));
 sky130_fd_sc_hd__a21bo_1 c53 (.A1(clknet_1_1__leaf_net23),
    .A2(clknet_1_1__leaf_net22),
    .B1_N(clknet_1_0__leaf_net42),
    .X(net29));
 sky130_fd_sc_hd__xnor2_2 c530 (.A(net519),
    .B(net518),
    .Y(net520));
 sky130_fd_sc_hd__xnor2_4 c531 (.A(net519),
    .B(net518),
    .Y(net521));
 sky130_fd_sc_hd__a21bo_1 c532 (.A1(net521),
    .A2(net519),
    .B1_N(net518),
    .X(net522));
 sky130_fd_sc_hd__buf_1 c533 (.A(net752),
    .X(net523));
 sky130_fd_sc_hd__xnor2_2 c534 (.A(net520),
    .B(net521),
    .Y(net524));
 sky130_fd_sc_hd__buf_2 c535 (.A(net793),
    .X(net525));
 sky130_fd_sc_hd__xnor2_4 c536 (.A(net1066),
    .B(net521),
    .Y(net526));
 sky130_fd_sc_hd__buf_1 c537 (.A(net787),
    .X(net527));
 sky130_fd_sc_hd__sdfxbp_1 c538 (.CLK(clknet_4_10_0_clk),
    .D(net524),
    .SCD(net527),
    .SCE(net526),
    .Q(net529),
    .Q_N(net528));
 sky130_fd_sc_hd__sdfxtp_1 c539 (.CLK(clknet_4_10_0_clk),
    .D(net521),
    .SCD(net525),
    .SCE(net526),
    .Q(net530));
 sky130_fd_sc_hd__buf_1 c54 (.A(net923),
    .X(net30));
 sky130_fd_sc_hd__a21bo_1 c540 (.A1(net518),
    .A2(net527),
    .B1_N(net525),
    .X(net531));
 sky130_fd_sc_hd__a21bo_1 c541 (.A1(net523),
    .A2(net1037),
    .B1_N(net531),
    .X(net532));
 sky130_fd_sc_hd__a21bo_1 c542 (.A1(net529),
    .A2(net1037),
    .B1_N(net520),
    .X(net533));
 sky130_fd_sc_hd__mux4_1 c543 (.A0(net526),
    .A1(net532),
    .A2(net524),
    .A3(net533),
    .S0(net530),
    .S1(net518),
    .X(net534));
 sky130_fd_sc_hd__a21bo_1 c544 (.A1(net533),
    .A2(net525),
    .B1_N(net529),
    .X(net535));
 sky130_fd_sc_hd__a21bo_1 c545 (.A1(net1037),
    .A2(net533),
    .B1_N(net532),
    .X(net536));
 sky130_fd_sc_hd__a41o_1 c546 (.A1(net533),
    .A2(net532),
    .A3(net885),
    .A4(clknet_1_0__leaf_net914),
    .B1(net924),
    .X(net537));
 sky130_fd_sc_hd__a21bo_1 c547 (.A1(net531),
    .A2(net532),
    .B1_N(net952),
    .X(net538));
 sky130_fd_sc_hd__mux4_1 c548 (.A0(net532),
    .A1(net538),
    .A2(net528),
    .A3(net526),
    .S0(net527),
    .S1(net924),
    .X(net539));
 sky130_fd_sc_hd__sdfbbp_1 c549 (.CLK(clknet_4_10_0_clk),
    .D(net538),
    .RESET_B(net526),
    .SCD(net884),
    .SCE(clknet_1_0__leaf_net914),
    .SET_B(net1048),
    .Q(net541),
    .Q_N(net540));
 sky130_fd_sc_hd__clkbuf_1 c55 (.A(net981),
    .X(net31));
 sky130_fd_sc_hd__xnor2_1 c550 (.A(net424),
    .B(net991),
    .Y(net542));
 sky130_fd_sc_hd__buf_1 c551 (.A(net542),
    .X(net543));
 sky130_fd_sc_hd__clkbuf_1 c552 (.A(net543),
    .X(net544));
 sky130_fd_sc_hd__clkbuf_1 c553 (.A(net543),
    .X(net545));
 sky130_fd_sc_hd__buf_1 c554 (.A(net972),
    .X(net546));
 sky130_fd_sc_hd__xnor2_1 c555 (.A(net542),
    .B(net525),
    .Y(net547));
 sky130_fd_sc_hd__buf_1 c556 (.A(net525),
    .X(net548));
 sky130_fd_sc_hd__clkbuf_2 c557 (.A(net972),
    .X(net549));
 sky130_fd_sc_hd__xnor2_1 c558 (.A(net547),
    .B(net549),
    .Y(net550));
 sky130_fd_sc_hd__xnor2_1 c559 (.A(net549),
    .B(net546),
    .Y(net551));
 sky130_fd_sc_hd__a41o_1 c56 (.A1(net31),
    .A2(clknet_1_0__leaf_net29),
    .A3(net30),
    .A4(net1006),
    .B1(clknet_1_1__leaf_net20),
    .X(net32));
 sky130_fd_sc_hd__xnor2_1 c560 (.A(net551),
    .B(net549),
    .Y(net552));
 sky130_fd_sc_hd__a21bo_1 c561 (.A1(net548),
    .A2(net552),
    .B1_N(net549),
    .X(net553));
 sky130_fd_sc_hd__xnor2_1 c562 (.A(net546),
    .B(net548),
    .Y(net554));
 sky130_fd_sc_hd__a21bo_1 c563 (.A1(net1056),
    .A2(net552),
    .B1_N(net404),
    .X(net555));
 sky130_fd_sc_hd__a21bo_1 c564 (.A1(net553),
    .A2(net525),
    .X(net873));
 sky130_fd_sc_hd__a21bo_1 c565 (.A1(net545),
    .A2(net549),
    .B1_N(net553),
    .X(net557));
 sky130_fd_sc_hd__buf_1 c566 (.A(clknet_1_1__leaf_net994),
    .X(net558));
 sky130_fd_sc_hd__xnor2_1 c567 (.A(clknet_1_1__leaf_net558),
    .B(net549),
    .Y(net559));
 sky130_fd_sc_hd__a21bo_1 c568 (.A1(net553),
    .A2(clknet_1_0__leaf_net558),
    .B1_N(net424),
    .X(net560));
 sky130_fd_sc_hd__xnor2_1 c569 (.A(net559),
    .B(net921),
    .Y(net561));
 sky130_fd_sc_hd__buf_6 c57 (.A(net902),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_1 c570 (.A(net921),
    .X(net562));
 sky130_fd_sc_hd__a21bo_1 c571 (.A1(net561),
    .A2(net562),
    .B1_N(net873),
    .X(net563));
 sky130_fd_sc_hd__buf_2 c572 (.A(net775),
    .X(net564));
 sky130_fd_sc_hd__xnor2_1 c573 (.A(net564),
    .B(net970),
    .Y(net565));
 sky130_fd_sc_hd__clkbuf_2 c574 (.A(net775),
    .X(net566));
 sky130_fd_sc_hd__clkbuf_1 c575 (.A(net566),
    .X(net567));
 sky130_fd_sc_hd__clkbuf_1 c576 (.A(net919),
    .X(net568));
 sky130_fd_sc_hd__xnor2_1 c577 (.A(net567),
    .B(net566),
    .Y(net569));
 sky130_fd_sc_hd__xnor2_1 c578 (.A(net568),
    .B(net564),
    .Y(net570));
 sky130_fd_sc_hd__buf_1 c579 (.A(net448),
    .X(net571));
 sky130_fd_sc_hd__a21bo_1 c58 (.A1(net33),
    .A2(clknet_1_0__leaf_net27),
    .B1_N(clknet_1_0__leaf_net23),
    .X(net34));
 sky130_fd_sc_hd__a21bo_1 c580 (.A1(net564),
    .A2(net571),
    .B1_N(net567),
    .X(net572));
 sky130_fd_sc_hd__clkbuf_1 c581 (.A(net978),
    .X(net573));
 sky130_fd_sc_hd__clkbuf_1 c582 (.A(net964),
    .X(net574));
 sky130_fd_sc_hd__a21bo_1 c583 (.A1(net571),
    .A2(net570),
    .B1_N(net564),
    .X(net575));
 sky130_fd_sc_hd__a21bo_1 c584 (.A1(net574),
    .A2(net566),
    .B1_N(net573),
    .X(net576));
 sky130_fd_sc_hd__xnor2_1 c585 (.A(net576),
    .B(net571),
    .Y(net577));
 sky130_fd_sc_hd__clkbuf_1 c586 (.A(net943),
    .X(net578));
 sky130_fd_sc_hd__a21bo_1 c587 (.A1(net573),
    .A2(net578),
    .B1_N(net574),
    .X(net579));
 sky130_fd_sc_hd__a21bo_1 c588 (.A1(net569),
    .A2(net570),
    .B1_N(net565),
    .X(net580));
 sky130_fd_sc_hd__a21bo_1 c589 (.A1(net580),
    .A2(net576),
    .B1_N(net577),
    .X(net581));
 sky130_fd_sc_hd__sdfbbn_1 c59 (.CLK_N(clknet_4_1_0_clk),
    .D(clknet_1_0__leaf_net26),
    .RESET_B(clknet_1_0__leaf_net34),
    .SCD(net13),
    .SCE(clknet_1_1__leaf_net27),
    .SET_B(clknet_1_0__leaf_net912),
    .Q(net36),
    .Q_N(net35));
 sky130_fd_sc_hd__a21bo_1 c590 (.A1(net1063),
    .A2(net580),
    .B1_N(net576),
    .X(net582));
 sky130_fd_sc_hd__a41o_1 c591 (.A1(net579),
    .A2(net572),
    .A3(net564),
    .A4(net566),
    .B1(net883),
    .X(net583));
 sky130_fd_sc_hd__a41o_1 c592 (.A1(net580),
    .A2(net576),
    .A3(net564),
    .A4(net883),
    .B1(net975),
    .X(net584));
 sky130_fd_sc_hd__xnor2_1 c593 (.A(net975),
    .B(net978),
    .Y(net585));
 sky130_fd_sc_hd__buf_2 c594 (.A(net939),
    .X(net586));
 sky130_fd_sc_hd__clkbuf_2 c595 (.A(net586),
    .X(net587));
 sky130_fd_sc_hd__buf_1 c596 (.A(net586),
    .X(net588));
 sky130_fd_sc_hd__xnor2_2 c597 (.A(net587),
    .B(net586),
    .Y(net589));
 sky130_fd_sc_hd__xnor2_1 c598 (.A(net587),
    .B(net586),
    .Y(net590));
 sky130_fd_sc_hd__buf_1 c599 (.A(net908),
    .X(net591));
 sky130_fd_sc_hd__a21bo_1 c60 (.A1(net30),
    .A2(clknet_1_1__leaf_net27),
    .B1_N(net35),
    .X(net37));
 sky130_fd_sc_hd__xnor2_1 c600 (.A(net460),
    .B(net588),
    .Y(net592));
 sky130_fd_sc_hd__sdfxtp_1 c601 (.CLK(clknet_4_13_0_clk),
    .D(net592),
    .SCD(net589),
    .SCE(net586),
    .Q(net593));
 sky130_fd_sc_hd__dlymetal6s2s_1 c602 (.A(net908),
    .X(net594));
 sky130_fd_sc_hd__a21bo_1 c603 (.A1(net588),
    .A2(net589),
    .B1_N(net594),
    .X(net595));
 sky130_fd_sc_hd__a21bo_1 c604 (.A1(net593),
    .A2(net594),
    .B1_N(net892),
    .X(net596));
 sky130_fd_sc_hd__xnor2_1 c605 (.A(net591),
    .B(net593),
    .Y(net597));
 sky130_fd_sc_hd__a21bo_1 c606 (.A1(net592),
    .A2(net591),
    .B1_N(net594),
    .X(net598));
 sky130_fd_sc_hd__buf_1 c607 (.A(net892),
    .X(net599));
 sky130_fd_sc_hd__xnor2_1 c608 (.A(net586),
    .B(net599),
    .Y(net600));
 sky130_fd_sc_hd__xnor2_1 c609 (.A(net600),
    .B(net597),
    .Y(net601));
 sky130_fd_sc_hd__a31o_1 c61 (.A1(net36),
    .A2(clknet_1_1__leaf_net27),
    .A3(clknet_1_0__leaf_net34),
    .B1(clknet_1_0__leaf_net912),
    .X(net38));
 sky130_fd_sc_hd__sdfxtp_1 c610 (.CLK(clknet_4_13_0_clk),
    .D(net590),
    .SCD(net594),
    .SCE(net587),
    .Q(net602));
 sky130_fd_sc_hd__a21bo_1 c611 (.A1(net597),
    .A2(net591),
    .B1_N(net602),
    .X(net603));
 sky130_fd_sc_hd__mux4_1 c612 (.A0(net603),
    .A1(net588),
    .A2(net594),
    .A3(net602),
    .S0(net592),
    .S1(net1067),
    .X(net604));
 sky130_fd_sc_hd__a21bo_1 c613 (.A1(net596),
    .A2(net602),
    .B1_N(net992),
    .X(net605));
 sky130_fd_sc_hd__a31o_1 c614 (.A1(net602),
    .A2(net605),
    .A3(net594),
    .B1(net1045),
    .X(net606));
 sky130_fd_sc_hd__a31o_1 c615 (.A1(net599),
    .A2(net606),
    .A3(net602),
    .B1(net1045),
    .X(net607));
 sky130_fd_sc_hd__dlymetal6s2s_1 c616 (.A(net978),
    .X(net608));
 sky130_fd_sc_hd__buf_1 c617 (.A(net608),
    .X(net609));
 sky130_fd_sc_hd__buf_1 c618 (.A(net609),
    .X(net610));
 sky130_fd_sc_hd__clkbuf_1 c619 (.A(net905),
    .X(net611));
 sky130_fd_sc_hd__a41o_1 c62 (.A1(clknet_1_1__leaf_net34),
    .A2(net31),
    .A3(clknet_1_0__leaf_net22),
    .A4(clknet_1_1__leaf_net20),
    .B1(net979),
    .X(net39));
 sky130_fd_sc_hd__buf_1 c620 (.A(net911),
    .X(net612));
 sky130_fd_sc_hd__buf_1 c621 (.A(net911),
    .X(net613));
 sky130_fd_sc_hd__clkbuf_4 c622 (.A(net905),
    .X(net614));
 sky130_fd_sc_hd__a21bo_1 c623 (.A1(net612),
    .A2(net613),
    .B1_N(net614),
    .X(net615));
 sky130_fd_sc_hd__xnor2_2 c624 (.A(net614),
    .B(net977),
    .Y(net616));
 sky130_fd_sc_hd__xnor2_2 c625 (.A(net615),
    .B(net608),
    .Y(net617));
 sky130_fd_sc_hd__xnor2_1 c626 (.A(net609),
    .B(net612),
    .Y(net618));
 sky130_fd_sc_hd__xnor2_1 c627 (.A(net616),
    .B(net614),
    .Y(net619));
 sky130_fd_sc_hd__xnor2_1 c628 (.A(net613),
    .B(net977),
    .Y(net1019));
 sky130_fd_sc_hd__buf_1 c629 (.A(net911),
    .X(net620));
 sky130_fd_sc_hd__a41o_1 c63 (.A1(net36),
    .A2(clknet_1_0__leaf_net34),
    .A3(clknet_1_1__leaf_net23),
    .A4(clknet_1_1__leaf_net912),
    .B1(net927),
    .X(net40));
 sky130_fd_sc_hd__xnor2_2 c630 (.A(net617),
    .B(net616),
    .Y(net621));
 sky130_fd_sc_hd__xnor2_1 c631 (.A(net615),
    .B(net620),
    .Y(net622));
 sky130_fd_sc_hd__xnor2_1 c632 (.A(net619),
    .B(net620),
    .Y(net623));
 sky130_fd_sc_hd__clkbuf_1 c633 (.A(net919),
    .X(net624));
 sky130_fd_sc_hd__a31o_1 c634 (.A1(net611),
    .A2(net623),
    .A3(net617),
    .B1(net621),
    .X(net625));
 sky130_fd_sc_hd__clkbuf_1 c635 (.A(net941),
    .X(net626));
 sky130_fd_sc_hd__a21bo_1 c636 (.A1(net622),
    .A2(net626),
    .B1_N(net868),
    .X(net627));
 sky130_fd_sc_hd__mux4_1 c637 (.A0(net627),
    .A1(net626),
    .A2(net611),
    .A3(net621),
    .S0(net610),
    .X(net868));
 sky130_fd_sc_hd__a31o_1 c64 (.A1(clknet_1_1__leaf_net26),
    .A2(net30),
    .A3(clknet_1_1__leaf_net34),
    .B1(net927),
    .X(net41));
 sky130_fd_sc_hd__buf_1 c65 (.A(clknet_1_1__leaf_net951),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_2 c651 (.A(net1021),
    .X(net1025));
 sky130_fd_sc_hd__clkbuf_2 c652 (.A(net1054),
    .X(net1022));
 sky130_fd_sc_hd__a21bo_1 c653 (.A1(net1022),
    .A2(net517),
    .B1_N(net867),
    .X(net1024));
 sky130_fd_sc_hd__a31o_1 c654 (.A1(net1024),
    .A2(net1025),
    .A3(net510),
    .B1(net1022),
    .X(net1027));
 sky130_fd_sc_hd__a21bo_1 c655 (.A1(net510),
    .A2(net1025),
    .B1_N(net1024),
    .X(net1030));
 sky130_fd_sc_hd__sdfrtp_1 c656 (.CLK(clknet_4_14_0_clk),
    .D(net1030),
    .RESET_B(net1022),
    .SCD(net1024),
    .SCE(net1025),
    .Q(net1023));
 sky130_fd_sc_hd__mux4_1 c657 (.A0(net1023),
    .A1(net1025),
    .A2(net1030),
    .A3(net1024),
    .S0(net1022),
    .S1(net510),
    .X(net629));
 sky130_fd_sc_hd__mux4_1 c658 (.A0(net621),
    .A1(net1022),
    .A2(net1023),
    .A3(net1024),
    .S0(net1025),
    .S1(clknet_1_0__leaf_net1020),
    .X(net630));
 sky130_fd_sc_hd__mux4_1 c659 (.A0(net1025),
    .A1(net1023),
    .A2(net1022),
    .A3(net1024),
    .S0(net1021),
    .S1(clknet_1_0__leaf_net1020),
    .X(net1018));
 sky130_fd_sc_hd__buf_2 c66 (.A(net948),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_2 c660 (.A(net541),
    .X(net631));
 sky130_fd_sc_hd__clkbuf_1 c661 (.A(net631),
    .X(net632));
 sky130_fd_sc_hd__clkbuf_2 c662 (.A(net631),
    .X(net633));
 sky130_fd_sc_hd__xnor2_2 c663 (.A(net633),
    .B(net631),
    .Y(net634));
 sky130_fd_sc_hd__clkbuf_1 c664 (.X(net635));
 sky130_fd_sc_hd__xnor2_1 c665 (.A(net633),
    .B(net631),
    .Y(net636));
 sky130_fd_sc_hd__clkbuf_1 c666 (.A(net769),
    .X(net637));
 sky130_fd_sc_hd__buf_1 c667 (.A(net1072),
    .X(net638));
 sky130_fd_sc_hd__clkbuf_8 c668 (.A(net803),
    .X(net639));
 sky130_fd_sc_hd__xnor2_2 c669 (.A(net638),
    .B(net639),
    .Y(net640));
 sky130_fd_sc_hd__clkbuf_2 c67 (.A(net43),
    .X(net44));
 sky130_fd_sc_hd__buf_1 c670 (.A(net1053),
    .X(net641));
 sky130_fd_sc_hd__xnor2_1 c671 (.A(net635),
    .B(net633),
    .Y(net642));
 sky130_fd_sc_hd__buf_1 c672 (.A(net819),
    .X(net643));
 sky130_fd_sc_hd__xnor2_1 c673 (.A(net643),
    .B(net641),
    .Y(net644));
 sky130_fd_sc_hd__xnor2_1 c674 (.A(net401),
    .B(net640),
    .Y(net645));
 sky130_fd_sc_hd__xnor2_1 c675 (.A(net640),
    .B(net643),
    .Y(net646));
 sky130_fd_sc_hd__a31o_1 c676 (.A1(net645),
    .A2(net646),
    .A3(net640),
    .B1(net1070),
    .X(net647));
 sky130_fd_sc_hd__xnor2_1 c677 (.A(net641),
    .B(net644),
    .Y(net648));
 sky130_fd_sc_hd__xnor2_1 c678 (.A(net644),
    .B(net646),
    .Y(net649));
 sky130_fd_sc_hd__clkbuf_1 c679 (.A(net824),
    .X(net650));
 sky130_fd_sc_hd__xnor2_2 c68 (.A(net1035),
    .B(net44),
    .Y(net45));
 sky130_fd_sc_hd__a31o_1 c680 (.A1(net648),
    .A2(net640),
    .A3(net645),
    .B1(net634),
    .X(net651));
 sky130_fd_sc_hd__xnor2_1 c681 (.A(net650),
    .B(net872),
    .Y(net652));
 sky130_fd_sc_hd__clkbuf_4 c682 (.X(net653));
 sky130_fd_sc_hd__clkbuf_4 c683 (.A(net758),
    .X(net654));
 sky130_fd_sc_hd__xnor2_4 c684 (.A(net639),
    .B(net654),
    .Y(net655));
 sky130_fd_sc_hd__xnor2_1 c685 (.A(net654),
    .B(net653),
    .Y(net656));
 sky130_fd_sc_hd__xnor2_1 c686 (.A(net654),
    .B(net653),
    .Y(net657));
 sky130_fd_sc_hd__xnor2_4 c687 (.A(net653),
    .B(net639),
    .Y(net658));
 sky130_fd_sc_hd__xnor2_4 c688 (.A(net655),
    .B(net639),
    .Y(net659));
 sky130_fd_sc_hd__buf_1 c689 (.A(net788),
    .X(net660));
 sky130_fd_sc_hd__clkbuf_1 c69 (.A(net44),
    .X(net46));
 sky130_fd_sc_hd__xnor2_4 c690 (.A(net658),
    .B(net659),
    .Y(net661));
 sky130_fd_sc_hd__xnor2_1 c691 (.A(net657),
    .B(net653),
    .Y(net662));
 sky130_fd_sc_hd__xnor2_1 c692 (.A(net653),
    .B(net662),
    .Y(net663));
 sky130_fd_sc_hd__clkbuf_1 c693 (.A(net964),
    .X(net664));
 sky130_fd_sc_hd__dfbbn_1 c694 (.CLK_N(clknet_4_8_0_clk),
    .D(net656),
    .RESET_B(net660),
    .SET_B(net661),
    .Q(net666),
    .Q_N(net665));
 sky130_fd_sc_hd__xnor2_1 c695 (.A(net659),
    .B(net654),
    .Y(net667));
 sky130_fd_sc_hd__clkbuf_1 c696 (.A(net802),
    .X(net668));
 sky130_fd_sc_hd__a21bo_1 c697 (.A1(net660),
    .A2(net668),
    .B1_N(net665),
    .X(net669));
 sky130_fd_sc_hd__a21bo_1 c698 (.A1(net658),
    .A2(net656),
    .B1_N(net669),
    .X(net670));
 sky130_fd_sc_hd__a21bo_1 c699 (.A1(net670),
    .A2(net669),
    .B1_N(net652),
    .X(net671));
 sky130_fd_sc_hd__xnor2_1 c70 (.A(net44),
    .B(net43),
    .Y(net47));
 sky130_fd_sc_hd__a21bo_1 c700 (.A1(net666),
    .A2(net668),
    .B1_N(net671),
    .X(net672));
 sky130_fd_sc_hd__dfbbn_1 c701 (.CLK_N(clknet_4_8_0_clk),
    .D(net671),
    .RESET_B(net670),
    .SET_B(net659),
    .Q(net674),
    .Q_N(net673));
 sky130_fd_sc_hd__a31o_1 c702 (.A1(net667),
    .A2(net674),
    .A3(net660),
    .B1(net654),
    .X(net675));
 sky130_fd_sc_hd__a31o_1 c703 (.A1(net655),
    .A2(net673),
    .A3(net659),
    .B1(net924),
    .X(net676));
 sky130_fd_sc_hd__clkbuf_2 c704 (.A(net762),
    .X(net677));
 sky130_fd_sc_hd__clkbuf_1 c705 (.A(net677),
    .X(net678));
 sky130_fd_sc_hd__clkbuf_1 c706 (.A(net762),
    .X(net679));
 sky130_fd_sc_hd__clkbuf_1 c707 (.A(net971),
    .X(net680));
 sky130_fd_sc_hd__clkbuf_1 c708 (.A(net971),
    .X(net681));
 sky130_fd_sc_hd__buf_1 c709 (.A(net680),
    .X(net682));
 sky130_fd_sc_hd__buf_1 c71 (.A(net777),
    .X(net48));
 sky130_fd_sc_hd__buf_4 c710 (.A(net1034),
    .X(net683));
 sky130_fd_sc_hd__xnor2_4 c711 (.A(net677),
    .B(net683),
    .Y(net684));
 sky130_fd_sc_hd__a21bo_1 c712 (.A1(net681),
    .A2(net683),
    .B1_N(net684),
    .X(net685));
 sky130_fd_sc_hd__buf_1 c713 (.A(net803),
    .X(net686));
 sky130_fd_sc_hd__xnor2_1 c714 (.A(net678),
    .B(net684),
    .Y(net687));
 sky130_fd_sc_hd__xnor2_1 c715 (.A(net662),
    .B(net683),
    .Y(net688));
 sky130_fd_sc_hd__xnor2_2 c716 (.A(net682),
    .B(net684),
    .Y(net689));
 sky130_fd_sc_hd__xnor2_1 c717 (.A(net687),
    .B(net686),
    .Y(net690));
 sky130_fd_sc_hd__clkbuf_1 c718 (.A(net978),
    .X(net691));
 sky130_fd_sc_hd__clkbuf_1 c719 (.A(net957),
    .X(net692));
 sky130_fd_sc_hd__dlymetal6s2s_1 c72 (.A(net901),
    .X(net49));
 sky130_fd_sc_hd__mux4_1 c720 (.A0(net692),
    .A1(net685),
    .A2(net688),
    .A3(net689),
    .S0(net684),
    .S1(net686),
    .X(net693));
 sky130_fd_sc_hd__a31o_1 c721 (.A1(net691),
    .A2(net684),
    .A3(net689),
    .B1(clknet_1_1__leaf_net993),
    .X(net694));
 sky130_fd_sc_hd__mux4_1 c722 (.A0(net679),
    .A1(clknet_1_0__leaf_net694),
    .A2(net661),
    .A3(net689),
    .S0(net683),
    .S1(clknet_1_0__leaf_net993),
    .X(net695));
 sky130_fd_sc_hd__a31o_1 c723 (.A1(clknet_1_1__leaf_net694),
    .A2(net689),
    .A3(net684),
    .B1(net968),
    .X(net696));
 sky130_fd_sc_hd__a31o_1 c724 (.A1(net686),
    .A2(clknet_1_0__leaf_net694),
    .A3(net689),
    .B1(net968),
    .X(net697));
 sky130_fd_sc_hd__a31o_1 c725 (.A1(net689),
    .A2(clknet_1_1__leaf_net694),
    .A3(net669),
    .B1(clknet_1_1__leaf_net914),
    .X(net698));
 sky130_fd_sc_hd__clkbuf_1 c726 (.A(net767),
    .X(net699));
 sky130_fd_sc_hd__buf_2 c727 (.A(net767),
    .X(net700));
 sky130_fd_sc_hd__clkbuf_4 c728 (.A(net699),
    .X(net701));
 sky130_fd_sc_hd__xnor2_4 c729 (.A(net700),
    .B(net701),
    .Y(net702));
 sky130_fd_sc_hd__clkbuf_1 c73 (.A(net777),
    .X(net50));
 sky130_fd_sc_hd__buf_1 c730 (.A(net701),
    .X(net703));
 sky130_fd_sc_hd__xnor2_1 c731 (.A(net702),
    .B(net701),
    .Y(net704));
 sky130_fd_sc_hd__xnor2_1 c732 (.A(net683),
    .B(net702),
    .Y(net705));
 sky130_fd_sc_hd__xnor2_2 c733 (.A(net701),
    .B(net700),
    .Y(net706));
 sky130_fd_sc_hd__clkbuf_1 c734 (.A(net961),
    .X(net707));
 sky130_fd_sc_hd__buf_1 c735 (.A(net964),
    .X(net708));
 sky130_fd_sc_hd__a21bo_1 c736 (.A1(net702),
    .A2(net708),
    .B1_N(net703),
    .X(net709));
 sky130_fd_sc_hd__buf_1 c737 (.A(clknet_1_1__leaf_net949),
    .X(net710));
 sky130_fd_sc_hd__xnor2_1 c738 (.A(net703),
    .B(net702),
    .Y(net711));
 sky130_fd_sc_hd__xnor2_1 c739 (.A(net706),
    .B(clknet_1_1__leaf_net710),
    .Y(net712));
 sky130_fd_sc_hd__xnor2_1 c74 (.A(net48),
    .B(net49),
    .Y(net51));
 sky130_fd_sc_hd__a21bo_1 c740 (.A1(net708),
    .A2(net711),
    .B1_N(net705),
    .X(net713));
 sky130_fd_sc_hd__a21bo_1 c741 (.A1(net585),
    .A2(net705),
    .B1_N(net706),
    .X(net714));
 sky130_fd_sc_hd__sdfbbn_1 c742 (.CLK_N(clknet_4_10_0_clk),
    .D(clknet_1_0__leaf_net710),
    .RESET_B(net683),
    .SCD(clknet_1_1__leaf_net712),
    .SCE(net953),
    .SET_B(net1041),
    .Q(net716),
    .Q_N(net715));
 sky130_fd_sc_hd__a21bo_1 c743 (.A1(clknet_1_0__leaf_net710),
    .A2(net716),
    .B1_N(net969),
    .X(net717));
 sky130_fd_sc_hd__buf_1 c744 (.A(net964),
    .X(net718));
 sky130_fd_sc_hd__a31o_1 c745 (.A1(net707),
    .A2(net716),
    .A3(clknet_1_1__leaf_net717),
    .B1(net702),
    .X(net719));
 sky130_fd_sc_hd__clkbuf_4 c746 (.A(net983),
    .X(net720));
 sky130_fd_sc_hd__mux4_1 c747 (.A0(clknet_1_1__leaf_net719),
    .A1(clknet_1_1__leaf_net717),
    .A2(net720),
    .A3(net683),
    .S0(net718),
    .S1(clknet_1_1__leaf_net914),
    .X(net721));
 sky130_fd_sc_hd__xnor2_2 c748 (.A(net614),
    .B(net867),
    .Y(net722));
 sky130_fd_sc_hd__xnor2_1 c749 (.A(net1031),
    .B(net614),
    .Y(net723));
 sky130_fd_sc_hd__clkbuf_1 c75 (.A(net855),
    .X(net52));
 sky130_fd_sc_hd__xnor2_1 c750 (.A(net718),
    .B(net1031),
    .Y(net724));
 sky130_fd_sc_hd__xnor2_2 c751 (.A(net720),
    .B(net953),
    .Y(net725));
 sky130_fd_sc_hd__xnor2_1 c752 (.A(net725),
    .B(net722),
    .Y(net1028));
 sky130_fd_sc_hd__xnor2_1 c753 (.A(net724),
    .B(net1031),
    .Y(net726));
 sky130_fd_sc_hd__xnor2_4 c754 (.A(net720),
    .B(net1031),
    .Y(net727));
 sky130_fd_sc_hd__xnor2_1 c755 (.A(net722),
    .B(net727),
    .Y(net728));
 sky130_fd_sc_hd__dfbbp_1 c756 (.CLK(clknet_4_11_0_clk),
    .D(net614),
    .RESET_B(net728),
    .SET_B(net727),
    .Q(net730),
    .Q_N(net729));
 sky130_fd_sc_hd__a31o_1 c757 (.A1(net723),
    .A2(net727),
    .A3(net729),
    .B1(clknet_1_1__leaf_net949),
    .X(net731));
 sky130_fd_sc_hd__buf_1 c758 (.A(net920),
    .X(net732));
 sky130_fd_sc_hd__xnor2_2 c759 (.A(net730),
    .B(net732),
    .Y(net1017));
 sky130_fd_sc_hd__xnor2_1 c76 (.A(net50),
    .B(net49),
    .Y(net53));
 sky130_fd_sc_hd__buf_1 c760 (.A(net920),
    .X(net733));
 sky130_fd_sc_hd__xnor2_1 c761 (.A(net725),
    .B(net733),
    .Y(net734));
 sky130_fd_sc_hd__a41o_1 c762 (.A1(net726),
    .A2(net728),
    .A3(net723),
    .A4(net1017),
    .B1(net1031),
    .X(net735));
 sky130_fd_sc_hd__a21bo_1 c763 (.A1(net733),
    .A2(net730),
    .B1_N(net727),
    .X(net736));
 sky130_fd_sc_hd__a21bo_2 c764 (.A1(net734),
    .A2(net1031),
    .B1_N(net727),
    .X(net737));
 sky130_fd_sc_hd__clkbuf_1 c765 (.A(net911),
    .X(net738));
 sky130_fd_sc_hd__clkbuf_1 c766 (.A(net961),
    .X(net739));
 sky130_fd_sc_hd__sdfbbn_1 c767 (.CLK_N(clknet_4_11_0_clk),
    .D(net732),
    .RESET_B(net736),
    .SCD(net727),
    .SCE(net737),
    .SET_B(net722),
    .Q(net1016),
    .Q_N(net740));
 sky130_fd_sc_hd__mux4_1 c768 (.A0(net728),
    .A1(net739),
    .A2(net1017),
    .A3(net740),
    .S0(net737),
    .S1(net727),
    .X(net741));
 sky130_fd_sc_hd__a21bo_1 c769 (.A1(net727),
    .A2(net725),
    .B1_N(net905),
    .X(net1029));
 sky130_fd_sc_hd__buf_1 c77 (.A(net976),
    .X(net54));
 sky130_fd_sc_hd__buf_1 c78 (.A(net900),
    .X(net55));
 sky130_fd_sc_hd__a21bo_1 c79 (.A1(net51),
    .A2(net53),
    .B1_N(net55),
    .X(net56));
 sky130_fd_sc_hd__a21bo_2 c80 (.A1(net56),
    .A2(net44),
    .B1_N(net53),
    .X(net57));
 sky130_fd_sc_hd__a21bo_1 c81 (.A1(net37),
    .A2(net56),
    .B1_N(net54),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_1 c82 (.A(net941),
    .X(net59));
 sky130_fd_sc_hd__a21bo_1 c83 (.A1(net52),
    .A2(net54),
    .B1_N(net55),
    .X(net60));
 sky130_fd_sc_hd__a21bo_1 c84 (.A1(net59),
    .A2(net55),
    .B1_N(net60),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_1 c85 (.A(net941),
    .X(net62));
 sky130_fd_sc_hd__a31o_1 c86 (.A1(net53),
    .A2(net60),
    .A3(net55),
    .B1(net57),
    .X(net63));
 sky130_fd_sc_hd__a41o_1 c87 (.A1(net62),
    .A2(net60),
    .A3(net57),
    .A4(net55),
    .X(net64));
 sky130_fd_sc_hd__buf_1 c88 (.A(net43),
    .X(net65));
 sky130_fd_sc_hd__buf_1 c89 (.A(net65),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_2 c90 (.A(net65),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_2 c91 (.A(net931),
    .X(net68));
 sky130_fd_sc_hd__buf_1 c92 (.A(net931),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_1 c93 (.A(net982),
    .X(net70));
 sky130_fd_sc_hd__xnor2_2 c94 (.A(net69),
    .B(net68),
    .Y(net71));
 sky130_fd_sc_hd__xnor2_1 c95 (.A(net71),
    .B(net68),
    .Y(net72));
 sky130_fd_sc_hd__clkbuf_2 c96 (.A(net808),
    .X(net73));
 sky130_fd_sc_hd__clkbuf_1 c97 (.A(net982),
    .X(net74));
 sky130_fd_sc_hd__dlymetal6s2s_1 c98 (.A(net928),
    .X(net75));
 sky130_fd_sc_hd__xnor2_2 c99 (.A(net75),
    .B(net71),
    .Y(net76));
 sky130_fd_sc_hd__mux4_1 merge782 (.A0(net7),
    .A1(net995),
    .A2(net3),
    .A3(net11),
    .S0(net12),
    .S1(net13),
    .X(net742));
 sky130_fd_sc_hd__a21bo_1 merge783 (.A1(clknet_1_1__leaf_net226),
    .A2(clknet_1_0__leaf_net325),
    .B1_N(net339),
    .X(net743));
 sky130_fd_sc_hd__a31o_1 merge784 (.A1(net252),
    .A2(net251),
    .A3(net256),
    .B1(net253),
    .X(net744));
 sky130_fd_sc_hd__a31o_1 merge785 (.A1(net118),
    .A2(net117),
    .A3(net122),
    .B1(net997),
    .X(net745));
 sky130_fd_sc_hd__a31o_1 merge786 (.A1(clknet_1_1__leaf_net89),
    .A2(net94),
    .A3(net93),
    .B1(clknet_1_0__leaf_net95),
    .X(net746));
 sky130_fd_sc_hd__buf_1 merge787 (.A(clknet_1_1__leaf_net950),
    .X(net747));
 sky130_fd_sc_hd__a21bo_1 merge788 (.A1(net430),
    .A2(net431),
    .B1_N(net432),
    .X(net748));
 sky130_fd_sc_hd__a31o_1 merge789 (.A1(net731),
    .A2(net729),
    .A3(net1017),
    .B1(net726),
    .X(net749));
 sky130_fd_sc_hd__a21bo_1 merge790 (.A1(net609),
    .A2(net610),
    .B1_N(net608),
    .X(net750));
 sky130_fd_sc_hd__clkbuf_1 merge791 (.A(net940),
    .X(net751));
 sky130_fd_sc_hd__sdfxbp_1 merge792 (.CLK(clknet_4_10_0_clk),
    .D(net405),
    .SCD(net522),
    .SCE(net519),
    .Q(net753),
    .Q_N(net752));
 sky130_fd_sc_hd__a21bo_1 merge793 (.A1(net139),
    .A2(net140),
    .B1_N(net142),
    .X(net754));
 sky130_fd_sc_hd__a31o_1 merge794 (.A1(clknet_1_1__leaf_net160),
    .A2(clknet_1_1__leaf_net161),
    .A3(clknet_1_0__leaf_net162),
    .B1(net13),
    .X(net755));
 sky130_fd_sc_hd__clkbuf_1 merge795 (.A(net781),
    .X(net756));
 sky130_fd_sc_hd__a31o_1 merge796 (.A1(clknet_1_1__leaf_net162),
    .A2(net181),
    .A3(net297),
    .B1(net956),
    .X(net757));
 sky130_fd_sc_hd__sdfxbp_2 merge797 (.CLK(clknet_4_8_0_clk),
    .D(net652),
    .SCD(clknet_1_0__leaf_net563),
    .Q(net653),
    .Q_N(net758));
 sky130_fd_sc_hd__clkbuf_1 merge798 (.A(net955),
    .X(net760));
 sky130_fd_sc_hd__buf_1 merge799 (.A(net929),
    .X(net761));
 sky130_fd_sc_hd__clkbuf_1 merge800 (.A(net940),
    .X(net762));
 sky130_fd_sc_hd__a21bo_1 merge801 (.A1(net544),
    .A2(net543),
    .B1_N(net991),
    .X(net763));
 sky130_fd_sc_hd__buf_1 merge802 (.A(clknet_1_0__leaf_net950),
    .X(net764));
 sky130_fd_sc_hd__a21bo_1 merge803 (.A1(net182),
    .A2(net184),
    .B1_N(net57),
    .X(net765));
 sky130_fd_sc_hd__a31o_1 merge804 (.A1(net65),
    .A2(net67),
    .A3(net66),
    .B1(net68),
    .X(net766));
 sky130_fd_sc_hd__clkbuf_1 merge805 (.A(net958),
    .X(net767));
 sky130_fd_sc_hd__a31o_1 merge806 (.A1(clknet_1_0__leaf_net226),
    .A2(net230),
    .A3(net231),
    .B1(net959),
    .X(net768));
 sky130_fd_sc_hd__sdfxtp_1 merge807 (.CLK(clknet_4_8_0_clk),
    .D(net634),
    .SCD(net525),
    .Q(net635));
 sky130_fd_sc_hd__a21bo_1 merge808 (.A1(net19),
    .A2(net1006),
    .B1_N(net13),
    .X(net770));
 sky130_fd_sc_hd__clkbuf_1 merge809 (.A(net980),
    .X(net771));
 sky130_fd_sc_hd__a31o_1 merge810 (.A1(net590),
    .A2(net460),
    .A3(net593),
    .B1(net575),
    .X(net772));
 sky130_fd_sc_hd__buf_1 merge811 (.A(net932),
    .X(net773));
 sky130_fd_sc_hd__a21bo_1 merge812 (.A1(clknet_1_0__leaf_net272),
    .A2(net264),
    .B1_N(net273),
    .X(net774));
 sky130_fd_sc_hd__clkbuf_1 merge813 (.A(net940),
    .X(net775));
 sky130_fd_sc_hd__mux4_1 merge814 (.A0(net589),
    .A1(net1019),
    .A2(net381),
    .A3(net517),
    .S0(net621),
    .S1(net1025),
    .X(net776));
 sky130_fd_sc_hd__clkbuf_1 merge815 (.A(net944),
    .X(net777));
 sky130_fd_sc_hd__sdfrtp_1 merge816 (.CLK(clknet_4_4_0_clk),
    .D(net359),
    .RESET_B(net358),
    .SCD(clknet_1_1__leaf_net213),
    .SCE(clknet_1_1__leaf_net207),
    .Q(net778));
 sky130_fd_sc_hd__a31o_1 merge817 (.A1(net601),
    .A2(net433),
    .A3(net439),
    .B1(clknet_1_0__leaf_net949),
    .X(net779));
 sky130_fd_sc_hd__a31o_1 merge818 (.A1(net119),
    .A2(net123),
    .A3(net140),
    .B1(net142),
    .X(net780));
 sky130_fd_sc_hd__clkbuf_1 merge819 (.A(net871),
    .X(net781));
 sky130_fd_sc_hd__a31o_1 merge820 (.A1(net176),
    .A2(clknet_1_1__leaf_net168),
    .A3(net169),
    .B1(net165),
    .X(net782));
 sky130_fd_sc_hd__a31o_1 merge821 (.A1(net389),
    .A2(net386),
    .A3(net434),
    .B1(net432),
    .X(net783));
 sky130_fd_sc_hd__a31o_1 merge822 (.A1(net300),
    .A2(net302),
    .A3(net138),
    .B1(net142),
    .X(net784));
 sky130_fd_sc_hd__a31o_1 merge823 (.A1(clknet_1_0__leaf_net317),
    .A2(clknet_1_1__leaf_net325),
    .A3(net45),
    .B1(net47),
    .X(net785));
 sky130_fd_sc_hd__a31o_1 merge824 (.A1(net296),
    .A2(net302),
    .A3(net336),
    .B1(net327),
    .X(net786));
 sky130_fd_sc_hd__sdfsbp_1 merge825 (.CLK(clknet_4_10_0_clk),
    .D(net659),
    .SCD(clknet_1_0__leaf_net563),
    .SCE(net522),
    .SET_B(net526),
    .Q(net788),
    .Q_N(net787));
 sky130_fd_sc_hd__a31o_1 merge826 (.A1(net190),
    .A2(net193),
    .A3(net165),
    .B1(clknet_1_0__leaf_net168),
    .X(net789));
 sky130_fd_sc_hd__a31o_1 merge827 (.A1(net349),
    .A2(net484),
    .A3(net346),
    .B1(net345),
    .X(net790));
 sky130_fd_sc_hd__a31o_1 merge828 (.A1(net453),
    .A2(net456),
    .A3(net435),
    .B1(net434),
    .X(net791));
 sky130_fd_sc_hd__sdfsbp_1 merge829 (.CLK(clknet_4_14_0_clk),
    .D(net524),
    .SCD(net523),
    .SCE(net261),
    .SET_B(net252),
    .Q(net793),
    .Q_N(net792));
 sky130_fd_sc_hd__a31o_1 merge830 (.A1(net690),
    .A2(net683),
    .A3(net565),
    .B1(net572),
    .X(net794));
 sky130_fd_sc_hd__a31o_1 merge831 (.A1(net189),
    .A2(net184),
    .A3(net461),
    .B1(net455),
    .X(net795));
 sky130_fd_sc_hd__a31o_1 merge832 (.A1(net301),
    .A2(net300),
    .A3(net451),
    .B1(net453),
    .X(net796));
 sky130_fd_sc_hd__a31o_1 merge833 (.A1(net322),
    .A2(clknet_1_0__leaf_net321),
    .A3(clknet_1_1__leaf_net29),
    .B1(clknet_1_1__leaf_net24),
    .X(net797));
 sky130_fd_sc_hd__a31o_1 merge834 (.A1(net260),
    .A2(net259),
    .A3(net281),
    .B1(net284),
    .X(net798));
 sky130_fd_sc_hd__a31o_1 merge835 (.A1(clknet_1_1__leaf_net272),
    .A2(net276),
    .A3(net577),
    .B1(net576),
    .X(net799));
 sky130_fd_sc_hd__a31o_1 merge836 (.A1(net566),
    .A2(clknet_1_1__leaf_net563),
    .A3(net610),
    .B1(net1019),
    .X(net800));
 sky130_fd_sc_hd__a31o_1 merge837 (.A1(net705),
    .A2(net701),
    .A3(net737),
    .B1(net738),
    .X(net801));
 sky130_fd_sc_hd__sdfstp_1 merge838 (.CLK(clknet_4_8_0_clk),
    .D(net664),
    .SCD(net661),
    .SCE(net632),
    .SET_B(net634),
    .Q(net802));
 sky130_fd_sc_hd__sdfstp_1 merge839 (.CLK(clknet_4_8_0_clk),
    .D(net636),
    .SCD(net634),
    .SCE(net661),
    .SET_B(net684),
    .Q(net803));
 sky130_fd_sc_hd__a31o_1 merge840 (.A1(net306),
    .A2(net302),
    .A3(net274),
    .B1(clknet_1_0__leaf_net272),
    .X(net804));
 sky130_fd_sc_hd__a31o_1 merge841 (.A1(net362),
    .A2(net365),
    .A3(clknet_1_0__leaf_net321),
    .B1(clknet_1_0__leaf_net324),
    .X(net805));
 sky130_fd_sc_hd__a31o_1 merge842 (.A1(net483),
    .A2(clknet_1_0__leaf_net482),
    .A3(net476),
    .B1(net478),
    .X(net806));
 sky130_fd_sc_hd__sdfstp_1 merge843 (.CLK(clknet_4_8_0_clk),
    .D(net637),
    .SCD(net634),
    .SCE(net421),
    .SET_B(net422),
    .Q(net807));
 sky130_fd_sc_hd__sedfxbp_1 merge844 (.CLK(clknet_4_1_0_clk),
    .D(net211),
    .DE(net66),
    .SCD(net71),
    .SCE(net1069),
    .Q(net809),
    .Q_N(net808));
 sky130_fd_sc_hd__a31o_1 merge845 (.A1(net572),
    .A2(net569),
    .A3(net704),
    .B1(net706),
    .X(net810));
 sky130_fd_sc_hd__a31o_1 merge846 (.A1(net65),
    .A2(net57),
    .A3(net68),
    .B1(net67),
    .X(net811));
 sky130_fd_sc_hd__a31o_1 merge847 (.A1(clknet_1_1__leaf_net197),
    .A2(clknet_1_0__leaf_net201),
    .A3(clknet_1_1__leaf_net162),
    .B1(net187),
    .X(net812));
 sky130_fd_sc_hd__a31o_1 merge848 (.A1(net165),
    .A2(clknet_1_0__leaf_net160),
    .A3(net45),
    .B1(net48),
    .X(net813));
 sky130_fd_sc_hd__a41o_1 merge849 (.A1(net608),
    .A2(net610),
    .A3(net609),
    .A4(net613),
    .B1(net943),
    .X(net814));
 sky130_fd_sc_hd__a31o_1 merge850 (.A1(net486),
    .A2(net478),
    .A3(net459),
    .B1(net965),
    .X(net815));
 sky130_fd_sc_hd__a31o_1 merge851 (.A1(net67),
    .A2(net68),
    .A3(clknet_1_1__leaf_net91),
    .B1(net231),
    .X(net816));
 sky130_fd_sc_hd__a31o_1 merge852 (.A1(net392),
    .A2(net386),
    .A3(clknet_1_0__leaf_net563),
    .B1(net924),
    .X(net817));
 sky130_fd_sc_hd__sedfxbp_1 merge853 (.CLK(clknet_4_8_0_clk),
    .D(net642),
    .DE(net639),
    .SCD(net424),
    .SCE(net434),
    .Q(net819),
    .Q_N(net818));
 sky130_fd_sc_hd__a31o_1 merge854 (.A1(net389),
    .A2(net392),
    .A3(clknet_1_1__leaf_net25),
    .B1(clknet_1_1__leaf_net912),
    .X(net820));
 sky130_fd_sc_hd__a31o_1 merge855 (.A1(net406),
    .A2(net414),
    .A3(clknet_1_0__leaf_net330),
    .B1(clknet_1_0__leaf_net329),
    .X(net821));
 sky130_fd_sc_hd__mux4_1 merge856 (.A0(net618),
    .A1(net613),
    .A2(net617),
    .A3(net728),
    .S0(net737),
    .S1(net905),
    .X(net822));
 sky130_fd_sc_hd__a31o_1 merge857 (.A1(clknet_1_1__leaf_net321),
    .A2(clknet_1_1__leaf_net317),
    .A3(net415),
    .B1(net420),
    .X(net823));
 sky130_fd_sc_hd__sedfxtp_1 merge858 (.CLK(clknet_4_8_0_clk),
    .D(net649),
    .DE(net419),
    .SCD(net414),
    .SCE(net872),
    .Q(net824));
 sky130_fd_sc_hd__a31o_1 merge859 (.A1(clknet_1_0__leaf_net21),
    .A2(clknet_1_0__leaf_net25),
    .A3(net408),
    .B1(net414),
    .X(net825));
 sky130_fd_sc_hd__a31o_1 merge860 (.A1(net219),
    .A2(net345),
    .A3(net13),
    .B1(clknet_1_1__leaf_net20),
    .X(net826));
 sky130_fd_sc_hd__sedfxtp_1 merge861 (.CLK(clknet_4_3_0_clk),
    .D(net369),
    .DE(net362),
    .SCD(net343),
    .SCE(net345),
    .Q(net827));
 sky130_fd_sc_hd__a41o_1 merge862 (.A1(net228),
    .A2(net365),
    .A3(net70),
    .A4(clknet_1_0__leaf_net81),
    .B1(net963),
    .X(net828));
 sky130_fd_sc_hd__a21bo_1 merge863 (.A1(net669),
    .A2(net575),
    .B1_N(net676),
    .X(net829));
 sky130_fd_sc_hd__a41o_1 merge864 (.A1(net394),
    .A2(net389),
    .A3(net392),
    .A4(net393),
    .B1(net397),
    .X(net830));
 sky130_fd_sc_hd__mux4_1 merge865 (.A0(net125),
    .A1(net123),
    .A2(net122),
    .A3(net140),
    .S0(net142),
    .S1(net870),
    .X(net831));
 sky130_fd_sc_hd__mux4_1 merge866 (.A0(clknet_1_1__leaf_net357),
    .A1(clknet_1_0__leaf_net353),
    .A2(net347),
    .A3(net188),
    .S0(net187),
    .S1(net183),
    .X(net832));
 sky130_fd_sc_hd__mux4_1 merge867 (.A0(net47),
    .A1(net43),
    .A2(net46),
    .A3(net49),
    .S0(net54),
    .S1(net979),
    .X(net833));
 sky130_fd_sc_hd__mux4_1 merge868 (.A0(clknet_1_1__leaf_net329),
    .A1(clknet_1_1__leaf_net324),
    .A2(net322),
    .A3(net488),
    .S0(net481),
    .S1(net478),
    .X(net834));
 sky130_fd_sc_hd__mux4_1 merge869 (.A0(clknet_1_1__leaf_net42),
    .A1(net47),
    .A2(net45),
    .A3(net509),
    .S0(net922),
    .S1(net958),
    .X(net835));
 sky130_fd_sc_hd__mux4_1 merge870 (.A0(net311),
    .A1(net305),
    .A2(net307),
    .A3(net249),
    .S0(net362),
    .S1(net365),
    .X(net836));
 sky130_fd_sc_hd__mux4_1 merge871 (.A0(net366),
    .A1(net365),
    .A2(clknet_1_0__leaf_net712),
    .A3(clknet_1_0__leaf_net717),
    .S0(clknet_1_0__leaf_net719),
    .S1(net945),
    .X(net837));
 sky130_fd_sc_hd__mux4_1 merge872 (.A0(net67),
    .A1(clknet_1_1__leaf_net210),
    .A2(clknet_1_0__leaf_net213),
    .A3(net130),
    .S0(net118),
    .S1(net124),
    .X(net838));
 sky130_fd_sc_hd__a41o_1 merge873 (.A1(net395),
    .A2(net399),
    .A3(net397),
    .A4(net398),
    .B1(net390),
    .X(net839));
 sky130_fd_sc_hd__mux4_1 merge874 (.A0(net151),
    .A1(net152),
    .A2(net142),
    .A3(net124),
    .S0(net131),
    .S1(net130),
    .X(net840));
 sky130_fd_sc_hd__mux4_1 merge875 (.A0(net554),
    .A1(net553),
    .A2(net252),
    .A3(net258),
    .S0(net254),
    .S1(net1064),
    .X(net841));
 sky130_fd_sc_hd__mux4_1 merge876 (.A0(net709),
    .A1(net708),
    .A2(net706),
    .A3(net439),
    .S0(net436),
    .S1(net970),
    .X(net842));
 sky130_fd_sc_hd__a41o_1 merge877 (.A1(net259),
    .A2(net257),
    .A3(net260),
    .A4(net263),
    .B1(net264),
    .X(net843));
 sky130_fd_sc_hd__mux4_1 merge878 (.A0(net663),
    .A1(net660),
    .A2(net661),
    .A3(clknet_1_0__leaf_net717),
    .S0(net715),
    .S1(net709),
    .X(net844));
 sky130_fd_sc_hd__mux4_1 merge879 (.A0(net428),
    .A1(clknet_1_1__leaf_net563),
    .A2(net564),
    .A3(net378),
    .S0(net248),
    .S1(net931),
    .X(net845));
 sky130_fd_sc_hd__mux4_1 merge880 (.A0(net688),
    .A1(net689),
    .A2(net683),
    .A3(net1012),
    .S0(clknet_1_0__leaf_net145),
    .S1(net140),
    .X(net846));
 sky130_fd_sc_hd__mux4_1 merge881 (.A0(net368),
    .A1(net366),
    .A2(net362),
    .A3(clknet_1_1__leaf_net81),
    .S0(net84),
    .S1(clknet_1_0__leaf_net85),
    .X(net847));
 sky130_fd_sc_hd__mux4_1 merge882 (.A0(net367),
    .A1(net509),
    .A2(net300),
    .A3(net303),
    .S0(net308),
    .S1(net965),
    .X(net848));
 sky130_fd_sc_hd__mux4_1 merge883 (.A0(net410),
    .A1(net1032),
    .A2(net409),
    .A3(net132),
    .S0(clknet_1_0__leaf_net127),
    .S1(net130),
    .X(net849));
 sky130_fd_sc_hd__mux4_1 merge884 (.A0(net307),
    .A1(net302),
    .A2(net477),
    .A3(net476),
    .S0(net478),
    .S1(net990),
    .X(net850));
 sky130_fd_sc_hd__mux4_1 merge885 (.A0(net624),
    .A1(net623),
    .A2(net620),
    .A3(net283),
    .S0(net278),
    .S1(net1058),
    .X(net851));
 sky130_fd_sc_hd__mux4_1 merge886 (.A0(net676),
    .A1(net575),
    .A2(net677),
    .A3(clknet_1_0__leaf_net498),
    .S0(clknet_1_0__leaf_net496),
    .S1(net481),
    .X(net852));
 sky130_fd_sc_hd__a41o_1 merge887 (.A1(net49),
    .A2(net57),
    .A3(net52),
    .A4(net61),
    .B1(net58),
    .X(net853));
 sky130_fd_sc_hd__xnor2_1 merge888 (.A(net696),
    .B(net697),
    .Y(net854));
 sky130_fd_sc_hd__dfrbp_1 merge889 (.CLK(clknet_4_6_0_clk),
    .D(net338),
    .RESET_B(net785),
    .Q(net856),
    .Q_N(net855));
 sky130_fd_sc_hd__xnor2_1 merge890 (.A(net714),
    .B(net721),
    .Y(net857));
 sky130_fd_sc_hd__xnor2_1 merge891 (.A(net38),
    .B(net40),
    .Y(net858));
 sky130_fd_sc_hd__xnor2_1 merge892 (.A(net462),
    .B(net464),
    .Y(net859));
 sky130_fd_sc_hd__xnor2_1 merge893 (.A(net154),
    .B(net157),
    .Y(net860));
 sky130_fd_sc_hd__xnor2_1 merge894 (.A(net78),
    .B(net83),
    .Y(net861));
 sky130_fd_sc_hd__xnor2_1 merge895 (.A(net672),
    .B(net675),
    .Y(net862));
 sky130_fd_sc_hd__xnor2_1 merge896 (.A(net173),
    .B(net174),
    .Y(net863));
 sky130_fd_sc_hd__xnor2_1 merge897 (.A(net288),
    .B(net289),
    .Y(net864));
 sky130_fd_sc_hd__xnor2_1 merge898 (.A(net417),
    .B(net426),
    .Y(net865));
 sky130_fd_sc_hd__xnor2_1 merge899 (.A(net348),
    .B(net351),
    .Y(net866));
 sky130_fd_sc_hd__dfrbp_1 merge900 (.CLK(clknet_4_14_0_clk),
    .D(net625),
    .Q(net868),
    .Q_N(net867));
 sky130_fd_sc_hd__xnor2_1 merge901 (.A(net111),
    .B(net115),
    .Y(net869));
 sky130_fd_sc_hd__dfrtn_1 merge902 (.CLK_N(clknet_4_13_0_clk),
    .D(net128),
    .RESET_B(net137),
    .Q(net870));
 sky130_fd_sc_hd__dfrtp_1 merge903 (.CLK(clknet_4_2_0_clk),
    .D(net403),
    .RESET_B(net783),
    .Q(net871));
 sky130_fd_sc_hd__dfrtp_1 merge904 (.CLK(clknet_4_8_0_clk),
    .D(net647),
    .RESET_B(net651),
    .Q(net872));
 sky130_fd_sc_hd__dfrtp_1 merge905 (.CLK(clknet_4_15_0_clk),
    .RESET_B(net1057),
    .Q(net873));
 sky130_fd_sc_hd__xnor2_1 merge906 (.A(net14),
    .B(net17),
    .Y(net874));
 sky130_fd_sc_hd__dfsbp_1 merge907 (.CLK(clknet_4_6_0_clk),
    .D(net310),
    .SET_B(net757),
    .Q(net876),
    .Q_N(net875));
 sky130_fd_sc_hd__xnor2_1 merge908 (.A(net196),
    .B(net198),
    .Y(net877));
 sky130_fd_sc_hd__dfsbp_1 merge909 (.CLK(clknet_4_4_0_clk),
    .D(net212),
    .SET_B(net223),
    .Q(net879),
    .Q_N(net878));
 sky130_fd_sc_hd__xnor2_1 merge910 (.A(net735),
    .B(net741),
    .Y(net880));
 sky130_fd_sc_hd__dfstp_1 merge911 (.CLK(clknet_4_14_0_clk),
    .D(net776),
    .SET_B(net630),
    .Q(net1021));
 sky130_fd_sc_hd__xnor2_1 merge912 (.A(net505),
    .B(net511),
    .Y(net881));
 sky130_fd_sc_hd__dfstp_1 merge913 (.CLK(clknet_4_5_0_clk),
    .D(net63),
    .Q(net64));
 sky130_fd_sc_hd__dfstp_1 merge914 (.CLK(clknet_4_14_0_clk),
    .D(net581),
    .SET_B(net582),
    .Q(net883));
 sky130_fd_sc_hd__dlrbn_1 merge915 (.D(net534),
    .GATE_N(clknet_4_10_0_clk),
    .RESET_B(net1060),
    .Q(net885),
    .Q_N(net884));
 sky130_fd_sc_hd__xnor2_1 merge916 (.A(net485),
    .B(net492),
    .Y(net886));
 sky130_fd_sc_hd__xnor2_1 merge917 (.A(net372),
    .B(net379),
    .Y(net887));
 sky130_fd_sc_hd__dlrbn_1 merge918 (.D(net245),
    .GATE_N(clknet_4_2_0_clk),
    .RESET_B(net238),
    .Q(net889),
    .Q_N(net888));
 sky130_fd_sc_hd__xnor2_1 merge919 (.A(net268),
    .B(net270),
    .Y(net890));
 sky130_fd_sc_hd__dlrbp_1 merge920 (.D(net595),
    .GATE(clknet_4_13_0_clk),
    .RESET_B(net598),
    .Q(net892),
    .Q_N(net891));
 sky130_fd_sc_hd__xnor2_1 merge921 (.A(net438),
    .B(net450),
    .Y(net893));
 sky130_fd_sc_hd__xnor2_1 merge922 (.A(net863),
    .B(net18),
    .Y(net894));
 sky130_fd_sc_hd__xnor2_1 merge923 (.A(net584),
    .B(net495),
    .Y(net895));
 sky130_fd_sc_hd__xnor2_1 merge924 (.A(net469),
    .B(net472),
    .Y(net896));
 sky130_fd_sc_hd__xnor2_1 merge925 (.A(net202),
    .B(net204),
    .Y(net897));
 sky130_fd_sc_hd__xnor2_1 merge926 (.A(net494),
    .B(net224),
    .Y(net898));
 sky130_fd_sc_hd__xnor2_1 merge927 (.A(net291),
    .B(net271),
    .Y(net899));
 sky130_fd_sc_hd__dlrbp_1 merge928 (.D(net225),
    .GATE(clknet_4_4_0_clk),
    .RESET_B(net833),
    .Q(net901),
    .Q_N(net900));
 sky130_fd_sc_hd__dlrtn_2 merge929 (.D(net817),
    .GATE_N(clknet_4_2_0_clk),
    .RESET_B(net820),
    .Q(net902));
 sky130_fd_sc_hd__xnor2_1 merge930 (.A(net355),
    .B(net383),
    .Y(net903));
 sky130_fd_sc_hd__dlrtn_1 merge931 (.D(net172),
    .GATE_N(clknet_4_7_0_clk),
    .RESET_B(net755),
    .Q(net904));
 sky130_fd_sc_hd__dlrtn_1 merge932 (.D(net814),
    .GATE_N(clknet_4_11_0_clk),
    .RESET_B(net880),
    .Q(net905));
 sky130_fd_sc_hd__dlrtp_1 merge933 (.D(net292),
    .GATE(clknet_4_15_0_clk),
    .RESET_B(net744),
    .Q(net906));
 sky130_fd_sc_hd__dlrtp_1 merge934 (.D(net860),
    .GATE(clknet_4_7_0_clk),
    .RESET_B(net745),
    .Q(net907));
 sky130_fd_sc_hd__dlrtp_1 merge935 (.D(net823),
    .GATE(clknet_4_13_0_clk),
    .RESET_B(net772),
    .Q(net908));
 sky130_fd_sc_hd__edfxbp_1 merge936 (.CLK(clknet_4_0_0_clk),
    .D(net746),
    .DE(net768),
    .Q(net910),
    .Q_N(net909));
 sky130_fd_sc_hd__edfxtp_1 merge937 (.CLK(clknet_4_11_0_clk),
    .D(net750),
    .DE(net822),
    .Q(net911));
 sky130_fd_sc_hd__sdlclkp_1 merge938 (.CLK(clknet_4_3_0_clk),
    .GATE(net28),
    .SCE(net32),
    .GCLK(net912));
 sky130_fd_sc_hd__xnor2_1 merge939 (.A(net512),
    .B(net513),
    .Y(net913));
 sky130_fd_sc_hd__sdlclkp_2 merge940 (.CLK(clknet_4_10_0_clk),
    .GATE(net854),
    .SCE(net535),
    .GCLK(net914));
 sky130_fd_sc_hd__sdlclkp_4 merge941 (.CLK(clknet_4_13_0_clk),
    .GATE(net780),
    .SCE(net831),
    .GCLK(net915));
 sky130_fd_sc_hd__dfrbp_1 merge942 (.CLK(clknet_4_6_0_clk),
    .D(net815),
    .RESET_B(net784),
    .Q(net917),
    .Q_N(net916));
 sky130_fd_sc_hd__xnor2_1 merge943 (.A(net514),
    .B(net913),
    .Y(net918));
 sky130_fd_sc_hd__dfrbp_1 merge944 (.CLK(clknet_4_11_0_clk),
    .D(net749),
    .RESET_B(net800),
    .Q(net920),
    .Q_N(net919));
 sky130_fd_sc_hd__dfrtn_1 merge945 (.CLK_N(clknet_4_15_0_clk),
    .D(net557),
    .RESET_B(net560),
    .Q(net921));
 sky130_fd_sc_hd__dfrtp_2 merge946 (.CLK(clknet_4_12_0_clk),
    .D(net515),
    .RESET_B(net791),
    .Q(net922));
 sky130_fd_sc_hd__dfrtp_1 merge947 (.CLK(clknet_4_3_0_clk),
    .D(net797),
    .RESET_B(net834),
    .Q(net923));
 sky130_fd_sc_hd__dfrtp_2 merge948 (.CLK(clknet_4_10_0_clk),
    .D(net862),
    .RESET_B(net1038),
    .Q(net924));
 sky130_fd_sc_hd__dfsbp_1 merge949 (.CLK(clknet_4_15_0_clk),
    .D(net798),
    .SET_B(net1050),
    .Q(net926),
    .Q_N(net925));
 sky130_fd_sc_hd__dfsbp_1 merge950 (.CLK(clknet_4_0_0_clk),
    .D(net816),
    .SET_B(net39),
    .Q(net928),
    .Q_N(net927));
 sky130_fd_sc_hd__dfstp_1 merge951 (.CLK(clknet_4_4_0_clk),
    .D(net836),
    .SET_B(net16),
    .Q(net929));
 sky130_fd_sc_hd__dfstp_1 merge952 (.CLK(clknet_4_5_0_clk),
    .D(net765),
    .SET_B(net742),
    .Q(net930));
 sky130_fd_sc_hd__dfstp_1 merge953 (.CLK(clknet_4_2_0_clk),
    .D(net887),
    .SET_B(net766),
    .Q(net931));
 sky130_fd_sc_hd__dlrbn_1 merge954 (.D(net774),
    .GATE_N(clknet_4_12_0_clk),
    .RESET_B(net849),
    .Q(net933),
    .Q_N(net932));
 sky130_fd_sc_hd__dlrbn_1 merge955 (.D(net821),
    .GATE_N(clknet_4_3_0_clk),
    .RESET_B(net748),
    .Q(net935),
    .Q_N(net934));
 sky130_fd_sc_hd__dlrbp_1 merge956 (.D(net830),
    .GATE(clknet_4_2_0_clk),
    .RESET_B(net839),
    .Q(net937),
    .Q_N(net936));
 sky130_fd_sc_hd__dlrbp_1 merge957 (.D(net896),
    .GATE(clknet_4_7_0_clk),
    .RESET_B(net155),
    .Q(net939),
    .Q_N(net938));
 sky130_fd_sc_hd__dlrtn_1 merge958 (.D(net845),
    .GATE_N(clknet_4_9_0_clk),
    .RESET_B(net852),
    .Q(net940));
 sky130_fd_sc_hd__dlrtn_2 merge959 (.D(net853),
    .GATE_N(clknet_4_14_0_clk),
    .RESET_B(net851),
    .Q(net941));
 sky130_fd_sc_hd__dlrtn_2 merge960 (.D(net789),
    .GATE_N(clknet_4_5_0_clk),
    .RESET_B(net898),
    .Q(net942));
 sky130_fd_sc_hd__dlrtp_1 merge961 (.D(net886),
    .GATE(clknet_4_14_0_clk),
    .RESET_B(net799),
    .Q(net943));
 sky130_fd_sc_hd__dlrtp_2 merge962 (.D(net835),
    .GATE(clknet_4_6_0_clk),
    .RESET_B(net795),
    .Q(net944));
 sky130_fd_sc_hd__dlrtp_2 merge963 (.D(net370),
    .GATE(clknet_4_3_0_clk),
    .RESET_B(net786),
    .Q(net945));
 sky130_fd_sc_hd__edfxbp_1 merge964 (.CLK(clknet_4_13_0_clk),
    .D(net782),
    .DE(net890),
    .Q(net947),
    .Q_N(net946));
 sky130_fd_sc_hd__edfxtp_1 merge965 (.CLK(clknet_4_1_0_clk),
    .D(net743),
    .DE(net41),
    .Q(net948));
 sky130_fd_sc_hd__sdlclkp_1 merge966 (.CLK(clknet_4_9_0_clk),
    .GATE(net698),
    .SCE(net842),
    .GCLK(net949));
 sky130_fd_sc_hd__sdlclkp_2 merge967 (.CLK(clknet_4_6_0_clk),
    .GATE(net850),
    .SCE(net805),
    .GCLK(net950));
 sky130_fd_sc_hd__sdlclkp_4 merge968 (.CLK(clknet_4_4_0_clk),
    .GATE(net826),
    .SCE(net770),
    .GCLK(net951));
 sky130_fd_sc_hd__dfrbp_1 merge969 (.CLK(clknet_4_11_0_clk),
    .D(net857),
    .RESET_B(net537),
    .Q(net953),
    .Q_N(net952));
 sky130_fd_sc_hd__dfrbp_1 merge970 (.CLK(clknet_4_5_0_clk),
    .D(net796),
    .RESET_B(net894),
    .Q(net955),
    .Q_N(net954));
 sky130_fd_sc_hd__dfrtn_1 merge971 (.CLK_N(clknet_4_7_0_clk),
    .D(net899),
    .RESET_B(net897),
    .Q(net956));
 sky130_fd_sc_hd__dfrtp_4 merge972 (.CLK(clknet_4_9_0_clk),
    .D(net449),
    .RESET_B(net846),
    .Q(net957));
 sky130_fd_sc_hd__dfrtp_2 merge973 (.CLK(clknet_4_12_0_clk),
    .D(net779),
    .RESET_B(net918),
    .Q(net958));
 sky130_fd_sc_hd__dfrtp_4 merge974 (.CLK(clknet_4_1_0_clk),
    .D(net869),
    .RESET_B(net1040),
    .Q(net959));
 sky130_fd_sc_hd__dfsbp_1 merge975 (.CLK(clknet_4_11_0_clk),
    .D(net801),
    .SET_B(net865),
    .Q(net961),
    .Q_N(net960));
 sky130_fd_sc_hd__dfsbp_1 merge976 (.CLK(clknet_4_4_0_clk),
    .D(net77),
    .SET_B(net874),
    .Q(net963),
    .Q_N(net962));
 sky130_fd_sc_hd__dfstp_1 merge977 (.CLK(clknet_4_11_0_clk),
    .D(net810),
    .SET_B(net844),
    .Q(net964));
 sky130_fd_sc_hd__dfstp_1 merge978 (.CLK(clknet_4_12_0_clk),
    .D(net859),
    .SET_B(net881),
    .Q(net965));
 sky130_fd_sc_hd__dfstp_1 merge979 (.CLK(clknet_4_12_0_clk),
    .D(net804),
    .SET_B(net806),
    .Q(net966));
 sky130_fd_sc_hd__dlrbn_1 merge980 (.D(net695),
    .GATE_N(clknet_4_9_0_clk),
    .RESET_B(net790),
    .Q(net968),
    .Q_N(net967));
 sky130_fd_sc_hd__dlrbn_1 merge981 (.D(net893),
    .GATE_N(clknet_4_11_0_clk),
    .RESET_B(net713),
    .Q(net970),
    .Q_N(net969));
 sky130_fd_sc_hd__dlrbp_1 merge982 (.D(net763),
    .GATE(clknet_4_14_0_clk),
    .RESET_B(net829),
    .Q(net972),
    .Q_N(net971));
 sky130_fd_sc_hd__dlrbp_1 merge983 (.D(net812),
    .GATE(clknet_4_7_0_clk),
    .RESET_B(net848),
    .Q(net974),
    .Q_N(net973));
 sky130_fd_sc_hd__dlrtn_2 merge984 (.D(net583),
    .GATE_N(clknet_4_13_0_clk),
    .RESET_B(net754),
    .Q(net975));
 sky130_fd_sc_hd__dlrtn_1 merge985 (.D(net840),
    .GATE_N(clknet_4_7_0_clk),
    .RESET_B(net813),
    .Q(net976));
 sky130_fd_sc_hd__dlrtn_2 merge986 (.D(net864),
    .GATE_N(clknet_4_13_0_clk),
    .RESET_B(net1046),
    .Q(net977));
 sky130_fd_sc_hd__dlrtp_1 merge987 (.D(net895),
    .GATE(clknet_4_9_0_clk),
    .RESET_B(net794),
    .Q(net978));
 sky130_fd_sc_hd__dlrtp_1 merge988 (.D(net877),
    .GATE(clknet_4_7_0_clk),
    .RESET_B(net858),
    .Q(net979));
 sky130_fd_sc_hd__dlrtp_2 merge989 (.D(net838),
    .GATE(clknet_4_1_0_clk),
    .RESET_B(net847),
    .Q(net980));
 sky130_fd_sc_hd__edfxbp_1 merge990 (.CLK(clknet_4_1_0_clk),
    .D(net811),
    .DE(net825),
    .Q(net982),
    .Q_N(net981));
 sky130_fd_sc_hd__edfxtp_1 merge991 (.CLK(clknet_4_3_0_clk),
    .D(net866),
    .DE(net837),
    .Q(net983));
 sky130_fd_sc_hd__sdlclkp_1 merge992 (.CLK(clknet_4_5_0_clk),
    .GATE(net903),
    .SCE(net832),
    .GCLK(net984));
 sky130_fd_sc_hd__sdlclkp_2 merge993 (.CLK(clknet_4_1_0_clk),
    .GATE(net861),
    .SCE(net828),
    .GCLK(net985));
 sky130_fd_sc_hd__dlclkp_2 s1000 (.CLK(clknet_4_9_0_clk),
    .GATE(net693),
    .GCLK(net993));
 sky130_fd_sc_hd__dlclkp_4 s1001 (.CLK(clknet_4_15_0_clk),
    .GATE(net841),
    .GCLK(net994));
 sky130_fd_sc_hd__dfxbp_1 s994 (.CLK(clknet_4_1_0_clk),
    .D(net82),
    .Q(net987),
    .Q_N(net986));
 sky130_fd_sc_hd__dfxbp_1 s995 (.CLK(clknet_4_2_0_clk),
    .D(net246),
    .Q(net989),
    .Q_N(net988));
 sky130_fd_sc_hd__dfxtp_2 s996 (.CLK(clknet_4_7_0_clk),
    .D(net314),
    .Q(net990));
 sky130_fd_sc_hd__dfxtp_1 s997 (.CLK(clknet_4_9_0_clk),
    .D(net427),
    .Q(net991));
 sky130_fd_sc_hd__dfxtp_1 s998 (.CLK(clknet_4_13_0_clk),
    .D(net604),
    .Q(net992));
 sky130_fd_sc_hd__dlclkp_1 s999 (.CLK(clknet_4_15_0_clk),
    .GATE(net629),
    .GCLK(net1020));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Right_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Right_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Right_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Right_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Right_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Right_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Right_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Right_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Right_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Right_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Right_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Right_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Right_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Right_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Right_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Right_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Right_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Right_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Right_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Right_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Right_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_161 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_162 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_163 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_164 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_165 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_166 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_167 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_168 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_169 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_170 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_171 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_172 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_173 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_174 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_175 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_176 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_177 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_178 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_179 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_180 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_181 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_182 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Left_183 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Left_184 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Left_185 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Left_186 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Left_187 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Left_188 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Left_189 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Left_190 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Left_191 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Left_192 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Left_193 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Left_194 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Left_195 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Left_196 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Left_197 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Left_198 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Left_199 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Left_200 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Left_201 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Left_202 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Left_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1347 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(in0),
    .X(net556));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(in1),
    .X(net628));
 sky130_fd_sc_hd__buf_1 input3 (.A(in10),
    .X(net759));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(in11),
    .X(net995));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(in12),
    .X(net996));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(in13),
    .X(net997));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(in14),
    .X(net998));
 sky130_fd_sc_hd__clkbuf_2 input8 (.A(in15),
    .X(net999));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(in16),
    .X(net1000));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(in17),
    .X(net1001));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(in19),
    .X(net1002));
 sky130_fd_sc_hd__buf_1 input12 (.A(in2),
    .X(net1003));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(in20),
    .X(net1004));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(in21),
    .X(net1005));
 sky130_fd_sc_hd__buf_4 input15 (.A(in22),
    .X(net1006));
 sky130_fd_sc_hd__buf_1 input16 (.A(in23),
    .X(net1007));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(in24),
    .X(net1008));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(in3),
    .X(net1009));
 sky130_fd_sc_hd__buf_1 input19 (.A(in4),
    .X(net1010));
 sky130_fd_sc_hd__clkbuf_1 input20 (.A(in5),
    .X(net1011));
 sky130_fd_sc_hd__buf_1 input21 (.A(in6),
    .X(net1012));
 sky130_fd_sc_hd__buf_1 input22 (.A(in7),
    .X(net1013));
 sky130_fd_sc_hd__clkbuf_1 input23 (.A(in8),
    .X(net1014));
 sky130_fd_sc_hd__buf_1 input24 (.A(in9),
    .X(net1015));
 sky130_fd_sc_hd__clkbuf_4 output25 (.A(net1016),
    .X(out0));
 sky130_fd_sc_hd__clkbuf_4 output26 (.A(net1017),
    .X(out1));
 sky130_fd_sc_hd__clkbuf_1 output27 (.A(net1018),
    .X(out12));
 sky130_fd_sc_hd__clkbuf_4 output28 (.A(net1019),
    .X(out13));
 sky130_fd_sc_hd__clkbuf_1 output29 (.A(clknet_1_1__leaf_net1020),
    .X(out14));
 sky130_fd_sc_hd__clkbuf_4 output30 (.A(net1021),
    .X(out16));
 sky130_fd_sc_hd__clkbuf_4 output31 (.A(net1022),
    .X(out19));
 sky130_fd_sc_hd__clkbuf_4 output32 (.A(net1023),
    .X(out21));
 sky130_fd_sc_hd__clkbuf_4 output33 (.A(net1024),
    .X(out22));
 sky130_fd_sc_hd__clkbuf_4 output34 (.A(net1025),
    .X(out23));
 sky130_fd_sc_hd__clkbuf_4 output35 (.A(net1026),
    .X(out24));
 sky130_fd_sc_hd__clkbuf_4 output36 (.A(net1027),
    .X(out4));
 sky130_fd_sc_hd__clkbuf_4 output37 (.A(net1028),
    .X(out5));
 sky130_fd_sc_hd__clkbuf_4 output38 (.A(net1029),
    .X(out7));
 sky130_fd_sc_hd__clkbuf_4 output39 (.A(net1030),
    .X(out9));
 sky130_fd_sc_hd__buf_4 max_cap40 (.A(net722),
    .X(net1031));
 sky130_fd_sc_hd__buf_4 max_cap41 (.A(net411),
    .X(net1032));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net1020 (.A(net1020),
    .X(clknet_0_net1020));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net1020 (.A(clknet_0_net1020),
    .X(clknet_1_0__leaf_net1020));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net1020 (.A(clknet_0_net1020),
    .X(clknet_1_1__leaf_net1020));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net994 (.A(net994),
    .X(clknet_0_net994));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net994 (.A(clknet_0_net994),
    .X(clknet_1_0__leaf_net994));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net994 (.A(clknet_0_net994),
    .X(clknet_1_1__leaf_net994));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net558 (.A(net558),
    .X(clknet_0_net558));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net558 (.A(clknet_0_net558),
    .X(clknet_1_0__leaf_net558));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net558 (.A(clknet_0_net558),
    .X(clknet_1_1__leaf_net558));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net563 (.A(net563),
    .X(clknet_0_net563));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net563 (.A(clknet_0_net563),
    .X(clknet_1_0__leaf_net563));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net563 (.A(clknet_0_net563),
    .X(clknet_1_1__leaf_net563));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net993 (.A(net993),
    .X(clknet_0_net993));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net993 (.A(clknet_0_net993),
    .X(clknet_1_0__leaf_net993));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net993 (.A(clknet_0_net993),
    .X(clknet_1_1__leaf_net993));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net694 (.A(net694),
    .X(clknet_0_net694));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net694 (.A(clknet_0_net694),
    .X(clknet_1_0__leaf_net694));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net694 (.A(clknet_0_net694),
    .X(clknet_1_1__leaf_net694));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net949 (.A(net949),
    .X(clknet_0_net949));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net949 (.A(clknet_0_net949),
    .X(clknet_1_0__leaf_net949));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net949 (.A(clknet_0_net949),
    .X(clknet_1_1__leaf_net949));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net710 (.A(net710),
    .X(clknet_0_net710));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net710 (.A(clknet_0_net710),
    .X(clknet_1_0__leaf_net710));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net710 (.A(clknet_0_net710),
    .X(clknet_1_1__leaf_net710));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net717 (.A(net717),
    .X(clknet_0_net717));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net717 (.A(clknet_0_net717),
    .X(clknet_1_0__leaf_net717));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net717 (.A(clknet_0_net717),
    .X(clknet_1_1__leaf_net717));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net719 (.A(net719),
    .X(clknet_0_net719));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net719 (.A(clknet_0_net719),
    .X(clknet_1_0__leaf_net719));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net719 (.A(clknet_0_net719),
    .X(clknet_1_1__leaf_net719));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net712 (.A(net712),
    .X(clknet_0_net712));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net712 (.A(clknet_0_net712),
    .X(clknet_1_0__leaf_net712));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net712 (.A(clknet_0_net712),
    .X(clknet_1_1__leaf_net712));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net442 (.A(net442),
    .X(clknet_0_net442));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net442 (.A(clknet_0_net442),
    .X(clknet_1_0__leaf_net442));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net442 (.A(clknet_0_net442),
    .X(clknet_1_1__leaf_net442));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net447 (.A(net447),
    .X(clknet_0_net447));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net447 (.A(clknet_0_net447),
    .X(clknet_1_0__leaf_net447));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net447 (.A(clknet_0_net447),
    .X(clknet_1_1__leaf_net447));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net914 (.A(net914),
    .X(clknet_0_net914));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net914 (.A(clknet_0_net914),
    .X(clknet_1_0__leaf_net914));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net914 (.A(clknet_0_net914),
    .X(clknet_1_1__leaf_net914));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net985 (.A(net985),
    .X(clknet_0_net985));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net985 (.A(clknet_0_net985),
    .X(clknet_1_0__leaf_net985));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net985 (.A(clknet_0_net985),
    .X(clknet_1_1__leaf_net985));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net984 (.A(net984),
    .X(clknet_0_net984));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net984 (.A(clknet_0_net984),
    .X(clknet_1_0__leaf_net984));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net984 (.A(clknet_0_net984),
    .X(clknet_1_1__leaf_net984));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net498 (.A(net498),
    .X(clknet_0_net498));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net498 (.A(clknet_0_net498),
    .X(clknet_1_0__leaf_net498));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net498 (.A(clknet_0_net498),
    .X(clknet_1_1__leaf_net498));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net357 (.A(net357),
    .X(clknet_0_net357));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net357 (.A(clknet_0_net357),
    .X(clknet_1_0__leaf_net357));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net357 (.A(clknet_0_net357),
    .X(clknet_1_1__leaf_net357));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net197 (.A(net197),
    .X(clknet_0_net197));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net197 (.A(clknet_0_net197),
    .X(clknet_1_0__leaf_net197));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net197 (.A(clknet_0_net197),
    .X(clknet_1_1__leaf_net197));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net201 (.A(net201),
    .X(clknet_0_net201));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net201 (.A(clknet_0_net201),
    .X(clknet_1_0__leaf_net201));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net201 (.A(clknet_0_net201),
    .X(clknet_1_1__leaf_net201));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net85 (.A(net85),
    .X(clknet_0_net85));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net85 (.A(clknet_0_net85),
    .X(clknet_1_0__leaf_net85));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net85 (.A(clknet_0_net85),
    .X(clknet_1_1__leaf_net85));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net205 (.A(net205),
    .X(clknet_0_net205));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net205 (.A(clknet_0_net205),
    .X(clknet_1_0__leaf_net205));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net205 (.A(clknet_0_net205),
    .X(clknet_1_1__leaf_net205));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net208 (.A(net208),
    .X(clknet_0_net208));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net208 (.A(clknet_0_net208),
    .X(clknet_1_0__leaf_net208));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net208 (.A(clknet_0_net208),
    .X(clknet_1_1__leaf_net208));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net226 (.A(net226),
    .X(clknet_0_net226));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net226 (.A(clknet_0_net226),
    .X(clknet_1_0__leaf_net226));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net226 (.A(clknet_0_net226),
    .X(clknet_1_1__leaf_net226));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net210 (.A(net210),
    .X(clknet_0_net210));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net210 (.A(clknet_0_net210),
    .X(clknet_1_0__leaf_net210));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net210 (.A(clknet_0_net210),
    .X(clknet_1_1__leaf_net210));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net207 (.A(net207),
    .X(clknet_0_net207));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net207 (.A(clknet_0_net207),
    .X(clknet_1_0__leaf_net207));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net207 (.A(clknet_0_net207),
    .X(clknet_1_1__leaf_net207));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net213 (.A(net213),
    .X(clknet_0_net213));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net213 (.A(clknet_0_net213),
    .X(clknet_1_0__leaf_net213));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net213 (.A(clknet_0_net213),
    .X(clknet_1_1__leaf_net213));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net87 (.A(net87),
    .X(clknet_0_net87));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net87 (.A(clknet_0_net87),
    .X(clknet_1_0__leaf_net87));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net87 (.A(clknet_0_net87),
    .X(clknet_1_1__leaf_net87));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net91 (.A(net91),
    .X(clknet_0_net91));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net91 (.A(clknet_0_net91),
    .X(clknet_1_0__leaf_net91));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net91 (.A(clknet_0_net91),
    .X(clknet_1_1__leaf_net91));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net89 (.A(net89),
    .X(clknet_0_net89));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net89 (.A(clknet_0_net89),
    .X(clknet_1_0__leaf_net89));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net89 (.A(clknet_0_net89),
    .X(clknet_1_1__leaf_net89));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net88 (.A(net88),
    .X(clknet_0_net88));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net88 (.A(clknet_0_net88),
    .X(clknet_1_0__leaf_net88));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net88 (.A(clknet_0_net88),
    .X(clknet_1_1__leaf_net88));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net95 (.A(net95),
    .X(clknet_0_net95));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net95 (.A(clknet_0_net95),
    .X(clknet_1_0__leaf_net95));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net95 (.A(clknet_0_net95),
    .X(clknet_1_1__leaf_net95));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net79 (.A(net79),
    .X(clknet_0_net79));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net79 (.A(clknet_0_net79),
    .X(clknet_1_0__leaf_net79));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net79 (.A(clknet_0_net79),
    .X(clknet_1_1__leaf_net79));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net81 (.A(net81),
    .X(clknet_0_net81));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net81 (.A(clknet_0_net81),
    .X(clknet_1_0__leaf_net81));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net81 (.A(clknet_0_net81),
    .X(clknet_1_1__leaf_net81));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net951 (.A(net951),
    .X(clknet_0_net951));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net951 (.A(clknet_0_net951),
    .X(clknet_1_0__leaf_net951));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net951 (.A(clknet_0_net951),
    .X(clknet_1_1__leaf_net951));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net42 (.A(net42),
    .X(clknet_0_net42));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net42 (.A(clknet_0_net42),
    .X(clknet_1_0__leaf_net42));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net42 (.A(clknet_0_net42),
    .X(clknet_1_1__leaf_net42));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net29 (.A(net29),
    .X(clknet_0_net29));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net29 (.A(clknet_0_net29),
    .X(clknet_1_0__leaf_net29));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net29 (.A(clknet_0_net29),
    .X(clknet_1_1__leaf_net29));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net912 (.A(net912),
    .X(clknet_0_net912));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net912 (.A(clknet_0_net912),
    .X(clknet_1_0__leaf_net912));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net912 (.A(clknet_0_net912),
    .X(clknet_1_1__leaf_net912));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net26 (.A(net26),
    .X(clknet_0_net26));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net26 (.A(clknet_0_net26),
    .X(clknet_1_0__leaf_net26));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net26 (.A(clknet_0_net26),
    .X(clknet_1_1__leaf_net26));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net21 (.A(net21),
    .X(clknet_0_net21));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net21 (.A(clknet_0_net21),
    .X(clknet_1_0__leaf_net21));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net21 (.A(clknet_0_net21),
    .X(clknet_1_1__leaf_net21));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net24 (.A(net24),
    .X(clknet_0_net24));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net24 (.A(clknet_0_net24),
    .X(clknet_1_0__leaf_net24));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net24 (.A(clknet_0_net24),
    .X(clknet_1_1__leaf_net24));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net20 (.A(net20),
    .X(clknet_0_net20));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net20 (.A(clknet_0_net20),
    .X(clknet_1_0__leaf_net20));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net20 (.A(clknet_0_net20),
    .X(clknet_1_1__leaf_net20));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net25 (.A(net25),
    .X(clknet_0_net25));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net25 (.A(clknet_0_net25),
    .X(clknet_1_0__leaf_net25));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net25 (.A(clknet_0_net25),
    .X(clknet_1_1__leaf_net25));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net23 (.A(net23),
    .X(clknet_0_net23));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net23 (.A(clknet_0_net23),
    .X(clknet_1_0__leaf_net23));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net23 (.A(clknet_0_net23),
    .X(clknet_1_1__leaf_net23));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net34 (.A(net34),
    .X(clknet_0_net34));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net34 (.A(clknet_0_net34),
    .X(clknet_1_0__leaf_net34));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net34 (.A(clknet_0_net34),
    .X(clknet_1_1__leaf_net34));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net161 (.A(net161),
    .X(clknet_0_net161));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net161 (.A(clknet_0_net161),
    .X(clknet_1_0__leaf_net161));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net161 (.A(clknet_0_net161),
    .X(clknet_1_1__leaf_net161));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net163 (.A(net163),
    .X(clknet_0_net163));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net163 (.A(clknet_0_net163),
    .X(clknet_1_0__leaf_net163));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net163 (.A(clknet_0_net163),
    .X(clknet_1_1__leaf_net163));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net168 (.A(net168),
    .X(clknet_0_net168));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net168 (.A(clknet_0_net168),
    .X(clknet_1_0__leaf_net168));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net168 (.A(clknet_0_net168),
    .X(clknet_1_1__leaf_net168));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net162 (.A(net162),
    .X(clknet_0_net162));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net162 (.A(clknet_0_net162),
    .X(clknet_1_0__leaf_net162));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net162 (.A(clknet_0_net162),
    .X(clknet_1_1__leaf_net162));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net27 (.A(net27),
    .X(clknet_0_net27));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net27 (.A(clknet_0_net27),
    .X(clknet_1_0__leaf_net27));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net27 (.A(clknet_0_net27),
    .X(clknet_1_1__leaf_net27));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net22 (.A(net22),
    .X(clknet_0_net22));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net22 (.A(clknet_0_net22),
    .X(clknet_1_0__leaf_net22));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net22 (.A(clknet_0_net22),
    .X(clknet_1_1__leaf_net22));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net352 (.A(net352),
    .X(clknet_0_net352));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net352 (.A(clknet_0_net352),
    .X(clknet_1_0__leaf_net352));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net352 (.A(clknet_0_net352),
    .X(clknet_1_1__leaf_net352));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net353 (.A(net353),
    .X(clknet_0_net353));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net353 (.A(clknet_0_net353),
    .X(clknet_1_0__leaf_net353));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net353 (.A(clknet_0_net353),
    .X(clknet_1_1__leaf_net353));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net950 (.A(net950),
    .X(clknet_0_net950));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net950 (.A(clknet_0_net950),
    .X(clknet_1_0__leaf_net950));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net950 (.A(clknet_0_net950),
    .X(clknet_1_1__leaf_net950));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net764 (.A(net764),
    .X(clknet_0_net764));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net764 (.A(clknet_0_net764),
    .X(clknet_1_0__leaf_net764));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net764 (.A(clknet_0_net764),
    .X(clknet_1_1__leaf_net764));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net482 (.A(net482),
    .X(clknet_0_net482));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net482 (.A(clknet_0_net482),
    .X(clknet_1_0__leaf_net482));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net482 (.A(clknet_0_net482),
    .X(clknet_1_1__leaf_net482));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net479 (.A(net479),
    .X(clknet_0_net479));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net479 (.A(clknet_0_net479),
    .X(clknet_1_0__leaf_net479));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net479 (.A(clknet_0_net479),
    .X(clknet_1_1__leaf_net479));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net491 (.A(net491),
    .X(clknet_0_net491));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net491 (.A(clknet_0_net491),
    .X(clknet_1_0__leaf_net491));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net491 (.A(clknet_0_net491),
    .X(clknet_1_1__leaf_net491));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net496 (.A(net496),
    .X(clknet_0_net496));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net496 (.A(clknet_0_net496),
    .X(clknet_1_0__leaf_net496));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net496 (.A(clknet_0_net496),
    .X(clknet_1_1__leaf_net496));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net493 (.A(net493),
    .X(clknet_0_net493));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net493 (.A(clknet_0_net493),
    .X(clknet_1_0__leaf_net493));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net493 (.A(clknet_0_net493),
    .X(clknet_1_1__leaf_net493));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net747 (.A(net747),
    .X(clknet_0_net747));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net747 (.A(clknet_0_net747),
    .X(clknet_1_0__leaf_net747));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net747 (.A(clknet_0_net747),
    .X(clknet_1_1__leaf_net747));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net318 (.A(net318),
    .X(clknet_0_net318));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net318 (.A(clknet_0_net318),
    .X(clknet_1_0__leaf_net318));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net318 (.A(clknet_0_net318),
    .X(clknet_1_1__leaf_net318));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net325 (.A(net325),
    .X(clknet_0_net325));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net325 (.A(clknet_0_net325),
    .X(clknet_1_0__leaf_net325));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net325 (.A(clknet_0_net325),
    .X(clknet_1_1__leaf_net325));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net320 (.A(net320),
    .X(clknet_0_net320));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net320 (.A(clknet_0_net320),
    .X(clknet_1_0__leaf_net320));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net320 (.A(clknet_0_net320),
    .X(clknet_1_1__leaf_net320));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net321 (.A(net321),
    .X(clknet_0_net321));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net321 (.A(clknet_0_net321),
    .X(clknet_1_0__leaf_net321));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net321 (.A(clknet_0_net321),
    .X(clknet_1_1__leaf_net321));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net317 (.A(net317),
    .X(clknet_0_net317));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net317 (.A(clknet_0_net317),
    .X(clknet_1_0__leaf_net317));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net317 (.A(clknet_0_net317),
    .X(clknet_1_1__leaf_net317));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net324 (.A(net324),
    .X(clknet_0_net324));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net324 (.A(clknet_0_net324),
    .X(clknet_1_0__leaf_net324));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net324 (.A(clknet_0_net324),
    .X(clknet_1_1__leaf_net324));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net329 (.A(net329),
    .X(clknet_0_net329));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net329 (.A(clknet_0_net329),
    .X(clknet_1_0__leaf_net329));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net329 (.A(clknet_0_net329),
    .X(clknet_1_1__leaf_net329));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net326 (.A(net326),
    .X(clknet_0_net326));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net326 (.A(clknet_0_net326),
    .X(clknet_1_0__leaf_net326));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net326 (.A(clknet_0_net326),
    .X(clknet_1_1__leaf_net326));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net330 (.A(net330),
    .X(clknet_0_net330));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net330 (.A(clknet_0_net330),
    .X(clknet_1_0__leaf_net330));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net330 (.A(clknet_0_net330),
    .X(clknet_1_1__leaf_net330));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net328 (.A(net328),
    .X(clknet_0_net328));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net328 (.A(clknet_0_net328),
    .X(clknet_1_0__leaf_net328));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net328 (.A(clknet_0_net328),
    .X(clknet_1_1__leaf_net328));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net915 (.A(net915),
    .X(clknet_0_net915));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net915 (.A(clknet_0_net915),
    .X(clknet_1_0__leaf_net915));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net915 (.A(clknet_0_net915),
    .X(clknet_1_1__leaf_net915));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net160 (.A(net160),
    .X(clknet_0_net160));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net160 (.A(clknet_0_net160),
    .X(clknet_1_0__leaf_net160));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net160 (.A(clknet_0_net160),
    .X(clknet_1_1__leaf_net160));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net144 (.A(net144),
    .X(clknet_0_net144));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net144 (.A(clknet_0_net144),
    .X(clknet_1_0__leaf_net144));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net144 (.A(clknet_0_net144),
    .X(clknet_1_1__leaf_net144));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net147 (.A(net147),
    .X(clknet_0_net147));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net147 (.A(clknet_0_net147),
    .X(clknet_1_0__leaf_net147));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net147 (.A(clknet_0_net147),
    .X(clknet_1_1__leaf_net147));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net145 (.A(net145),
    .X(clknet_0_net145));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net145 (.A(clknet_0_net145),
    .X(clknet_1_0__leaf_net145));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net145 (.A(clknet_0_net145),
    .X(clknet_1_1__leaf_net145));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net272 (.A(net272),
    .X(clknet_0_net272));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net272 (.A(clknet_0_net272),
    .X(clknet_1_0__leaf_net272));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net272 (.A(clknet_0_net272),
    .X(clknet_1_1__leaf_net272));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net126 (.A(net126),
    .X(clknet_0_net126));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net126 (.A(clknet_0_net126),
    .X(clknet_1_0__leaf_net126));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net126 (.A(clknet_0_net126),
    .X(clknet_1_1__leaf_net126));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net129 (.A(net129),
    .X(clknet_0_net129));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net129 (.A(clknet_0_net129),
    .X(clknet_1_0__leaf_net129));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net129 (.A(clknet_0_net129),
    .X(clknet_1_1__leaf_net129));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net127 (.A(net127),
    .X(clknet_0_net127));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net127 (.A(clknet_0_net127),
    .X(clknet_1_0__leaf_net127));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net127 (.A(clknet_0_net127),
    .X(clknet_1_1__leaf_net127));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer1 (.A(net902),
    .X(net1033));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer2 (.A(net902),
    .X(net1034));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer3 (.A(net33),
    .X(net1035));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(net102),
    .X(net1036));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(net530),
    .X(net1037));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(net536),
    .X(net1038));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(net980),
    .X(net1039));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(net114),
    .X(net1040));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(net969),
    .X(net1041));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(net222),
    .X(net1042));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(net824),
    .X(net1043));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(net962),
    .X(net1044));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(net992),
    .X(net1045));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(net607),
    .X(net1046));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(net228),
    .X(net1047));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(net952),
    .X(net1048));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(net792),
    .X(net1049));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(net843),
    .X(net1050));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(net99),
    .X(net1051));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(net105),
    .X(net1052));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(net807),
    .X(net1053));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(net1021),
    .X(net1054));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(net550),
    .X(net1056));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(net555),
    .X(net1057));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(net280),
    .X(net1058));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(net539),
    .X(net1060));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(net889),
    .X(net1061));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(net235),
    .X(net1062));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(net578),
    .X(net1063));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(net873),
    .X(net1064));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(net818),
    .X(net1065));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(net518),
    .X(net1066));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(net891),
    .X(net1067));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(net229),
    .X(net1068));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(net986),
    .X(net1069));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(net540),
    .X(net1070));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(net958),
    .X(net1071));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(net802),
    .X(net1072));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_A (.DIODE(clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(in0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(in1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(in10));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(in11));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(in12));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(in13));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(in14));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(in15));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(in16));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(in17));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_A (.DIODE(in18));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(in19));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(in2));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(in20));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(in21));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(in22));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(in23));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(in24));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(in3));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(in4));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(in5));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(in6));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_A (.DIODE(in7));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_A (.DIODE(in8));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_A (.DIODE(in9));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge872_S0 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge785_A1 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_c134_X (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge874_A3 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge872_S1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c140_X (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge860_A3 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge808_B1_N (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge794_B1 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge782_S1 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c59_SCD (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c42_A2 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c41_A3 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c38_B1 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c37_X (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_S0 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge883_S1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge874_S1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge872_A3 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_S0 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_A2 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_X (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge880_S1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge865_A3 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge818_A3 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge793_A2 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_A3 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_SET_B (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_Y (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge877_B1 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge812_A2 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_A (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_A3 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_B (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA_c286_A (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA_c283_A1 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_B1_N (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA_c278_X (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge884_A1 (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge840_A2 (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge824_A2 (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge822_A2 (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_S1 (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA_c323_S0 (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_Y (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge868_A2 (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge833_A1 (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_B1 (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_A (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_B1_N (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_X (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_S0 (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_B1_N (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_A0 (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_A3 (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_B1_N (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA_c346_X (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_A3 (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_B (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_A (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA_c373_X (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge881_A2 (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge870_S0 (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge861_DE (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge841_A1 (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA_c395_S1 (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA_c392_A4 (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA_c385_A3 (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA_c383_A1 (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA_c375_X (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge871_A1 (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge870_S1 (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge862_A2 (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge841_A2 (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA_c385_A2 (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA_c378_Y (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge814_A2 (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA_c507_B (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA_c394_Q_N (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA_c513_A2 (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA_c511_A (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA_c395_A3 (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA_c394_Q (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA_c404_B (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA_c403_A (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA_c397_A (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_X (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA_c563_B1_N (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_A (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA_c416_X (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge792_D (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_X (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge855_A1 (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_B (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_B (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_A (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_X (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_A3 (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_B1_N (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA_c431_A (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_A2 (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_B (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_B (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_B (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_A (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_X (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge859_B1 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge858_SCD (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge855_A2 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_A1 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_Y (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge853_SCD (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_B1_N (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_A (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_S0 (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_S0 (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_X (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge867_A1 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_c88_A (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_c70_B (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_c67_A (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_c66_X (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_A (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_c107_A2 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_c105_S1 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge853_SCE (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge828_B1 (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge821_A3 (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_A3 (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA_c446_Y (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge831_B1 (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_B1 (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_S1 (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_B (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_A2 (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_A1 (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_A (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_A (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_A2 (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_X (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge882_A1 (.DIODE(net509));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge869_A3 (.DIODE(net509));
 sky130_fd_sc_hd__diode_2 ANTENNA_c525_A2 (.DIODE(net509));
 sky130_fd_sc_hd__diode_2 ANTENNA_c523_A2 (.DIODE(net509));
 sky130_fd_sc_hd__diode_2 ANTENNA_c522_B1_N (.DIODE(net509));
 sky130_fd_sc_hd__diode_2 ANTENNA_c521_A1 (.DIODE(net509));
 sky130_fd_sc_hd__diode_2 ANTENNA_c519_Y (.DIODE(net509));
 sky130_fd_sc_hd__diode_2 ANTENNA_c657_S1 (.DIODE(net510));
 sky130_fd_sc_hd__diode_2 ANTENNA_c655_A1 (.DIODE(net510));
 sky130_fd_sc_hd__diode_2 ANTENNA_c654_A3 (.DIODE(net510));
 sky130_fd_sc_hd__diode_2 ANTENNA_c527_B1_N (.DIODE(net510));
 sky130_fd_sc_hd__diode_2 ANTENNA_c524_A2 (.DIODE(net510));
 sky130_fd_sc_hd__diode_2 ANTENNA_c521_B1_N (.DIODE(net510));
 sky130_fd_sc_hd__diode_2 ANTENNA_c520_X (.DIODE(net510));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge829_SCD (.DIODE(net523));
 sky130_fd_sc_hd__diode_2 ANTENNA_c541_A1 (.DIODE(net523));
 sky130_fd_sc_hd__diode_2 ANTENNA_c533_X (.DIODE(net523));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge829_D (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA_c543_A2 (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA_c538_D (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA_c534_Y (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge807_SCD (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA_c564_A2 (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA_c556_A (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA_c555_B (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA_c544_A2 (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA_c540_B1_N (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA_c539_SCD (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA_c535_X (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net563_A (.DIODE(net563));
 sky130_fd_sc_hd__diode_2 ANTENNA_c571_X (.DIODE(net563));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge879_A2 (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_A3 (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_A3 (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_B1_N (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_A1 (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_B (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_A (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_X (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge887_A2 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge846_A2 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge803_B1_N (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_c87_A3 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_c86_B1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_c80_X (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_c101_A1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge814_A0 (.DIODE(net589));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_A2 (.DIODE(net589));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_SCD (.DIODE(net589));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_Y (.DIODE(net589));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge817_A1 (.DIODE(net601));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_Y (.DIODE(net601));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge863_A1 (.DIODE(net669));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_A3 (.DIODE(net669));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_A2 (.DIODE(net669));
 sky130_fd_sc_hd__diode_2 ANTENNA_c698_B1_N (.DIODE(net669));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_X (.DIODE(net669));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge886_A0 (.DIODE(net676));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge863_B1_N (.DIODE(net676));
 sky130_fd_sc_hd__diode_2 ANTENNA_c703_X (.DIODE(net676));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge880_A2 (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge830_A2 (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA_c747_A3 (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA_c742_RESET_B (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_A (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_S0 (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_B (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_A2 (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_B (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_X (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A (.DIODE(net720));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_A (.DIODE(net720));
 sky130_fd_sc_hd__diode_2 ANTENNA_c747_A2 (.DIODE(net720));
 sky130_fd_sc_hd__diode_2 ANTENNA_c746_X (.DIODE(net720));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge964_D (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge820_X (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge959_D (.DIODE(net853));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge887_X (.DIODE(net853));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge971_D (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge927_Y (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge946_Q (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge869_S0 (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_A (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_A (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_c546_B1 (.DIODE(net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_c548_S1 (.DIODE(net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge948_Q (.DIODE(net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge852_B1 (.DIODE(net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_c703_B1 (.DIODE(net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge951_Q (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge799_A (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c42_A4 (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c41_S1 (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_A (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge959_Q (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c85_A (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c82_A (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_A (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_A (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge960_Q (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c513_B1_N (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c240_B1_N (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_A (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_A (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge961_Q (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge849_B1 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c586_A (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_B1 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_A (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge962_Q (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge815_A (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_c526_A (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_A (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_A (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge964_Q (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c194_A (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_A (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge972_Q (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_A (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_B (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_S1 (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_A (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold39_A (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge973_Q (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge869_S1 (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge805_A (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_A (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge982_Q_N (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_A (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_A (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge984_Q (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_A (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_B1 (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c159_A (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_A (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge985_Q (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_c77_A (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_A (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_A (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_c148_A (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge986_Q (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_B (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_B (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_B1 (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_S1 (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge988_Q (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge867_S1 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c62_B1 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_B1 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_B1_N (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold7_A (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge989_Q (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge809_A (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c382_A (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_A (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge991_Q (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c746_A (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c384_A (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c369_A (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_B (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_s996_Q (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge884_S1 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_B (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_B1 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_B1 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_s997_Q (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge801_B1_N (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_B (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_A (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_X (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge808_A2 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c56_A4 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c42_A3 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c37_B1_N (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c34_SCE (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c32_B1 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c27_B (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c25_B (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_A (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_X (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge880_A3 (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_output35_A (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c514_Y (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap41_X (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge883_A1 (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_B (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_A1 (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_A2 (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_B (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_A3 (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_A (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_15_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_14_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_13_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_12_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_11_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_10_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_9_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_8_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_7_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_6_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_5_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_4_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_3_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_2_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_1_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_0_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_X (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c121_CLK_N (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c122_CLK_N (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c123_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c124_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c125_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c127_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c129_CLK_N (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c250_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c254_CLK_N (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c255_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge936_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge950_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_0_0_clk_X (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c59_CLK_N (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge844_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge965_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge974_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge989_GATE (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge990_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge993_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s994_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_1_0_clk_X (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c494_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge889_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge907_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge942_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge962_GATE (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge967_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_6_0_clk_X (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge931_GATE_N (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge934_GATE (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge957_GATE (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge971_CLK_N (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge983_GATE (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge985_GATE_N (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge988_GATE (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s996_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_7_0_clk_X (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c767_CLK_N (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge932_GATE_N (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge937_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge944_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge969_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge975_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge977_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge981_GATE_N (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_11_0_clk_X (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c610_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge902_CLK_N (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge920_GATE (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge935_GATE (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge941_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge964_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge984_GATE_N (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge986_GATE_N (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s998_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_13_0_clk_X (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge797_SCD (.DIODE(clknet_1_0__leaf_net563));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge825_SCD (.DIODE(clknet_1_0__leaf_net563));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge852_A3 (.DIODE(clknet_1_0__leaf_net563));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net563_X (.DIODE(clknet_1_0__leaf_net563));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge836_A2 (.DIODE(clknet_1_1__leaf_net563));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge879_A1 (.DIODE(clknet_1_1__leaf_net563));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net563_X (.DIODE(clknet_1_1__leaf_net563));
 sky130_fd_sc_hd__diode_2 ANTENNA_c212_A (.DIODE(clknet_1_1__leaf_net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c508_B (.DIODE(clknet_1_1__leaf_net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net984_X (.DIODE(clknet_1_1__leaf_net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c286_B (.DIODE(clknet_1_0__leaf_net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge880_S0 (.DIODE(clknet_1_0__leaf_net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net145_X (.DIODE(clknet_1_0__leaf_net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(net140));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_478 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_379 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_242 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_260 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_490 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_364 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_482 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_228 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_271 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_466 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_366 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_275 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_548 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_428 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_527 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_539 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_520 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_479 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_441 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_535 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_543 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_566 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_546 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_548 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_608 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_354 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_507 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_538 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_599 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_336 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_504 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_582 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_554 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_508 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_532 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_385 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_187 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_403 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_476 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_532 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_547 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_283 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_584 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_274 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_411 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_566 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_395 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_245 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_392 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_494 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_506 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_518 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_267 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_283 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_327 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_423 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_522 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_387 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_536 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_467 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_395 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_439 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_617 ();
endmodule
