module netlist_1 (clk,
    in0,
    in1,
    in10,
    in11,
    in12,
    in13,
    in14,
    in15,
    in16,
    in17,
    in18,
    in19,
    in2,
    in20,
    in21,
    in22,
    in23,
    in24,
    in3,
    in4,
    in5,
    in6,
    in7,
    in8,
    in9,
    out0,
    out1,
    out10,
    out11,
    out12,
    out13,
    out14,
    out15,
    out16,
    out17,
    out18,
    out19,
    out2,
    out20,
    out21,
    out22,
    out23,
    out24,
    out3,
    out4,
    out5,
    out6,
    out7,
    out8,
    out9,
    rst);
 input clk;
 input in0;
 input in1;
 input in10;
 input in11;
 input in12;
 input in13;
 input in14;
 input in15;
 input in16;
 input in17;
 input in18;
 input in19;
 input in2;
 input in20;
 input in21;
 input in22;
 input in23;
 input in24;
 input in3;
 input in4;
 input in5;
 input in6;
 input in7;
 input in8;
 input in9;
 output out0;
 output out1;
 output out10;
 output out11;
 output out12;
 output out13;
 output out14;
 output out15;
 output out16;
 output out17;
 output out18;
 output out19;
 output out2;
 output out20;
 output out21;
 output out22;
 output out23;
 output out24;
 output out3;
 output out4;
 output out5;
 output out6;
 output out7;
 output out8;
 output out9;
 input rst;

 wire net0;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net63;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net64;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net65;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net66;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net67;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net68;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net69;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net7;
 wire net70;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net71;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net72;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net73;
 wire net730;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_0_net716;
 wire clknet_1_0__leaf_net716;
 wire clknet_1_1__leaf_net716;
 wire clknet_0_net64;
 wire clknet_1_0__leaf_net64;
 wire clknet_1_1__leaf_net64;
 wire clknet_0_net68;
 wire clknet_1_0__leaf_net68;
 wire clknet_1_1__leaf_net68;
 wire clknet_0_net79;
 wire clknet_1_0__leaf_net79;
 wire clknet_1_1__leaf_net79;
 wire clknet_0_net82;
 wire clknet_1_0__leaf_net82;
 wire clknet_1_1__leaf_net82;
 wire clknet_0_net84;
 wire clknet_1_0__leaf_net84;
 wire clknet_1_1__leaf_net84;
 wire clknet_0_net219;
 wire clknet_1_0__leaf_net219;
 wire clknet_1_1__leaf_net219;
 wire clknet_0_net85;
 wire clknet_1_0__leaf_net85;
 wire clknet_1_1__leaf_net85;
 wire clknet_0_net92;
 wire clknet_1_0__leaf_net92;
 wire clknet_1_1__leaf_net92;
 wire clknet_0_net102;
 wire clknet_1_0__leaf_net102;
 wire clknet_1_1__leaf_net102;
 wire clknet_0_net87;
 wire clknet_1_0__leaf_net87;
 wire clknet_1_1__leaf_net87;
 wire clknet_0_net91;
 wire clknet_1_0__leaf_net91;
 wire clknet_1_1__leaf_net91;
 wire clknet_0_net90;
 wire clknet_1_0__leaf_net90;
 wire clknet_1_1__leaf_net90;
 wire clknet_0_net89;
 wire clknet_1_0__leaf_net89;
 wire clknet_1_1__leaf_net89;
 wire clknet_0_net88;
 wire clknet_1_0__leaf_net88;
 wire clknet_1_1__leaf_net88;
 wire clknet_0_net72;
 wire clknet_1_0__leaf_net72;
 wire clknet_1_1__leaf_net72;
 wire clknet_0_net76;
 wire clknet_1_0__leaf_net76;
 wire clknet_1_1__leaf_net76;
 wire clknet_0_net78;
 wire clknet_1_0__leaf_net78;
 wire clknet_1_1__leaf_net78;
 wire clknet_0_net336;
 wire clknet_1_0__leaf_net336;
 wire clknet_1_1__leaf_net336;
 wire clknet_0_net337;
 wire clknet_1_0__leaf_net337;
 wire clknet_1_1__leaf_net337;
 wire clknet_0_net355;
 wire clknet_1_0__leaf_net355;
 wire clknet_1_1__leaf_net355;
 wire clknet_0_net361;
 wire clknet_1_0__leaf_net361;
 wire clknet_1_1__leaf_net361;
 wire clknet_0_net356;
 wire clknet_1_0__leaf_net356;
 wire clknet_1_1__leaf_net356;
 wire clknet_0_net340;
 wire clknet_1_0__leaf_net340;
 wire clknet_1_1__leaf_net340;
 wire clknet_0_net341;
 wire clknet_1_0__leaf_net341;
 wire clknet_1_1__leaf_net341;
 wire clknet_0_net215;
 wire clknet_1_0__leaf_net215;
 wire clknet_1_1__leaf_net215;
 wire clknet_0_net210;
 wire clknet_1_0__leaf_net210;
 wire clknet_1_1__leaf_net210;
 wire clknet_0_net216;
 wire clknet_1_0__leaf_net216;
 wire clknet_1_1__leaf_net216;
 wire clknet_0_net223;
 wire clknet_1_0__leaf_net223;
 wire clknet_1_1__leaf_net223;
 wire clknet_0_net218;
 wire clknet_1_0__leaf_net218;
 wire clknet_1_1__leaf_net218;
 wire clknet_0_net211;
 wire clknet_1_0__leaf_net211;
 wire clknet_1_1__leaf_net211;
 wire clknet_0_net195;
 wire clknet_1_0__leaf_net195;
 wire clknet_1_1__leaf_net195;
 wire clknet_0_net198;
 wire clknet_1_0__leaf_net198;
 wire clknet_1_1__leaf_net198;
 wire clknet_0_net202;
 wire clknet_1_0__leaf_net202;
 wire clknet_1_1__leaf_net202;
 wire clknet_0_net206;
 wire clknet_1_0__leaf_net206;
 wire clknet_1_1__leaf_net206;
 wire clknet_0_net205;
 wire clknet_1_0__leaf_net205;
 wire clknet_1_1__leaf_net205;
 wire clknet_0_net207;
 wire clknet_1_0__leaf_net207;
 wire clknet_1_1__leaf_net207;
 wire clknet_0_net200;
 wire clknet_1_0__leaf_net200;
 wire clknet_1_1__leaf_net200;
 wire clknet_0_net196;
 wire clknet_1_0__leaf_net196;
 wire clknet_1_1__leaf_net196;
 wire clknet_0_net65;
 wire clknet_1_0__leaf_net65;
 wire clknet_1_1__leaf_net65;
 wire clknet_0_net71;
 wire clknet_1_0__leaf_net71;
 wire clknet_1_1__leaf_net71;
 wire clknet_0_net77;
 wire clknet_1_0__leaf_net77;
 wire clknet_1_1__leaf_net77;
 wire clknet_0_net70;
 wire clknet_1_0__leaf_net70;
 wire clknet_1_1__leaf_net70;
 wire clknet_0_net67;
 wire clknet_1_0__leaf_net67;
 wire clknet_1_1__leaf_net67;
 wire clknet_0_net66;
 wire clknet_1_0__leaf_net66;
 wire clknet_1_1__leaf_net66;
 wire clknet_0_net69;
 wire clknet_1_0__leaf_net69;
 wire clknet_1_1__leaf_net69;
 wire clknet_0_net192;
 wire clknet_1_0__leaf_net192;
 wire clknet_1_1__leaf_net192;
 wire clknet_0_net650;
 wire clknet_1_0__leaf_net650;
 wire clknet_1_1__leaf_net650;
 wire clknet_0_net652;
 wire clknet_1_0__leaf_net652;
 wire clknet_1_1__leaf_net652;
 wire clknet_0_net680;
 wire clknet_1_0__leaf_net680;
 wire clknet_1_1__leaf_net680;
 wire clknet_0_net681;
 wire clknet_1_0__leaf_net681;
 wire clknet_1_1__leaf_net681;
 wire clknet_0_net664;
 wire clknet_1_0__leaf_net664;
 wire clknet_1_1__leaf_net664;
 wire clknet_0_net672;
 wire clknet_1_0__leaf_net672;
 wire clknet_1_1__leaf_net672;
 wire clknet_0_net673;
 wire clknet_1_0__leaf_net673;
 wire clknet_1_1__leaf_net673;
 wire clknet_0_net698;
 wire clknet_1_0__leaf_net698;
 wire clknet_1_1__leaf_net698;
 wire clknet_0_net692;
 wire clknet_1_0__leaf_net692;
 wire clknet_1_1__leaf_net692;
 wire clknet_0_net677;
 wire clknet_1_0__leaf_net677;
 wire clknet_1_1__leaf_net677;
 wire clknet_0_net659;
 wire clknet_1_0__leaf_net659;
 wire clknet_1_1__leaf_net659;
 wire clknet_0_net662;
 wire clknet_1_0__leaf_net662;
 wire clknet_1_1__leaf_net662;
 wire clknet_0_net663;
 wire clknet_1_0__leaf_net663;
 wire clknet_1_1__leaf_net663;
 wire clknet_0_net655;
 wire clknet_1_0__leaf_net655;
 wire clknet_1_1__leaf_net655;
 wire clknet_0_net654;
 wire clknet_1_0__leaf_net654;
 wire clknet_1_1__leaf_net654;
 wire clknet_0_net656;
 wire clknet_1_0__leaf_net656;
 wire clknet_1_1__leaf_net656;
 wire clknet_0_net668;
 wire clknet_1_0__leaf_net668;
 wire clknet_1_1__leaf_net668;
 wire clknet_0_net676;
 wire clknet_1_0__leaf_net676;
 wire clknet_1_1__leaf_net676;
 wire clknet_0_net653;
 wire clknet_1_0__leaf_net653;
 wire clknet_1_1__leaf_net653;
 wire clknet_0_net660;
 wire clknet_1_0__leaf_net660;
 wire clknet_1_1__leaf_net660;
 wire clknet_0_net651;
 wire clknet_1_0__leaf_net651;
 wire clknet_1_1__leaf_net651;
 wire clknet_0_net647;
 wire clknet_1_0__leaf_net647;
 wire clknet_1_1__leaf_net647;
 wire clknet_0_net648;
 wire clknet_1_0__leaf_net648;
 wire clknet_1_1__leaf_net648;
 wire clknet_0_net559;
 wire clknet_1_0__leaf_net559;
 wire clknet_1_1__leaf_net559;
 wire clknet_0_net573;
 wire clknet_1_0__leaf_net573;
 wire clknet_1_1__leaf_net573;
 wire clknet_0_net669;
 wire clknet_1_0__leaf_net669;
 wire clknet_1_1__leaf_net669;
 wire clknet_0_net581;
 wire clknet_1_0__leaf_net581;
 wire clknet_1_1__leaf_net581;
 wire clknet_0_net582;
 wire clknet_1_0__leaf_net582;
 wire clknet_1_1__leaf_net582;
 wire clknet_0_net756;
 wire clknet_1_0__leaf_net756;
 wire clknet_1_1__leaf_net756;
 wire clknet_0_net705;
 wire clknet_1_0__leaf_net705;
 wire clknet_1_1__leaf_net705;
 wire clknet_0_net757;
 wire clknet_1_0__leaf_net757;
 wire clknet_1_1__leaf_net757;
 wire clknet_0_net585;
 wire clknet_1_0__leaf_net585;
 wire clknet_1_1__leaf_net585;
 wire clknet_0_net578;
 wire clknet_1_0__leaf_net578;
 wire clknet_1_1__leaf_net578;
 wire clknet_0_net580;
 wire clknet_1_0__leaf_net580;
 wire clknet_1_1__leaf_net580;
 wire clknet_0_net584;
 wire clknet_1_0__leaf_net584;
 wire clknet_1_1__leaf_net584;
 wire clknet_0_net761;
 wire clknet_1_0__leaf_net761;
 wire clknet_1_1__leaf_net761;
 wire clknet_0_net564;
 wire clknet_1_0__leaf_net564;
 wire clknet_1_1__leaf_net564;
 wire clknet_0_net565;
 wire clknet_1_0__leaf_net565;
 wire clknet_1_1__leaf_net565;
 wire clknet_0_net558;
 wire clknet_1_0__leaf_net558;
 wire clknet_1_1__leaf_net558;
 wire clknet_0_net562;
 wire clknet_1_0__leaf_net562;
 wire clknet_1_1__leaf_net562;
 wire clknet_0_net280;
 wire clknet_1_0__leaf_net280;
 wire clknet_1_1__leaf_net280;
 wire clknet_0_net398;
 wire clknet_1_0__leaf_net398;
 wire clknet_1_1__leaf_net398;
 wire clknet_0_net404;
 wire clknet_1_0__leaf_net404;
 wire clknet_1_1__leaf_net404;
 wire clknet_0_net408;
 wire clknet_1_0__leaf_net408;
 wire clknet_1_1__leaf_net408;
 wire clknet_0_net413;
 wire clknet_1_0__leaf_net413;
 wire clknet_1_1__leaf_net413;
 wire clknet_0_net411;
 wire clknet_1_0__leaf_net411;
 wire clknet_1_1__leaf_net411;
 wire clknet_0_net409;
 wire clknet_1_0__leaf_net409;
 wire clknet_1_1__leaf_net409;
 wire clknet_0_net530;
 wire clknet_1_0__leaf_net530;
 wire clknet_1_1__leaf_net530;
 wire clknet_0_net426;
 wire clknet_1_0__leaf_net426;
 wire clknet_1_1__leaf_net426;
 wire clknet_0_net441;
 wire clknet_1_0__leaf_net441;
 wire clknet_1_1__leaf_net441;
 wire clknet_0_net410;
 wire clknet_1_0__leaf_net410;
 wire clknet_1_1__leaf_net410;
 wire clknet_0_net407;
 wire clknet_1_0__leaf_net407;
 wire clknet_1_1__leaf_net407;
 wire clknet_0_net401;
 wire clknet_1_0__leaf_net401;
 wire clknet_1_1__leaf_net401;
 wire clknet_0_net402;
 wire clknet_1_0__leaf_net402;
 wire clknet_1_1__leaf_net402;
 wire clknet_0_net406;
 wire clknet_1_0__leaf_net406;
 wire clknet_1_1__leaf_net406;
 wire clknet_0_net405;
 wire clknet_1_0__leaf_net405;
 wire clknet_1_1__leaf_net405;
 wire clknet_0_net403;
 wire clknet_1_0__leaf_net403;
 wire clknet_1_1__leaf_net403;
 wire clknet_0_net437;
 wire clknet_1_0__leaf_net437;
 wire clknet_1_1__leaf_net437;
 wire clknet_0_net439;
 wire clknet_1_0__leaf_net439;
 wire clknet_1_1__leaf_net439;
 wire clknet_0_net571;
 wire clknet_1_0__leaf_net571;
 wire clknet_1_1__leaf_net571;
 wire clknet_0_net440;
 wire clknet_1_0__leaf_net440;
 wire clknet_1_1__leaf_net440;
 wire clknet_0_net270;
 wire clknet_1_0__leaf_net270;
 wire clknet_1_1__leaf_net270;
 wire clknet_0_net272;
 wire clknet_1_0__leaf_net272;
 wire clknet_1_1__leaf_net272;
 wire clknet_0_net275;
 wire clknet_1_0__leaf_net275;
 wire clknet_1_1__leaf_net275;
 wire clknet_0_net273;
 wire clknet_1_0__leaf_net273;
 wire clknet_1_1__leaf_net273;
 wire clknet_0_net285;
 wire clknet_1_0__leaf_net285;
 wire clknet_1_1__leaf_net285;
 wire clknet_0_net300;
 wire clknet_1_0__leaf_net300;
 wire clknet_1_1__leaf_net300;
 wire clknet_0_net287;
 wire clknet_1_0__leaf_net287;
 wire clknet_1_1__leaf_net287;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;

 sky130_fd_sc_hd__a21bo_1 c100 (.A1(clknet_1_1__leaf_net76),
    .A2(net75),
    .B1_N(clknet_1_1__leaf_net79),
    .X(net80));
 sky130_fd_sc_hd__a21bo_1 c101 (.A1(clknet_1_1__leaf_net64),
    .A2(clknet_1_0__leaf_net76),
    .B1_N(clknet_1_0__leaf_net72),
    .X(net81));
 sky130_fd_sc_hd__a21bo_1 c102 (.A1(net81),
    .A2(clknet_1_0__leaf_net79),
    .B1_N(clknet_1_1__leaf_net77),
    .X(net82));
 sky130_fd_sc_hd__a31o_1 c103 (.A1(net80),
    .A2(clknet_1_1__leaf_net69),
    .A3(clknet_1_0__leaf_net82),
    .B1(clknet_1_0__leaf_net78),
    .X(net83));
 sky130_fd_sc_hd__a21bo_1 c104 (.A1(clknet_1_1__leaf_net72),
    .A2(clknet_1_1__leaf_net82),
    .B1_N(net83),
    .X(net84));
 sky130_fd_sc_hd__buf_1 c105 (.A(clknet_1_0__leaf_net84),
    .X(net85));
 sky130_fd_sc_hd__buf_1 c106 (.A(net57),
    .X(net86));
 sky130_fd_sc_hd__buf_1 c107 (.A(clknet_1_1__leaf_net85),
    .X(net87));
 sky130_fd_sc_hd__xnor2_1 c108 (.A(clknet_1_0__leaf_net87),
    .B(net86),
    .Y(net88));
 sky130_fd_sc_hd__xnor2_1 c109 (.A(clknet_1_0__leaf_net88),
    .B(clknet_1_0__leaf_net87),
    .Y(net89));
 sky130_fd_sc_hd__xnor2_1 c110 (.A(clknet_1_1__leaf_net88),
    .B(clknet_1_0__leaf_net87),
    .Y(net90));
 sky130_fd_sc_hd__xnor2_1 c111 (.A(clknet_1_1__leaf_net89),
    .B(clknet_1_0__leaf_net87),
    .Y(net91));
 sky130_fd_sc_hd__xnor2_1 c112 (.A(clknet_1_0__leaf_net85),
    .B(clknet_1_1__leaf_net87),
    .Y(net92));
 sky130_fd_sc_hd__xnor2_1 c113 (.A(net86),
    .B(clknet_1_0__leaf_net89),
    .Y(net93));
 sky130_fd_sc_hd__xnor2_1 c114 (.A(clknet_1_1__leaf_net87),
    .B(clknet_1_1__leaf_net92),
    .Y(net94));
 sky130_fd_sc_hd__sdfxbp_1 c115 (.CLK(clknet_4_5_0_clk),
    .D(clknet_1_0__leaf_net91),
    .SCD(clknet_1_0__leaf_net92),
    .SCE(clknet_1_1__leaf_net89),
    .Q(net95));
 sky130_fd_sc_hd__a21bo_1 c116 (.A1(clknet_1_0__leaf_net92),
    .A2(clknet_1_0__leaf_net90),
    .B1_N(clknet_1_0__leaf_net89),
    .X(net96));
 sky130_fd_sc_hd__dfrtp_1 c117 (.CLK(clknet_4_5_0_clk),
    .D(net96),
    .RESET_B(clknet_1_0__leaf_net84),
    .Q(net97));
 sky130_fd_sc_hd__dfsbp_1 c118 (.CLK(clknet_4_5_0_clk),
    .D(net794),
    .SET_B(clknet_1_1__leaf_net91),
    .Q(net99),
    .Q_N(net98));
 sky130_fd_sc_hd__dfsbp_1 c119 (.CLK(clknet_4_5_0_clk),
    .D(net93),
    .SET_B(clknet_1_0__leaf_net92),
    .Q(net100));
 sky130_fd_sc_hd__xnor2_1 c120 (.A(net833),
    .B(net99),
    .Y(net101));
 sky130_fd_sc_hd__a31o_1 c121 (.A1(net94),
    .A2(net101),
    .A3(net99),
    .B1(clknet_1_1__leaf_net87),
    .X(net102));
 sky130_fd_sc_hd__sdfxbp_1 c122 (.CLK(clknet_4_5_0_clk),
    .D(clknet_1_1__leaf_net90),
    .SCD(net99),
    .SCE(clknet_1_0__leaf_net102),
    .Q(net103));
 sky130_fd_sc_hd__sdfxtp_1 c123 (.CLK(clknet_4_5_0_clk),
    .D(net101),
    .SCD(clknet_1_1__leaf_net102),
    .SCE(net812),
    .Q(net104));
 sky130_fd_sc_hd__mux4_1 c124 (.A0(net100),
    .A1(net103),
    .A2(net104),
    .A3(net98),
    .S0(clknet_1_1__leaf_net92),
    .S1(clknet_1_1__leaf_net87),
    .X(net105));
 sky130_fd_sc_hd__a21bo_1 c125 (.A1(net105),
    .A2(net104),
    .B1_N(clknet_1_1__leaf_net92),
    .X(net106));
 sky130_fd_sc_hd__xnor2_1 c126 (.A(net732),
    .B(net741),
    .Y(net107));
 sky130_fd_sc_hd__xnor2_1 c127 (.A(net107),
    .B(net754),
    .Y(net108));
 sky130_fd_sc_hd__xnor2_1 c128 (.A(net108),
    .B(net736),
    .Y(net109));
 sky130_fd_sc_hd__xnor2_4 c129 (.A(net735),
    .B(net734),
    .Y(net110));
 sky130_fd_sc_hd__xnor2_1 c130 (.A(net110),
    .B(net750),
    .Y(net111));
 sky130_fd_sc_hd__xnor2_4 c131 (.A(net737),
    .B(net110),
    .Y(net112));
 sky130_fd_sc_hd__xnor2_1 c132 (.A(net111),
    .B(net743),
    .Y(net113));
 sky130_fd_sc_hd__xnor2_1 c133 (.A(net748),
    .B(net112),
    .Y(net114));
 sky130_fd_sc_hd__xnor2_1 c134 (.A(net114),
    .B(net110),
    .Y(net115));
 sky130_fd_sc_hd__xnor2_1 c135 (.A(net110),
    .B(net731),
    .Y(net116));
 sky130_fd_sc_hd__xnor2_4 c136 (.A(net112),
    .B(net740),
    .Y(net117));
 sky130_fd_sc_hd__xnor2_1 c137 (.A(net109),
    .B(net117),
    .Y(net118));
 sky130_fd_sc_hd__xnor2_2 c138 (.A(net115),
    .B(net117),
    .Y(net119));
 sky130_fd_sc_hd__xnor2_1 c139 (.A(net117),
    .B(net119),
    .Y(net120));
 sky130_fd_sc_hd__a21bo_2 c140 (.A1(net120),
    .A2(net119),
    .B1_N(net110),
    .X(net121));
 sky130_fd_sc_hd__a21bo_1 c141 (.A1(net118),
    .A2(net119),
    .B1_N(net112),
    .X(net122));
 sky130_fd_sc_hd__a21bo_1 c142 (.A1(net116),
    .A2(net117),
    .B1_N(net119),
    .X(net123));
 sky130_fd_sc_hd__a21bo_1 c143 (.A1(net119),
    .A2(net122),
    .B1_N(net123),
    .X(net124));
 sky130_fd_sc_hd__a41o_1 c144 (.A1(net113),
    .A2(net123),
    .A3(net121),
    .A4(net122),
    .B1(net110),
    .X(net125));
 sky130_fd_sc_hd__a41o_1 c145 (.A1(net124),
    .A2(net112),
    .A3(net123),
    .A4(net119),
    .B1(net110),
    .X(net126));
 sky130_fd_sc_hd__mux4_2 c146 (.A0(net125),
    .A1(net126),
    .A2(net117),
    .A3(net123),
    .S0(net110),
    .S1(net121),
    .X(net127));
 sky130_fd_sc_hd__dlymetal6s2s_1 c147 (.A(net121),
    .X(net128));
 sky130_fd_sc_hd__clkbuf_2 c148 (.A(net128),
    .X(net129));
 sky130_fd_sc_hd__clkbuf_1 c149 (.A(net129),
    .X(net130));
 sky130_fd_sc_hd__xnor2_1 c150 (.A(net16),
    .B(net128),
    .Y(net131));
 sky130_fd_sc_hd__buf_4 c151 (.A(net128),
    .X(net132));
 sky130_fd_sc_hd__xnor2_1 c152 (.A(net128),
    .B(net132),
    .Y(net133));
 sky130_fd_sc_hd__a21bo_1 c153 (.A1(net131),
    .A2(net753),
    .B1_N(net132),
    .X(net134));
 sky130_fd_sc_hd__xnor2_2 c154 (.A(net132),
    .B(net14),
    .Y(net135));
 sky130_fd_sc_hd__xnor2_4 c155 (.A(net129),
    .B(net132),
    .Y(net136));
 sky130_fd_sc_hd__xnor2_4 c156 (.A(net136),
    .B(net132),
    .Y(net137));
 sky130_fd_sc_hd__xnor2_4 c157 (.A(net2),
    .B(net136),
    .Y(net138));
 sky130_fd_sc_hd__xnor2_4 c158 (.A(net135),
    .B(net138),
    .Y(net139));
 sky130_fd_sc_hd__a21bo_1 c159 (.A1(net134),
    .A2(net139),
    .B1_N(net138),
    .X(net140));
 sky130_fd_sc_hd__xnor2_1 c160 (.A(net138),
    .B(net139),
    .Y(net141));
 sky130_fd_sc_hd__xnor2_1 c161 (.A(net140),
    .B(net141),
    .Y(net142));
 sky130_fd_sc_hd__mux4_1 c162 (.A0(net133),
    .A1(net141),
    .A2(net127),
    .A3(net138),
    .S0(net137),
    .S1(net139),
    .X(net143));
 sky130_fd_sc_hd__a21bo_1 c163 (.A1(net129),
    .A2(net138),
    .B1_N(net137),
    .X(net144));
 sky130_fd_sc_hd__xnor2_1 c164 (.A(net142),
    .B(net143),
    .Y(net145));
 sky130_fd_sc_hd__dfstp_1 c165 (.CLK(clknet_4_0_0_clk),
    .D(net141),
    .SET_B(net145),
    .Q(net146));
 sky130_fd_sc_hd__xnor2_1 c166 (.A(net130),
    .B(net146),
    .Y(net147));
 sky130_fd_sc_hd__xnor2_2 c167 (.A(net147),
    .B(net139),
    .Y(net148));
 sky130_fd_sc_hd__buf_1 c168 (.A(net26),
    .X(net149));
 sky130_fd_sc_hd__buf_1 c169 (.A(net149),
    .X(net150));
 sky130_fd_sc_hd__xnor2_1 c170 (.A(net149),
    .B(net150),
    .Y(net151));
 sky130_fd_sc_hd__clkbuf_2 c171 (.A(net150),
    .X(net152));
 sky130_fd_sc_hd__buf_2 c172 (.A(net149),
    .X(net153));
 sky130_fd_sc_hd__clkbuf_2 c173 (.A(net149),
    .X(net154));
 sky130_fd_sc_hd__xnor2_4 c174 (.A(net152),
    .B(net153),
    .Y(net155));
 sky130_fd_sc_hd__xnor2_1 c175 (.A(net154),
    .B(net155),
    .Y(net156));
 sky130_fd_sc_hd__a21bo_1 c176 (.A1(net150),
    .A2(net156),
    .B1_N(net154),
    .X(net157));
 sky130_fd_sc_hd__xnor2_2 c177 (.A(net154),
    .B(net155),
    .Y(net158));
 sky130_fd_sc_hd__a31o_1 c178 (.A1(net150),
    .A2(net158),
    .A3(net155),
    .B1(net156),
    .X(net159));
 sky130_fd_sc_hd__a31o_2 c179 (.A1(net156),
    .A2(net154),
    .A3(net773),
    .B1(net158),
    .X(net160));
 sky130_fd_sc_hd__xnor2_1 c180 (.A(net153),
    .B(net160),
    .Y(net161));
 sky130_fd_sc_hd__a21bo_1 c181 (.A1(net157),
    .A2(net158),
    .B1_N(net154),
    .X(net162));
 sky130_fd_sc_hd__a21bo_1 c182 (.A1(net155),
    .A2(net158),
    .B1_N(net160),
    .X(net163));
 sky130_fd_sc_hd__dfstp_1 c183 (.CLK(clknet_4_1_0_clk),
    .D(net159),
    .SET_B(net163),
    .Q(net164));
 sky130_fd_sc_hd__sdfxtp_1 c184 (.CLK(clknet_4_4_0_clk),
    .D(net151),
    .SCD(net152),
    .SCE(net162),
    .Q(net165));
 sky130_fd_sc_hd__dfstp_1 c185 (.CLK(clknet_4_4_0_clk),
    .D(net161),
    .SET_B(net787),
    .Q(net166));
 sky130_fd_sc_hd__sdfrbp_1 c186 (.CLK(clknet_4_4_0_clk),
    .D(net158),
    .RESET_B(net163),
    .SCD(net166),
    .SCE(net152),
    .Q(net167));
 sky130_fd_sc_hd__a21bo_1 c187 (.A1(net167),
    .A2(net153),
    .B1_N(net165),
    .X(net168));
 sky130_fd_sc_hd__mux4_1 c188 (.A0(net166),
    .A1(net168),
    .A2(net163),
    .A3(net165),
    .S0(net158),
    .S1(net160),
    .X(net169));
 sky130_fd_sc_hd__dlrbn_2 c189 (.D(net162),
    .GATE_N(clknet_4_4_0_clk),
    .RESET_B(net160),
    .Q(net171),
    .Q_N(net170));
 sky130_fd_sc_hd__xnor2_1 c190 (.A(net171),
    .B(net42),
    .Y(net172));
 sky130_fd_sc_hd__dlrbn_2 c191 (.D(net171),
    .GATE_N(clknet_4_4_0_clk),
    .RESET_B(net172),
    .Q(net174),
    .Q_N(net173));
 sky130_fd_sc_hd__dlrbp_1 c192 (.D(net172),
    .GATE(clknet_4_4_0_clk),
    .RESET_B(net174),
    .Q(net176),
    .Q_N(net175));
 sky130_fd_sc_hd__dlrbp_2 c193 (.D(net171),
    .GATE(clknet_4_5_0_clk),
    .RESET_B(net172),
    .Q(net178),
    .Q_N(net177));
 sky130_fd_sc_hd__xnor2_4 c194 (.A(net175),
    .B(net170),
    .Y(net179));
 sky130_fd_sc_hd__xnor2_4 c195 (.A(net179),
    .B(net178),
    .Y(net180));
 sky130_fd_sc_hd__xnor2_4 c196 (.A(net179),
    .B(net178),
    .Y(net181));
 sky130_fd_sc_hd__xnor2_4 c197 (.A(net180),
    .B(net181),
    .Y(net182));
 sky130_fd_sc_hd__a21bo_4 c198 (.A1(net178),
    .A2(net179),
    .B1_N(net182),
    .X(net183));
 sky130_fd_sc_hd__xnor2_1 c199 (.A(net182),
    .B(net173),
    .Y(net184));
 sky130_fd_sc_hd__xnor2_4 c200 (.A(net782),
    .B(net183),
    .Y(net185));
 sky130_fd_sc_hd__xnor2_4 c201 (.A(net174),
    .B(net178),
    .Y(net186));
 sky130_fd_sc_hd__a41o_4 c202 (.A1(net185),
    .A2(net183),
    .A3(net186),
    .A4(net170),
    .B1(net182),
    .X(net187));
 sky130_fd_sc_hd__xnor2_4 c203 (.A(net186),
    .B(net780),
    .Y(net188));
 sky130_fd_sc_hd__a31o_1 c204 (.A1(net187),
    .A2(net182),
    .A3(net177),
    .B1(clknet_1_1__leaf_net716),
    .X(net189));
 sky130_fd_sc_hd__a21bo_1 c205 (.A1(net187),
    .A2(net776),
    .B1_N(net177),
    .X(net190));
 sky130_fd_sc_hd__a41o_1 c206 (.A1(net176),
    .A2(net186),
    .A3(net776),
    .A4(net173),
    .B1(net177),
    .X(net191));
 sky130_fd_sc_hd__a31o_1 c207 (.A1(net189),
    .A2(net185),
    .A3(net191),
    .B1(net776),
    .X(net192));
 sky130_fd_sc_hd__a41o_1 c208 (.A1(net190),
    .A2(net191),
    .A3(clknet_1_0__leaf_net192),
    .A4(net186),
    .B1(net781),
    .X(net193));
 sky130_fd_sc_hd__a31o_1 c209 (.A1(net183),
    .A2(net193),
    .A3(net174),
    .B1(net188),
    .X(net194));
 sky130_fd_sc_hd__xnor2_1 c210 (.A(clknet_1_0__leaf_net78),
    .B(clknet_1_0__leaf_net70),
    .Y(net195));
 sky130_fd_sc_hd__xnor2_4 c211 (.A(clknet_1_0__leaf_net195),
    .B(clknet_1_1__leaf_net192),
    .Y(net196));
 sky130_fd_sc_hd__buf_1 c212 (.A(clknet_1_0__leaf_net196),
    .X(net197));
 sky130_fd_sc_hd__xnor2_4 c213 (.A(clknet_1_0__leaf_net196),
    .B(clknet_1_0__leaf_net195),
    .Y(net198));
 sky130_fd_sc_hd__xnor2_1 c214 (.A(net197),
    .B(clknet_1_1__leaf_net198),
    .Y(net199));
 sky130_fd_sc_hd__xnor2_4 c215 (.A(net785),
    .B(clknet_1_0__leaf_net198),
    .Y(net200));
 sky130_fd_sc_hd__xnor2_1 c216 (.A(clknet_1_1__leaf_net196),
    .B(clknet_1_0__leaf_net200),
    .Y(net201));
 sky130_fd_sc_hd__xnor2_1 c217 (.A(net199),
    .B(clknet_1_0__leaf_net198),
    .Y(net202));
 sky130_fd_sc_hd__xnor2_1 c218 (.A(clknet_1_0__leaf_net78),
    .B(clknet_1_1__leaf_net195),
    .Y(net203));
 sky130_fd_sc_hd__xnor2_4 c219 (.A(net188),
    .B(clknet_1_0__leaf_net200),
    .Y(net204));
 sky130_fd_sc_hd__xnor2_1 c220 (.A(clknet_1_0__leaf_net202),
    .B(clknet_1_1__leaf_net196),
    .Y(net205));
 sky130_fd_sc_hd__xnor2_1 c221 (.A(net201),
    .B(clknet_1_0__leaf_net202),
    .Y(net206));
 sky130_fd_sc_hd__xnor2_1 c222 (.A(clknet_1_1__leaf_net70),
    .B(clknet_1_1__leaf_net205),
    .Y(net207));
 sky130_fd_sc_hd__xnor2_1 c223 (.A(clknet_1_0__leaf_net205),
    .B(clknet_1_0__leaf_net207),
    .Y(net208));
 sky130_fd_sc_hd__sdfxtp_1 c224 (.CLK(clknet_4_6_0_clk),
    .D(net208),
    .SCD(clknet_1_0__leaf_net205),
    .SCE(clknet_1_1__leaf_net195),
    .Q(net209));
 sky130_fd_sc_hd__xnor2_4 c225 (.A(net203),
    .B(net204),
    .Y(net210));
 sky130_fd_sc_hd__a21bo_1 c226 (.A1(clknet_1_0__leaf_net206),
    .A2(net209),
    .B1_N(clknet_1_0__leaf_net210),
    .X(net211));
 sky130_fd_sc_hd__a21bo_1 c227 (.A1(clknet_1_0__leaf_net211),
    .A2(clknet_1_0__leaf_net210),
    .B1_N(clknet_1_1__leaf_net206),
    .X(net212));
 sky130_fd_sc_hd__dfbbn_1 c228 (.CLK_N(clknet_4_7_0_clk),
    .D(clknet_1_1__leaf_net200),
    .RESET_B(net212),
    .SET_B(clknet_1_0__leaf_net210),
    .Q(net213));
 sky130_fd_sc_hd__mux4_1 c229 (.A0(net184),
    .A1(net213),
    .A2(clknet_1_0__leaf_net206),
    .A3(clknet_1_1__leaf_net202),
    .S0(clknet_1_1__leaf_net78),
    .S1(clknet_1_1__leaf_net205),
    .X(net214));
 sky130_fd_sc_hd__a21bo_1 c230 (.A1(net214),
    .A2(clknet_1_1__leaf_net211),
    .B1_N(clknet_1_1__leaf_net196),
    .X(net215));
 sky130_fd_sc_hd__buf_6 c231 (.A(clknet_1_0__leaf_net210),
    .X(net216));
 sky130_fd_sc_hd__dfxbp_1 c232 (.CLK(clknet_4_7_0_clk),
    .D(net106),
    .Q(net217));
 sky130_fd_sc_hd__buf_1 c233 (.A(clknet_1_1__leaf_net216),
    .X(net769));
 sky130_fd_sc_hd__xnor2_1 c234 (.A(net194),
    .B(clknet_1_0__leaf_net216),
    .Y(net218));
 sky130_fd_sc_hd__xnor2_1 c235 (.A(clknet_1_0__leaf_net216),
    .B(clknet_1_1__leaf_net84),
    .Y(net219));
 sky130_fd_sc_hd__dlrtn_1 c236 (.D(clknet_1_0__leaf_net218),
    .GATE_N(clknet_4_7_0_clk),
    .RESET_B(clknet_1_0__leaf_net219),
    .Q(net220));
 sky130_fd_sc_hd__dlrtn_1 c237 (.D(net220),
    .GATE_N(clknet_4_7_0_clk),
    .RESET_B(clknet_1_0__leaf_net219),
    .Q(net221));
 sky130_fd_sc_hd__dlrtn_1 c238 (.D(clknet_1_0__leaf_net218),
    .GATE_N(clknet_4_7_0_clk),
    .RESET_B(clknet_1_0__leaf_net219),
    .Q(net222));
 sky130_fd_sc_hd__xnor2_4 c239 (.A(net221),
    .B(clknet_1_1__leaf_net216),
    .Y(net223));
 sky130_fd_sc_hd__dlrtp_1 c240 (.D(net222),
    .GATE(clknet_4_7_0_clk),
    .RESET_B(clknet_1_1__leaf_net223),
    .Q(net224));
 sky130_fd_sc_hd__dfbbn_1 c241 (.CLK_N(clknet_4_7_0_clk),
    .D(net217),
    .RESET_B(clknet_1_0__leaf_net223),
    .SET_B(clknet_1_0__leaf_net218),
    .Q(net226),
    .Q_N(net225));
 sky130_fd_sc_hd__sdfbbn_1 c242 (.CLK_N(clknet_4_7_0_clk),
    .D(clknet_1_1__leaf_net219),
    .RESET_B(net226),
    .SCD(net222),
    .SCE(clknet_1_0__leaf_net223),
    .SET_B(clknet_1_1__leaf_net218),
    .Q(net227));
 sky130_fd_sc_hd__xnor2_1 c243 (.A(net224),
    .B(net222),
    .Y(net228));
 sky130_fd_sc_hd__xnor2_1 c244 (.A(net227),
    .B(net222),
    .Y(net229));
 sky130_fd_sc_hd__a21bo_1 c245 (.A1(net228),
    .A2(net226),
    .B1_N(net222),
    .X(net230));
 sky130_fd_sc_hd__dfbbp_1 c246 (.CLK(clknet_4_7_0_clk),
    .D(net229),
    .RESET_B(clknet_1_1__leaf_net218),
    .SET_B(net225),
    .Q(net231));
 sky130_fd_sc_hd__dlrtp_1 c247 (.D(net231),
    .GATE(clknet_4_7_0_clk),
    .RESET_B(clknet_1_1__leaf_net215),
    .Q(net232));
 sky130_fd_sc_hd__sdfxbp_1 c248 (.CLK(clknet_4_7_0_clk),
    .D(net226),
    .SCD(clknet_1_1__leaf_net218),
    .SCE(net222),
    .Q(net234),
    .Q_N(net233));
 sky130_fd_sc_hd__sdfxbp_1 c249 (.CLK(clknet_4_7_0_clk),
    .D(net797),
    .SCD(clknet_1_1__leaf_net219),
    .SCE(net821),
    .Q(net235));
 sky130_fd_sc_hd__xnor2_1 c25 (.A(net739),
    .B(net745),
    .Y(net0));
 sky130_fd_sc_hd__dlrtp_1 c250 (.D(clknet_1_1__leaf_net223),
    .GATE(clknet_4_7_0_clk),
    .RESET_B(net234),
    .Q(net236));
 sky130_fd_sc_hd__a21bo_1 c251 (.A1(net236),
    .A2(net234),
    .B1_N(net225),
    .X(net237));
 sky130_fd_sc_hd__buf_4 c252 (.A(net121),
    .X(net238));
 sky130_fd_sc_hd__xnor2_4 c253 (.A(net238),
    .B(net121),
    .Y(net239));
 sky130_fd_sc_hd__xnor2_4 c254 (.A(net239),
    .B(net127),
    .Y(net240));
 sky130_fd_sc_hd__xnor2_2 c255 (.A(net239),
    .B(net238),
    .Y(net241));
 sky130_fd_sc_hd__xnor2_2 c256 (.A(net238),
    .B(net241),
    .Y(net242));
 sky130_fd_sc_hd__xnor2_4 c257 (.A(net775),
    .B(net240),
    .Y(net243));
 sky130_fd_sc_hd__xnor2_4 c258 (.A(net243),
    .B(net775),
    .Y(net244));
 sky130_fd_sc_hd__xnor2_4 c259 (.A(net244),
    .B(net238),
    .Y(net245));
 sky130_fd_sc_hd__xnor2_1 c26 (.A(net744),
    .B(net745),
    .Y(net1));
 sky130_fd_sc_hd__xnor2_2 c260 (.A(net240),
    .B(net245),
    .Y(net246));
 sky130_fd_sc_hd__xnor2_4 c261 (.A(net245),
    .B(net246),
    .Y(net247));
 sky130_fd_sc_hd__xnor2_1 c262 (.A(net244),
    .B(net240),
    .Y(net248));
 sky130_fd_sc_hd__edfxbp_1 c263 (.CLK(clknet_4_0_0_clk),
    .D(net246),
    .DE(net247),
    .Q(net250),
    .Q_N(net249));
 sky130_fd_sc_hd__a31o_1 c264 (.A1(net241),
    .A2(net250),
    .A3(net242),
    .B1(net239),
    .X(net251));
 sky130_fd_sc_hd__a21bo_1 c265 (.A1(net121),
    .A2(net251),
    .B1_N(net241),
    .X(net252));
 sky130_fd_sc_hd__a31o_1 c266 (.A1(net242),
    .A2(net248),
    .A3(net245),
    .B1(net775),
    .X(net253));
 sky130_fd_sc_hd__xnor2_1 c267 (.A(net243),
    .B(net248),
    .Y(net254));
 sky130_fd_sc_hd__a31o_1 c268 (.A1(net245),
    .A2(net252),
    .A3(net249),
    .B1(net242),
    .X(net255));
 sky130_fd_sc_hd__a21bo_1 c269 (.A1(net254),
    .A2(net255),
    .B1_N(net243),
    .X(net256));
 sky130_fd_sc_hd__a21bo_2 c27 (.A1(net746),
    .A2(net749),
    .B1_N(net744),
    .X(net2));
 sky130_fd_sc_hd__sdfbbn_1 c270 (.CLK_N(clknet_4_0_0_clk),
    .D(net252),
    .RESET_B(net256),
    .SCD(net242),
    .SCE(net775),
    .SET_B(net247),
    .Q(net258),
    .Q_N(net257));
 sky130_fd_sc_hd__mux4_1 c271 (.A0(net253),
    .A1(net251),
    .A2(net254),
    .A3(net257),
    .S0(net775),
    .S1(net256),
    .X(net259));
 sky130_fd_sc_hd__a21bo_1 c272 (.A1(net258),
    .A2(net255),
    .B1_N(net718),
    .X(net260));
 sky130_fd_sc_hd__edfxtp_1 c273 (.CLK(clknet_4_0_0_clk),
    .D(net260),
    .DE(net773),
    .Q(net261));
 sky130_fd_sc_hd__xnor2_4 c274 (.A(net148),
    .B(net137),
    .Y(net262));
 sky130_fd_sc_hd__xnor2_1 c275 (.A(net261),
    .B(net262),
    .Y(net263));
 sky130_fd_sc_hd__sdlclkp_1 c276 (.CLK(clknet_4_0_0_clk),
    .GATE(net263),
    .SCE(net261),
    .GCLK(net264));
 sky130_fd_sc_hd__xnor2_1 c277 (.A(net773),
    .B(net261),
    .Y(net265));
 sky130_fd_sc_hd__xnor2_2 c278 (.A(net127),
    .B(net249),
    .Y(net266));
 sky130_fd_sc_hd__a21bo_1 c279 (.A1(net264),
    .A2(net261),
    .B1_N(net262),
    .X(net267));
 sky130_fd_sc_hd__xnor2_1 c28 (.A(net1),
    .B(net745),
    .Y(net3));
 sky130_fd_sc_hd__xnor2_1 c280 (.A(net144),
    .B(net261),
    .Y(net268));
 sky130_fd_sc_hd__xnor2_1 c281 (.A(net268),
    .B(net773),
    .Y(net269));
 sky130_fd_sc_hd__sdlclkp_2 c282 (.CLK(clknet_4_0_0_clk),
    .GATE(net269),
    .SCE(net263),
    .GCLK(net270));
 sky130_fd_sc_hd__xnor2_1 c283 (.A(net261),
    .B(net266),
    .Y(net271));
 sky130_fd_sc_hd__xnor2_1 c284 (.A(net266),
    .B(clknet_1_0__leaf_net270),
    .Y(net272));
 sky130_fd_sc_hd__a21bo_1 c285 (.A1(net265),
    .A2(net266),
    .B1_N(clknet_1_1__leaf_net272),
    .X(net273));
 sky130_fd_sc_hd__a21bo_1 c286 (.A1(clknet_1_1__leaf_net270),
    .A2(clknet_1_1__leaf_net272),
    .B1_N(net262),
    .X(net274));
 sky130_fd_sc_hd__xnor2_1 c287 (.A(clknet_1_0__leaf_net272),
    .B(net262),
    .Y(net275));
 sky130_fd_sc_hd__sdfrbp_1 c288 (.CLK(clknet_4_0_0_clk),
    .D(net274),
    .RESET_B(clknet_1_1__leaf_net272),
    .SCD(clknet_1_0__leaf_net273),
    .SCE(net265),
    .Q(net277),
    .Q_N(net276));
 sky130_fd_sc_hd__sdfxtp_1 c289 (.CLK(clknet_4_1_0_clk),
    .D(clknet_1_0__leaf_net275),
    .SCD(clknet_1_0__leaf_net270),
    .SCE(clknet_1_0__leaf_net272),
    .Q(net278));
 sky130_fd_sc_hd__xnor2_1 c29 (.A(net745),
    .B(net744),
    .Y(net4));
 sky130_fd_sc_hd__sdfbbp_1 c290 (.CLK(clknet_4_1_0_clk),
    .D(net271),
    .RESET_B(clknet_1_0__leaf_net275),
    .SCD(net818),
    .SCE(clknet_1_0__leaf_net272),
    .SET_B(net262),
    .Q(net279));
 sky130_fd_sc_hd__sdlclkp_4 c291 (.CLK(clknet_4_1_0_clk),
    .GATE(net262),
    .SCE(clknet_1_1__leaf_net275),
    .GCLK(net280));
 sky130_fd_sc_hd__mux4_1 c292 (.A0(clknet_1_1__leaf_net280),
    .A1(net271),
    .A2(net276),
    .A3(clknet_1_1__leaf_net270),
    .S0(net278),
    .S1(clknet_1_1__leaf_net275),
    .X(net281));
 sky130_fd_sc_hd__a31o_1 c293 (.A1(net279),
    .A2(net818),
    .A3(clknet_1_1__leaf_net270),
    .B1(clknet_1_0__leaf_net280),
    .X(net282));
 sky130_fd_sc_hd__buf_1 c294 (.A(net160),
    .X(net283));
 sky130_fd_sc_hd__buf_1 c295 (.A(net717),
    .X(net284));
 sky130_fd_sc_hd__xnor2_1 c296 (.A(clknet_1_1__leaf_net273),
    .B(net284),
    .Y(net285));
 sky130_fd_sc_hd__clkbuf_2 c297 (.A(net720),
    .X(net286));
 sky130_fd_sc_hd__xnor2_1 c298 (.A(clknet_1_0__leaf_net285),
    .B(net286),
    .Y(net287));
 sky130_fd_sc_hd__dfrbp_2 c299 (.CLK(clknet_4_3_0_clk),
    .D(net283),
    .RESET_B(net786),
    .Q(net289),
    .Q_N(net288));
 sky130_fd_sc_hd__xnor2_1 c30 (.A(net747),
    .B(net744),
    .Y(net5));
 sky130_fd_sc_hd__xnor2_2 c300 (.A(net286),
    .B(net289),
    .Y(net290));
 sky130_fd_sc_hd__xnor2_1 c301 (.A(net290),
    .B(net286),
    .Y(net291));
 sky130_fd_sc_hd__dfrbp_1 c302 (.CLK(clknet_4_1_0_clk),
    .D(net284),
    .RESET_B(net283),
    .Q(net292));
 sky130_fd_sc_hd__dfrtn_1 c303 (.CLK_N(clknet_4_1_0_clk),
    .D(net292),
    .RESET_B(clknet_1_0__leaf_net287),
    .Q(net293));
 sky130_fd_sc_hd__xnor2_1 c304 (.A(net291),
    .B(net293),
    .Y(net294));
 sky130_fd_sc_hd__dfrtp_1 c305 (.CLK(clknet_4_4_0_clk),
    .D(clknet_1_1__leaf_net287),
    .RESET_B(net160),
    .Q(net295));
 sky130_fd_sc_hd__xnor2_1 c306 (.A(net295),
    .B(net289),
    .Y(net296));
 sky130_fd_sc_hd__xnor2_1 c307 (.A(net164),
    .B(net294),
    .Y(net297));
 sky130_fd_sc_hd__xnor2_1 c308 (.A(net293),
    .B(net296),
    .Y(net298));
 sky130_fd_sc_hd__xnor2_1 c309 (.A(net298),
    .B(net788),
    .Y(net299));
 sky130_fd_sc_hd__xnor2_2 c31 (.A(net8),
    .B(net744),
    .Y(net6));
 sky130_fd_sc_hd__xnor2_1 c310 (.A(clknet_1_0__leaf_net285),
    .B(net290),
    .Y(net300));
 sky130_fd_sc_hd__dfrtp_1 c311 (.CLK(clknet_4_6_0_clk),
    .D(clknet_1_0__leaf_net300),
    .RESET_B(net789),
    .Q(net301));
 sky130_fd_sc_hd__a41o_1 c312 (.A1(net291),
    .A2(net298),
    .A3(net296),
    .A4(net290),
    .B1(clknet_1_1__leaf_net285),
    .X(net302));
 sky130_fd_sc_hd__sdfxtp_2 c313 (.CLK(clknet_4_6_0_clk),
    .D(net799),
    .SCD(clknet_1_1__leaf_net300),
    .SCE(net299),
    .Q(net303));
 sky130_fd_sc_hd__sdfxtp_1 c314 (.CLK(clknet_4_3_0_clk),
    .D(net302),
    .SCD(net297),
    .SCE(net294),
    .Q(net304));
 sky130_fd_sc_hd__xnor2_4 c315 (.A(net790),
    .B(net188),
    .Y(net305));
 sky130_fd_sc_hd__xnor2_4 c316 (.A(net305),
    .B(net777),
    .Y(net306));
 sky130_fd_sc_hd__xnor2_4 c317 (.A(net42),
    .B(net188),
    .Y(net307));
 sky130_fd_sc_hd__xnor2_1 c318 (.A(net305),
    .B(net306),
    .Y(net308));
 sky130_fd_sc_hd__dfrtp_4 c319 (.CLK(clknet_4_6_0_clk),
    .D(net307),
    .RESET_B(net305),
    .Q(net309));
 sky130_fd_sc_hd__xnor2_1 c32 (.A(net3),
    .B(net6),
    .Y(net7));
 sky130_fd_sc_hd__xnor2_4 c320 (.A(net309),
    .B(net306),
    .Y(net310));
 sky130_fd_sc_hd__dfbbn_1 c321 (.CLK_N(clknet_4_6_0_clk),
    .D(net305),
    .RESET_B(net307),
    .SET_B(net310),
    .Q(net312),
    .Q_N(net311));
 sky130_fd_sc_hd__a21bo_1 c322 (.A1(net310),
    .A2(net306),
    .B1_N(net309),
    .X(net313));
 sky130_fd_sc_hd__dfsbp_1 c323 (.CLK(clknet_4_6_0_clk),
    .D(net790),
    .SET_B(net307),
    .Q(net314));
 sky130_fd_sc_hd__a21bo_1 c324 (.A1(net306),
    .A2(net310),
    .B1_N(net313),
    .X(net315));
 sky130_fd_sc_hd__a21bo_1 c325 (.A1(net308),
    .A2(net306),
    .B1_N(net311),
    .X(net316));
 sky130_fd_sc_hd__xnor2_1 c326 (.A(net309),
    .B(net312),
    .Y(net317));
 sky130_fd_sc_hd__dfbbn_1 c327 (.CLK_N(clknet_4_6_0_clk),
    .D(net307),
    .RESET_B(net316),
    .SET_B(net310),
    .Q(net319),
    .Q_N(net318));
 sky130_fd_sc_hd__xnor2_1 c328 (.A(net316),
    .B(net313),
    .Y(net320));
 sky130_fd_sc_hd__dfbbp_1 c329 (.CLK(clknet_4_6_0_clk),
    .D(net317),
    .RESET_B(net316),
    .SET_B(net307),
    .Q(net322),
    .Q_N(net321));
 sky130_fd_sc_hd__a21bo_1 c33 (.A1(net751),
    .A2(net752),
    .B1_N(net742),
    .X(net8));
 sky130_fd_sc_hd__a21bo_1 c330 (.A1(net320),
    .A2(net310),
    .B1_N(net321),
    .X(net323));
 sky130_fd_sc_hd__a21bo_1 c331 (.A1(net778),
    .A2(net323),
    .B1_N(net316),
    .X(net324));
 sky130_fd_sc_hd__mux4_1 c332 (.A0(net313),
    .A1(net322),
    .A2(net324),
    .A3(net316),
    .S0(net310),
    .S1(net288),
    .X(net325));
 sky130_fd_sc_hd__mux4_1 c333 (.A0(net319),
    .A1(net325),
    .A2(net320),
    .A3(net307),
    .S0(net779),
    .S1(net306),
    .X(net326));
 sky130_fd_sc_hd__mux4_1 c334 (.A0(net315),
    .A1(net320),
    .A2(net318),
    .A3(net316),
    .S0(net307),
    .S1(net721),
    .X(net327));
 sky130_fd_sc_hd__mux4_1 c335 (.A0(net324),
    .A1(net322),
    .A2(net306),
    .A3(net313),
    .S0(net721),
    .S1(net722),
    .X(net328));
 sky130_fd_sc_hd__dfsbp_2 c336 (.CLK(clknet_4_6_0_clk),
    .D(clknet_1_1__leaf_net207),
    .SET_B(clknet_1_0__leaf_net215),
    .Q(net330),
    .Q_N(net329));
 sky130_fd_sc_hd__buf_4 c337 (.A(net330),
    .X(net331));
 sky130_fd_sc_hd__xnor2_4 c338 (.A(net331),
    .B(net330),
    .Y(net332));
 sky130_fd_sc_hd__xnor2_4 c339 (.A(net332),
    .B(net331),
    .Y(net333));
 sky130_fd_sc_hd__xnor2_1 c34 (.A(net4),
    .B(net6),
    .Y(net9));
 sky130_fd_sc_hd__sdfxbp_1 c340 (.CLK(clknet_4_7_0_clk),
    .D(net333),
    .SCD(clknet_1_0__leaf_net215),
    .SCE(net332),
    .Q(net334));
 sky130_fd_sc_hd__xnor2_2 c341 (.A(net333),
    .B(net311),
    .Y(net335));
 sky130_fd_sc_hd__xnor2_1 c342 (.A(net333),
    .B(clknet_1_1__leaf_net78),
    .Y(net336));
 sky130_fd_sc_hd__xnor2_1 c343 (.A(clknet_1_0__leaf_net336),
    .B(net329),
    .Y(net337));
 sky130_fd_sc_hd__xnor2_1 c344 (.A(net335),
    .B(net329),
    .Y(net338));
 sky130_fd_sc_hd__xnor2_1 c345 (.A(net330),
    .B(net332),
    .Y(net339));
 sky130_fd_sc_hd__xnor2_1 c346 (.A(net339),
    .B(clknet_1_0__leaf_net337),
    .Y(net340));
 sky130_fd_sc_hd__xnor2_1 c347 (.A(net332),
    .B(clknet_1_0__leaf_net340),
    .Y(net341));
 sky130_fd_sc_hd__a31o_1 c348 (.A1(net335),
    .A2(clknet_1_0__leaf_net341),
    .A3(net332),
    .B1(net333),
    .X(net342));
 sky130_fd_sc_hd__a21bo_1 c349 (.A1(clknet_1_1__leaf_net336),
    .A2(clknet_1_0__leaf_net340),
    .B1_N(net339),
    .X(net343));
 sky130_fd_sc_hd__a21bo_1 c35 (.A1(net5),
    .A2(net744),
    .B1_N(net7),
    .X(net10));
 sky130_fd_sc_hd__a21bo_1 c350 (.A1(net342),
    .A2(clknet_1_0__leaf_net341),
    .B1_N(clknet_1_0__leaf_net336),
    .X(net344));
 sky130_fd_sc_hd__xnor2_1 c351 (.A(net334),
    .B(clknet_1_1__leaf_net341),
    .Y(net345));
 sky130_fd_sc_hd__xnor2_1 c352 (.A(clknet_1_1__leaf_net337),
    .B(net331),
    .Y(net346));
 sky130_fd_sc_hd__xnor2_1 c353 (.A(net338),
    .B(clknet_1_0__leaf_net341),
    .Y(net347));
 sky130_fd_sc_hd__xnor2_1 c354 (.A(net346),
    .B(clknet_1_1__leaf_net340),
    .Y(net348));
 sky130_fd_sc_hd__xnor2_1 c355 (.A(net344),
    .B(net335),
    .Y(net349));
 sky130_fd_sc_hd__a21bo_1 c356 (.A1(net349),
    .A2(clknet_1_0__leaf_net341),
    .B1_N(net333),
    .X(net350));
 sky130_fd_sc_hd__buf_2 c357 (.A(net235),
    .X(net351));
 sky130_fd_sc_hd__dfstp_1 c358 (.CLK(clknet_4_7_0_clk),
    .D(clknet_1_1__leaf_net219),
    .SET_B(clknet_1_1__leaf_net215),
    .Q(net352));
 sky130_fd_sc_hd__xnor2_4 c359 (.A(net237),
    .B(net351),
    .Y(net353));
 sky130_fd_sc_hd__a21bo_1 c36 (.A1(net9),
    .A2(net10),
    .B1_N(net745),
    .X(net11));
 sky130_fd_sc_hd__xnor2_1 c360 (.A(net351),
    .B(net331),
    .Y(net354));
 sky130_fd_sc_hd__a31o_1 c361 (.A1(net348),
    .A2(net353),
    .A3(clknet_1_1__leaf_net210),
    .B1(net351),
    .X(net355));
 sky130_fd_sc_hd__a21bo_1 c362 (.A1(net354),
    .A2(clknet_1_0__leaf_net355),
    .B1_N(net351),
    .X(net356));
 sky130_fd_sc_hd__dfstp_1 c363 (.CLK(clknet_4_13_0_clk),
    .D(clknet_1_0__leaf_net355),
    .SET_B(clknet_1_0__leaf_net356),
    .Q(net357));
 sky130_fd_sc_hd__xnor2_2 c364 (.A(net828),
    .B(net353),
    .Y(net358));
 sky130_fd_sc_hd__sdfxbp_1 c365 (.CLK(clknet_4_13_0_clk),
    .D(net345),
    .SCD(net358),
    .SCE(clknet_1_0__leaf_net356),
    .Q(net360),
    .Q_N(net359));
 sky130_fd_sc_hd__a21bo_1 c366 (.A1(net353),
    .A2(clknet_1_1__leaf_net355),
    .B1_N(net359),
    .X(net361));
 sky130_fd_sc_hd__dfstp_1 c367 (.CLK(clknet_4_13_0_clk),
    .D(net343),
    .SET_B(clknet_1_0__leaf_net361),
    .Q(net362));
 sky130_fd_sc_hd__sdfxtp_1 c368 (.CLK(clknet_4_13_0_clk),
    .D(net230),
    .SCD(clknet_1_0__leaf_net356),
    .SCE(net809),
    .Q(net363));
 sky130_fd_sc_hd__dlrbn_1 c369 (.D(net822),
    .GATE_N(clknet_4_13_0_clk),
    .RESET_B(clknet_1_1__leaf_net356),
    .Q(net365),
    .Q_N(net364));
 sky130_fd_sc_hd__xnor2_1 c37 (.A(net11),
    .B(net10),
    .Y(net12));
 sky130_fd_sc_hd__dlrbn_1 c370 (.D(clknet_1_1__leaf_net361),
    .GATE_N(clknet_4_13_0_clk),
    .RESET_B(net358),
    .Q(net367),
    .Q_N(net366));
 sky130_fd_sc_hd__sdfrtn_1 c371 (.CLK_N(clknet_4_13_0_clk),
    .D(net801),
    .RESET_B(clknet_1_1__leaf_net356),
    .SCD(net358),
    .SCE(net353),
    .Q(net368));
 sky130_fd_sc_hd__sdfrtp_1 c372 (.CLK(clknet_4_13_0_clk),
    .D(net809),
    .RESET_B(net368),
    .SCD(net358),
    .SCE(clknet_1_1__leaf_net356),
    .Q(net369));
 sky130_fd_sc_hd__mux4_1 c373 (.A0(net367),
    .A1(net353),
    .A2(net362),
    .A3(net351),
    .S0(clknet_1_1__leaf_net355),
    .S1(clknet_1_1__leaf_net356),
    .X(net370));
 sky130_fd_sc_hd__xnor2_1 c374 (.A(net369),
    .B(net362),
    .Y(net371));
 sky130_fd_sc_hd__a21bo_1 c375 (.A1(net362),
    .A2(net364),
    .B1_N(net723),
    .X(net372));
 sky130_fd_sc_hd__a21bo_1 c376 (.A1(net371),
    .A2(net372),
    .B1_N(net723),
    .X(net373));
 sky130_fd_sc_hd__a31o_1 c377 (.A1(net363),
    .A2(net373),
    .A3(net366),
    .B1(clknet_1_1__leaf_net355),
    .X(net374));
 sky130_fd_sc_hd__dfxbp_1 c378 (.CLK(clknet_4_0_0_clk),
    .D(net247),
    .Q(net376),
    .Q_N(net375));
 sky130_fd_sc_hd__clkbuf_1 c379 (.A(net376),
    .X(net377));
 sky130_fd_sc_hd__a21bo_1 c38 (.A1(net12),
    .A2(net10),
    .B1_N(net7),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 c380 (.A(net377),
    .X(net378));
 sky130_fd_sc_hd__dlrbp_2 c381 (.D(net260),
    .GATE(clknet_4_0_0_clk),
    .RESET_B(net375),
    .Q(net380),
    .Q_N(net379));
 sky130_fd_sc_hd__sdfxtp_2 c382 (.CLK(clknet_4_0_0_clk),
    .D(net378),
    .SCD(net380),
    .SCE(net247),
    .Q(net381));
 sky130_fd_sc_hd__xnor2_4 c383 (.A(net376),
    .B(net381),
    .Y(net382));
 sky130_fd_sc_hd__xnor2_4 c384 (.A(net381),
    .B(net379),
    .Y(net383));
 sky130_fd_sc_hd__a21bo_1 c385 (.A1(net381),
    .A2(net380),
    .B1_N(net382),
    .X(net384));
 sky130_fd_sc_hd__a21bo_1 c386 (.A1(net377),
    .A2(net382),
    .B1_N(net383),
    .X(net385));
 sky130_fd_sc_hd__a21bo_2 c387 (.A1(net378),
    .A2(net383),
    .B1_N(net379),
    .X(net386));
 sky130_fd_sc_hd__xnor2_1 c388 (.A(net384),
    .B(net385),
    .Y(net387));
 sky130_fd_sc_hd__xnor2_4 c389 (.A(net382),
    .B(net386),
    .Y(net388));
 sky130_fd_sc_hd__a21bo_1 c39 (.A1(net0),
    .A2(net11),
    .B1_N(net744),
    .X(net14));
 sky130_fd_sc_hd__xnor2_4 c390 (.A(net250),
    .B(net388),
    .Y(net389));
 sky130_fd_sc_hd__xnor2_1 c391 (.A(net388),
    .B(net384),
    .Y(net390));
 sky130_fd_sc_hd__a21bo_1 c392 (.A1(net385),
    .A2(net389),
    .B1_N(net383),
    .X(net391));
 sky130_fd_sc_hd__a21bo_1 c393 (.A1(net391),
    .A2(net390),
    .B1_N(net383),
    .X(net392));
 sky130_fd_sc_hd__xnor2_2 c394 (.A(net383),
    .B(net386),
    .Y(net393));
 sky130_fd_sc_hd__xnor2_1 c395 (.A(net387),
    .B(net391),
    .Y(net394));
 sky130_fd_sc_hd__a21bo_1 c396 (.A1(net380),
    .A2(net387),
    .B1_N(net385),
    .X(net395));
 sky130_fd_sc_hd__a41o_1 c397 (.A1(net390),
    .A2(net395),
    .A3(net394),
    .A4(net389),
    .B1(net379),
    .X(net396));
 sky130_fd_sc_hd__mux4_2 c398 (.A0(net396),
    .A1(net394),
    .A2(net390),
    .A3(net383),
    .S0(net395),
    .S1(net389),
    .X(net397));
 sky130_fd_sc_hd__xnor2_1 c399 (.A(net282),
    .B(net389),
    .Y(net398));
 sky130_fd_sc_hd__a41o_1 c40 (.A1(net744),
    .A2(net12),
    .A3(net11),
    .A4(net14),
    .B1(net745),
    .X(net15));
 sky130_fd_sc_hd__xnor2_1 c400 (.A(net389),
    .B(net393),
    .Y(net399));
 sky130_fd_sc_hd__xnor2_1 c401 (.A(net397),
    .B(net399),
    .Y(net400));
 sky130_fd_sc_hd__xnor2_1 c402 (.A(clknet_1_0__leaf_net398),
    .B(net389),
    .Y(net401));
 sky130_fd_sc_hd__xnor2_1 c403 (.A(clknet_1_0__leaf_net401),
    .B(net397),
    .Y(net402));
 sky130_fd_sc_hd__xnor2_1 c404 (.A(net400),
    .B(clknet_1_1__leaf_net402),
    .Y(net403));
 sky130_fd_sc_hd__xnor2_1 c405 (.A(clknet_1_1__leaf_net398),
    .B(clknet_1_0__leaf_net402),
    .Y(net404));
 sky130_fd_sc_hd__xnor2_1 c406 (.A(clknet_1_0__leaf_net402),
    .B(net389),
    .Y(net405));
 sky130_fd_sc_hd__xnor2_1 c407 (.A(clknet_1_0__leaf_net402),
    .B(net719),
    .Y(net406));
 sky130_fd_sc_hd__xnor2_1 c408 (.A(clknet_1_1__leaf_net404),
    .B(clknet_1_0__leaf_net406),
    .Y(net407));
 sky130_fd_sc_hd__xnor2_1 c409 (.A(net400),
    .B(clknet_1_0__leaf_net404),
    .Y(net408));
 sky130_fd_sc_hd__a41o_1 c41 (.A1(net6),
    .A2(net15),
    .A3(net738),
    .A4(net745),
    .B1(net4),
    .X(net16));
 sky130_fd_sc_hd__xnor2_1 c410 (.A(clknet_1_0__leaf_net405),
    .B(clknet_1_1__leaf_net408),
    .Y(net409));
 sky130_fd_sc_hd__a21bo_1 c411 (.A1(clknet_1_1__leaf_net406),
    .A2(clknet_1_0__leaf_net409),
    .B1_N(clknet_1_0__leaf_net405),
    .X(net410));
 sky130_fd_sc_hd__a21bo_1 c412 (.A1(clknet_1_0__leaf_net408),
    .A2(clknet_1_0__leaf_net410),
    .B1_N(clknet_1_0__leaf_net405),
    .X(net411));
 sky130_fd_sc_hd__sdfxtp_1 c413 (.CLK(clknet_4_1_0_clk),
    .D(clknet_1_1__leaf_net411),
    .SCD(clknet_1_1__leaf_net407),
    .SCE(clknet_1_0__leaf_net409),
    .Q(net412));
 sky130_fd_sc_hd__a21bo_1 c414 (.A1(clknet_1_1__leaf_net410),
    .A2(clknet_1_1__leaf_net405),
    .B1_N(clknet_1_0__leaf_net408),
    .X(net413));
 sky130_fd_sc_hd__sdfbbn_1 c415 (.CLK_N(clknet_4_1_0_clk),
    .D(net399),
    .RESET_B(clknet_1_0__leaf_net411),
    .SCD(net412),
    .SCE(clknet_1_1__leaf_net413),
    .SET_B(clknet_1_1__leaf_net402),
    .Q(net415),
    .Q_N(net414));
 sky130_fd_sc_hd__dfbbn_1 c416 (.CLK_N(clknet_4_3_0_clk),
    .D(clknet_1_0__leaf_net407),
    .RESET_B(net415),
    .SET_B(clknet_1_1__leaf_net413),
    .Q(net417),
    .Q_N(net416));
 sky130_fd_sc_hd__sdfbbn_2 c417 (.CLK_N(clknet_4_3_0_clk),
    .D(net412),
    .RESET_B(clknet_1_1__leaf_net413),
    .SCD(net819),
    .SCE(clknet_1_1__leaf_net405),
    .SET_B(clknet_1_1__leaf_net402),
    .Q(net419),
    .Q_N(net418));
 sky130_fd_sc_hd__mux4_1 c418 (.A0(net417),
    .A1(net412),
    .A2(net418),
    .A3(clknet_1_1__leaf_net405),
    .S0(net414),
    .S1(clknet_1_0__leaf_net413),
    .X(net420));
 sky130_fd_sc_hd__sdfrtp_1 c419 (.CLK(clknet_4_3_0_clk),
    .D(clknet_1_1__leaf_net401),
    .RESET_B(net415),
    .SCD(clknet_1_0__leaf_net413),
    .SCE(net724),
    .Q(net421));
 sky130_fd_sc_hd__buf_2 c42 (.A(in14),
    .X(net17));
 sky130_fd_sc_hd__xnor2_2 c420 (.A(net304),
    .B(net288),
    .Y(net422));
 sky130_fd_sc_hd__buf_1 c421 (.A(net289),
    .X(net423));
 sky130_fd_sc_hd__clkbuf_1 c422 (.A(net423),
    .X(net424));
 sky130_fd_sc_hd__xnor2_1 c423 (.A(net423),
    .B(net422),
    .Y(net425));
 sky130_fd_sc_hd__xnor2_1 c424 (.A(net304),
    .B(clknet_1_1__leaf_net409),
    .Y(net426));
 sky130_fd_sc_hd__buf_1 c425 (.A(net805),
    .X(net427));
 sky130_fd_sc_hd__a21bo_1 c426 (.A1(net427),
    .A2(net425),
    .B1_N(net423),
    .X(net428));
 sky130_fd_sc_hd__dlrbp_1 c427 (.D(clknet_1_1__leaf_net413),
    .GATE(clknet_4_3_0_clk),
    .RESET_B(clknet_1_0__leaf_net426),
    .Q(net430),
    .Q_N(net429));
 sky130_fd_sc_hd__a21bo_1 c428 (.A1(net424),
    .A2(net429),
    .B1_N(net428),
    .X(net431));
 sky130_fd_sc_hd__a21bo_1 c429 (.A1(net427),
    .A2(net431),
    .B1_N(net423),
    .X(net432));
 sky130_fd_sc_hd__clkbuf_4 c43 (.A(net17),
    .X(net18));
 sky130_fd_sc_hd__xnor2_2 c430 (.A(net428),
    .B(net432),
    .Y(net433));
 sky130_fd_sc_hd__xnor2_1 c431 (.A(net432),
    .B(net429),
    .Y(net434));
 sky130_fd_sc_hd__xnor2_2 c432 (.A(net433),
    .B(net430),
    .Y(net435));
 sky130_fd_sc_hd__xnor2_1 c433 (.A(net435),
    .B(net434),
    .Y(net436));
 sky130_fd_sc_hd__a21bo_1 c434 (.A1(clknet_1_1__leaf_net403),
    .A2(net435),
    .B1_N(net433),
    .X(net437));
 sky130_fd_sc_hd__a21bo_1 c435 (.A1(net430),
    .A2(clknet_1_1__leaf_net437),
    .B1_N(net436),
    .X(net438));
 sky130_fd_sc_hd__xnor2_1 c436 (.A(clknet_1_0__leaf_net437),
    .B(net436),
    .Y(net439));
 sky130_fd_sc_hd__a21bo_1 c437 (.A1(net434),
    .A2(net428),
    .B1_N(clknet_1_0__leaf_net439),
    .X(net440));
 sky130_fd_sc_hd__a21bo_1 c438 (.A1(clknet_1_1__leaf_net426),
    .A2(net438),
    .B1_N(clknet_1_0__leaf_net440),
    .X(net441));
 sky130_fd_sc_hd__sdfbbp_1 c439 (.CLK(clknet_4_12_0_clk),
    .D(clknet_1_1__leaf_net440),
    .RESET_B(net423),
    .SCD(clknet_1_0__leaf_net441),
    .SCE(net435),
    .SET_B(net427),
    .Q(net442));
 sky130_fd_sc_hd__xnor2_1 c44 (.A(net14),
    .B(net18),
    .Y(net19));
 sky130_fd_sc_hd__dfbbn_2 c440 (.CLK_N(clknet_4_3_0_clk),
    .D(net425),
    .RESET_B(net430),
    .SET_B(clknet_1_0__leaf_net441),
    .Q(net443));
 sky130_fd_sc_hd__clkbuf_4 c441 (.A(net431),
    .X(net444));
 sky130_fd_sc_hd__buf_2 c442 (.A(net444),
    .X(net445));
 sky130_fd_sc_hd__clkbuf_4 c443 (.A(net445),
    .X(net446));
 sky130_fd_sc_hd__xnor2_4 c444 (.A(net444),
    .B(net446),
    .Y(net447));
 sky130_fd_sc_hd__xnor2_4 c445 (.A(net443),
    .B(net447),
    .Y(net448));
 sky130_fd_sc_hd__a21bo_2 c446 (.A1(net445),
    .A2(net448),
    .B1_N(net446),
    .X(net449));
 sky130_fd_sc_hd__xnor2_4 c447 (.A(net445),
    .B(net449),
    .Y(net450));
 sky130_fd_sc_hd__xnor2_1 c448 (.A(net314),
    .B(net447),
    .Y(net451));
 sky130_fd_sc_hd__xnor2_1 c449 (.A(net446),
    .B(net450),
    .Y(net452));
 sky130_fd_sc_hd__xnor2_4 c45 (.A(net18),
    .B(net17),
    .Y(net20));
 sky130_fd_sc_hd__a21bo_1 c450 (.A1(net449),
    .A2(net446),
    .B1_N(net450),
    .X(net453));
 sky130_fd_sc_hd__a21bo_1 c451 (.A1(net451),
    .A2(net450),
    .B1_N(net447),
    .X(net454));
 sky130_fd_sc_hd__xnor2_4 c452 (.A(net450),
    .B(net444),
    .Y(net455));
 sky130_fd_sc_hd__xnor2_4 c453 (.A(net442),
    .B(net455),
    .Y(net456));
 sky130_fd_sc_hd__xnor2_4 c454 (.A(net456),
    .B(net455),
    .Y(net457));
 sky130_fd_sc_hd__a21bo_1 c455 (.A1(net453),
    .A2(net454),
    .B1_N(net449),
    .X(net458));
 sky130_fd_sc_hd__mux4_1 c456 (.A0(net449),
    .A1(net457),
    .A2(net456),
    .A3(clknet_1_0__leaf_net441),
    .S0(net448),
    .S1(net450),
    .X(net459));
 sky130_fd_sc_hd__a31o_1 c457 (.A1(net445),
    .A2(net451),
    .A3(net450),
    .B1(net811),
    .X(net460));
 sky130_fd_sc_hd__a21bo_1 c458 (.A1(net312),
    .A2(net452),
    .B1_N(net460),
    .X(net461));
 sky130_fd_sc_hd__a21bo_1 c459 (.A1(net460),
    .A2(net461),
    .B1_N(net453),
    .X(net462));
 sky130_fd_sc_hd__xnor2_2 c46 (.A(net18),
    .B(net20),
    .Y(net21));
 sky130_fd_sc_hd__a21bo_1 c460 (.A1(net458),
    .A2(net462),
    .B1_N(net452),
    .X(net463));
 sky130_fd_sc_hd__dlrtn_1 c461 (.D(net454),
    .GATE_N(clknet_4_14_0_clk),
    .RESET_B(net463),
    .Q(net464));
 sky130_fd_sc_hd__dfxtp_1 c462 (.CLK(clknet_4_6_0_clk),
    .D(net328),
    .Q(net465));
 sky130_fd_sc_hd__buf_1 c463 (.A(net465),
    .X(net466));
 sky130_fd_sc_hd__xnor2_1 c464 (.A(net448),
    .B(net457),
    .Y(net467));
 sky130_fd_sc_hd__xnor2_1 c465 (.A(net466),
    .B(net457),
    .Y(net468));
 sky130_fd_sc_hd__dlrtn_1 c466 (.D(net331),
    .GATE_N(clknet_4_12_0_clk),
    .RESET_B(net467),
    .Q(net469));
 sky130_fd_sc_hd__dfbbp_1 c467 (.CLK(clknet_4_12_0_clk),
    .D(net467),
    .RESET_B(net468),
    .SET_B(net448),
    .Q(net471),
    .Q_N(net470));
 sky130_fd_sc_hd__buf_1 c468 (.A(net450),
    .X(net755));
 sky130_fd_sc_hd__xnor2_1 c469 (.A(net422),
    .B(net465),
    .Y(net472));
 sky130_fd_sc_hd__xnor2_2 c47 (.A(net21),
    .B(net20),
    .Y(net22));
 sky130_fd_sc_hd__clkbuf_1 c470 (.A(net469),
    .X(net473));
 sky130_fd_sc_hd__clkbuf_1 c471 (.A(net465),
    .X(net474));
 sky130_fd_sc_hd__dlrtn_2 c472 (.D(net347),
    .GATE_N(clknet_4_12_0_clk),
    .RESET_B(net468),
    .Q(net475));
 sky130_fd_sc_hd__xnor2_1 c473 (.A(net471),
    .B(net475),
    .Y(net476));
 sky130_fd_sc_hd__a21bo_1 c474 (.A1(net466),
    .A2(net475),
    .B1_N(net457),
    .X(net477));
 sky130_fd_sc_hd__sdfxbp_1 c475 (.CLK(clknet_4_15_0_clk),
    .D(net477),
    .SCD(net468),
    .SCE(net475),
    .Q(net478));
 sky130_fd_sc_hd__a21bo_1 c476 (.A1(net447),
    .A2(net473),
    .B1_N(net475),
    .X(net479));
 sky130_fd_sc_hd__sdfxbp_1 c477 (.CLK(clknet_4_12_0_clk),
    .D(net350),
    .SCD(net475),
    .SCE(net755),
    .Q(net480));
 sky130_fd_sc_hd__a21bo_1 c478 (.A1(net480),
    .A2(net474),
    .B1_N(net475),
    .X(net481));
 sky130_fd_sc_hd__a31o_1 c479 (.A1(net472),
    .A2(net479),
    .A3(net481),
    .B1(net475),
    .X(net482));
 sky130_fd_sc_hd__xnor2_1 c48 (.A(net13),
    .B(net21),
    .Y(net23));
 sky130_fd_sc_hd__a41o_1 c480 (.A1(net482),
    .A2(net476),
    .A3(net479),
    .A4(net481),
    .B1(net475),
    .X(net483));
 sky130_fd_sc_hd__a41o_1 c481 (.A1(net476),
    .A2(net470),
    .A3(net481),
    .A4(net475),
    .B1(net448),
    .X(net484));
 sky130_fd_sc_hd__a21bo_1 c482 (.A1(net481),
    .A2(net483),
    .B1_N(net484),
    .X(net762));
 sky130_fd_sc_hd__clkbuf_2 c487 (.A(net464),
    .X(net760));
 sky130_fd_sc_hd__dlrtp_1 c488 (.D(net374),
    .GATE(clknet_4_15_0_clk),
    .RESET_B(net832),
    .Q(net485));
 sky130_fd_sc_hd__xnor2_1 c489 (.A(net352),
    .B(net485),
    .Y(net486));
 sky130_fd_sc_hd__xnor2_1 c49 (.A(net20),
    .B(net18),
    .Y(net24));
 sky130_fd_sc_hd__buf_1 c490 (.A(net486),
    .X(net487));
 sky130_fd_sc_hd__xnor2_1 c491 (.A(net760),
    .B(net485),
    .Y(net488));
 sky130_fd_sc_hd__buf_2 c492 (.A(net487),
    .X(net489));
 sky130_fd_sc_hd__a21bo_1 c493 (.A1(net485),
    .A2(net488),
    .B1_N(net489),
    .X(net490));
 sky130_fd_sc_hd__xnor2_2 c494 (.A(net487),
    .B(net489),
    .Y(net491));
 sky130_fd_sc_hd__a21bo_2 c495 (.A1(net488),
    .A2(net490),
    .B1_N(net491),
    .X(net766));
 sky130_fd_sc_hd__a31o_1 c496 (.A1(net485),
    .A2(net491),
    .A3(net766),
    .B1(net489),
    .X(net765));
 sky130_fd_sc_hd__a31o_2 c497 (.A1(net766),
    .A2(net489),
    .A3(net487),
    .B1(net491),
    .X(net758));
 sky130_fd_sc_hd__a41o_1 c498 (.A1(net488),
    .A2(net486),
    .A3(net766),
    .A4(net758),
    .B1(net489),
    .X(net767));
 sky130_fd_sc_hd__a31o_1 c499 (.A1(net489),
    .A2(net758),
    .A3(net766),
    .B1(net491),
    .X(net764));
 sky130_fd_sc_hd__xnor2_1 c50 (.A(net7),
    .B(net22),
    .Y(net25));
 sky130_fd_sc_hd__a41o_1 c500 (.A1(net491),
    .A2(net490),
    .A3(net765),
    .A4(net758),
    .B1(net766),
    .X(net759));
 sky130_fd_sc_hd__mux4_1 c501 (.A0(net486),
    .A1(net767),
    .A2(net765),
    .A3(net764),
    .S0(net758),
    .S1(net491),
    .X(net768));
 sky130_fd_sc_hd__mux4_1 c502 (.A0(net491),
    .A1(net764),
    .A2(net489),
    .A3(net768),
    .S0(net766),
    .S1(net758),
    .X(net492));
 sky130_fd_sc_hd__mux4_1 c503 (.A0(net490),
    .A1(net492),
    .A2(net767),
    .A3(net758),
    .S0(net766),
    .S1(net489),
    .X(net763));
 sky130_fd_sc_hd__xnor2_2 c504 (.A(net392),
    .B(net389),
    .Y(net493));
 sky130_fd_sc_hd__xnor2_2 c505 (.A(net493),
    .B(net389),
    .Y(net494));
 sky130_fd_sc_hd__dlrtp_2 c506 (.D(net494),
    .GATE(clknet_4_3_0_clk),
    .RESET_B(net247),
    .Q(net495));
 sky130_fd_sc_hd__xnor2_4 c507 (.A(net495),
    .B(net774),
    .Y(net496));
 sky130_fd_sc_hd__xnor2_2 c508 (.A(net493),
    .B(net494),
    .Y(net497));
 sky130_fd_sc_hd__xnor2_4 c509 (.A(net495),
    .B(net397),
    .Y(net498));
 sky130_fd_sc_hd__xnor2_1 c51 (.A(net19),
    .B(net17),
    .Y(net26));
 sky130_fd_sc_hd__xnor2_1 c510 (.A(net774),
    .B(net772),
    .Y(net499));
 sky130_fd_sc_hd__xnor2_4 c511 (.A(net498),
    .B(net774),
    .Y(net500));
 sky130_fd_sc_hd__xnor2_1 c512 (.A(net499),
    .B(net498),
    .Y(net501));
 sky130_fd_sc_hd__xnor2_1 c513 (.A(net500),
    .B(net774),
    .Y(net502));
 sky130_fd_sc_hd__xnor2_1 c514 (.A(net501),
    .B(net499),
    .Y(net503));
 sky130_fd_sc_hd__xnor2_4 c515 (.A(net497),
    .B(net500),
    .Y(net504));
 sky130_fd_sc_hd__xnor2_1 c516 (.A(net503),
    .B(net504),
    .Y(net505));
 sky130_fd_sc_hd__xnor2_1 c517 (.A(net393),
    .B(net504),
    .Y(net506));
 sky130_fd_sc_hd__a41o_1 c518 (.A1(net505),
    .A2(net503),
    .A3(net504),
    .A4(net772),
    .B1(net774),
    .X(net507));
 sky130_fd_sc_hd__dlrtp_1 c519 (.D(net507),
    .GATE(clknet_4_2_0_clk),
    .RESET_B(net502),
    .Q(net508));
 sky130_fd_sc_hd__a21bo_1 c52 (.A1(net24),
    .A2(net20),
    .B1_N(net18),
    .X(net27));
 sky130_fd_sc_hd__xnor2_1 c520 (.A(net392),
    .B(net504),
    .Y(net509));
 sky130_fd_sc_hd__a21bo_2 c521 (.A1(net509),
    .A2(net792),
    .B1_N(net506),
    .X(net510));
 sky130_fd_sc_hd__a41o_1 c522 (.A1(net506),
    .A2(net502),
    .A3(net510),
    .A4(net504),
    .B1(net772),
    .X(net511));
 sky130_fd_sc_hd__edfxbp_1 c523 (.CLK(clknet_4_2_0_clk),
    .D(net511),
    .DE(net505),
    .Q(net512));
 sky130_fd_sc_hd__xnor2_4 c524 (.A(net791),
    .B(net510),
    .Y(net513));
 sky130_fd_sc_hd__xnor2_4 c525 (.A(net397),
    .B(net724),
    .Y(net514));
 sky130_fd_sc_hd__clkbuf_2 c526 (.A(net514),
    .X(net515));
 sky130_fd_sc_hd__xnor2_4 c527 (.A(net514),
    .B(net773),
    .Y(net516));
 sky130_fd_sc_hd__edfxtp_1 c528 (.CLK(clknet_4_2_0_clk),
    .D(net513),
    .DE(net516),
    .Q(net517));
 sky130_fd_sc_hd__xnor2_4 c529 (.A(net517),
    .B(net514),
    .Y(net518));
 sky130_fd_sc_hd__a21bo_1 c53 (.A1(net25),
    .A2(net22),
    .B1_N(net27),
    .X(net28));
 sky130_fd_sc_hd__xnor2_2 c530 (.A(net277),
    .B(net517),
    .Y(net519));
 sky130_fd_sc_hd__xnor2_1 c531 (.A(net514),
    .B(net516),
    .Y(net520));
 sky130_fd_sc_hd__xnor2_1 c532 (.A(net516),
    .B(net519),
    .Y(net521));
 sky130_fd_sc_hd__sdlclkp_1 c533 (.CLK(clknet_4_3_0_clk),
    .GATE(net267),
    .SCE(net519),
    .GCLK(net522));
 sky130_fd_sc_hd__xnor2_1 c534 (.A(net519),
    .B(net518),
    .Y(net523));
 sky130_fd_sc_hd__a21bo_1 c535 (.A1(net521),
    .A2(net496),
    .B1_N(net518),
    .X(net524));
 sky130_fd_sc_hd__xnor2_4 c536 (.A(net515),
    .B(net518),
    .Y(net525));
 sky130_fd_sc_hd__xnor2_1 c537 (.A(net517),
    .B(net771),
    .Y(net526));
 sky130_fd_sc_hd__a21bo_1 c538 (.A1(net522),
    .A2(net525),
    .B1_N(net516),
    .X(net527));
 sky130_fd_sc_hd__sdfxtp_1 c539 (.CLK(clknet_4_3_0_clk),
    .D(net524),
    .SCD(net526),
    .SCE(clknet_1_0__leaf_net413),
    .Q(net528));
 sky130_fd_sc_hd__a21bo_1 c54 (.A1(net20),
    .A2(net24),
    .B1_N(net22),
    .X(net29));
 sky130_fd_sc_hd__a21bo_1 c540 (.A1(net527),
    .A2(net514),
    .B1_N(net519),
    .X(net529));
 sky130_fd_sc_hd__a21bo_1 c541 (.A1(clknet_1_1__leaf_net409),
    .A2(net525),
    .B1_N(net518),
    .X(net530));
 sky130_fd_sc_hd__a31o_1 c542 (.A1(net520),
    .A2(clknet_1_0__leaf_net530),
    .A3(net517),
    .B1(net525),
    .X(net531));
 sky130_fd_sc_hd__sdfrtp_1 c543 (.CLK(clknet_4_2_0_clk),
    .D(net518),
    .RESET_B(net531),
    .SCD(clknet_1_0__leaf_net530),
    .SCE(net517),
    .Q(net532));
 sky130_fd_sc_hd__a31o_1 c544 (.A1(net532),
    .A2(clknet_1_1__leaf_net530),
    .A3(net519),
    .B1(net516),
    .X(net533));
 sky130_fd_sc_hd__sdfsbp_1 c545 (.CLK(clknet_4_3_0_clk),
    .D(net533),
    .SCD(net529),
    .SCE(clknet_1_0__leaf_net403),
    .SET_B(clknet_1_1__leaf_net530),
    .Q(net534));
 sky130_fd_sc_hd__dfxtp_2 c546 (.CLK(clknet_4_9_0_clk),
    .D(clknet_1_0__leaf_net441),
    .Q(net535));
 sky130_fd_sc_hd__clkbuf_4 c547 (.A(net535),
    .X(net536));
 sky130_fd_sc_hd__xnor2_1 c548 (.A(net536),
    .B(net535),
    .Y(net537));
 sky130_fd_sc_hd__xnor2_4 c549 (.A(net419),
    .B(net496),
    .Y(net538));
 sky130_fd_sc_hd__xnor2_1 c55 (.A(net28),
    .B(net733),
    .Y(net30));
 sky130_fd_sc_hd__a21bo_2 c550 (.A1(net535),
    .A2(net538),
    .B1_N(net536),
    .X(net539));
 sky130_fd_sc_hd__xnor2_1 c551 (.A(net536),
    .B(net535),
    .Y(net540));
 sky130_fd_sc_hd__xnor2_2 c552 (.A(net539),
    .B(net536),
    .Y(net541));
 sky130_fd_sc_hd__a21bo_1 c553 (.A1(net537),
    .A2(net541),
    .B1_N(net539),
    .X(net542));
 sky130_fd_sc_hd__xnor2_1 c554 (.A(net538),
    .B(net539),
    .Y(net543));
 sky130_fd_sc_hd__xnor2_1 c555 (.A(net541),
    .B(net539),
    .Y(net544));
 sky130_fd_sc_hd__xnor2_1 c556 (.A(net542),
    .B(net539),
    .Y(net545));
 sky130_fd_sc_hd__a21bo_1 c557 (.A1(net544),
    .A2(net538),
    .B1_N(net536),
    .X(net546));
 sky130_fd_sc_hd__mux4_1 c558 (.A0(net546),
    .A1(net538),
    .A2(clknet_1_0__leaf_net439),
    .A3(net539),
    .S0(net525),
    .S1(net535),
    .X(net547));
 sky130_fd_sc_hd__a21bo_2 c559 (.A1(net523),
    .A2(net542),
    .B1_N(net536),
    .X(net548));
 sky130_fd_sc_hd__a21bo_1 c56 (.A1(net23),
    .A2(net27),
    .B1_N(net25),
    .X(net31));
 sky130_fd_sc_hd__sdfxtp_1 c560 (.CLK(clknet_4_9_0_clk),
    .D(net543),
    .SCD(net541),
    .SCE(net548),
    .Q(net549));
 sky130_fd_sc_hd__sdfxtp_1 c561 (.CLK(clknet_4_9_0_clk),
    .D(net796),
    .SCD(net548),
    .SCE(net805),
    .Q(net550));
 sky130_fd_sc_hd__dfbbn_1 c562 (.CLK_N(clknet_4_9_0_clk),
    .D(net538),
    .RESET_B(net550),
    .SET_B(net548),
    .Q(net551));
 sky130_fd_sc_hd__dfbbn_1 c563 (.CLK_N(clknet_4_9_0_clk),
    .D(net550),
    .RESET_B(net546),
    .SET_B(net548),
    .Q(net553),
    .Q_N(net552));
 sky130_fd_sc_hd__a21bo_1 c564 (.A1(net553),
    .A2(net535),
    .B1_N(net541),
    .X(net554));
 sky130_fd_sc_hd__a21bo_1 c565 (.A1(net525),
    .A2(net553),
    .B1_N(net550),
    .X(net555));
 sky130_fd_sc_hd__a41o_1 c566 (.A1(net554),
    .A2(net555),
    .A3(net552),
    .A4(net539),
    .B1(net538),
    .X(net556));
 sky130_fd_sc_hd__clkbuf_1 c567 (.A(net457),
    .X(net557));
 sky130_fd_sc_hd__sdlclkp_2 c568 (.CLK(clknet_4_9_0_clk),
    .GATE(net548),
    .SCE(net536),
    .GCLK(net558));
 sky130_fd_sc_hd__sdlclkp_4 c569 (.CLK(clknet_4_9_0_clk),
    .GATE(net545),
    .SCE(net447),
    .GCLK(net559));
 sky130_fd_sc_hd__a21bo_1 c57 (.A1(net31),
    .A2(net29),
    .B1_N(net19),
    .X(net32));
 sky130_fd_sc_hd__xnor2_1 c570 (.A(clknet_1_0__leaf_net559),
    .B(net525),
    .Y(net560));
 sky130_fd_sc_hd__xnor2_1 c571 (.A(clknet_1_1__leaf_net558),
    .B(net446),
    .Y(net561));
 sky130_fd_sc_hd__xnor2_1 c572 (.A(net561),
    .B(clknet_1_0__leaf_net558),
    .Y(net562));
 sky130_fd_sc_hd__xnor2_1 c573 (.A(net446),
    .B(clknet_1_0__leaf_net559),
    .Y(net563));
 sky130_fd_sc_hd__xnor2_1 c574 (.A(net563),
    .B(net536),
    .Y(net564));
 sky130_fd_sc_hd__xnor2_1 c575 (.A(clknet_1_1__leaf_net564),
    .B(clknet_1_1__leaf_net562),
    .Y(net565));
 sky130_fd_sc_hd__xnor2_1 c576 (.A(clknet_1_0__leaf_net565),
    .B(clknet_1_0__leaf_net562),
    .Y(net770));
 sky130_fd_sc_hd__dfrbp_1 c577 (.CLK(clknet_4_14_0_clk),
    .D(net557),
    .RESET_B(clknet_1_1__leaf_net565),
    .Q(net567),
    .Q_N(net566));
 sky130_fd_sc_hd__xnor2_1 c578 (.A(net560),
    .B(clknet_1_0__leaf_net558),
    .Y(net568));
 sky130_fd_sc_hd__dfbbp_1 c579 (.CLK(clknet_4_9_0_clk),
    .D(net568),
    .RESET_B(net826),
    .SET_B(net548),
    .Q(net570),
    .Q_N(net569));
 sky130_fd_sc_hd__a21bo_1 c58 (.A1(net22),
    .A2(net24),
    .B1_N(net25),
    .X(net33));
 sky130_fd_sc_hd__xnor2_1 c580 (.A(clknet_1_1__leaf_net439),
    .B(net569),
    .Y(net571));
 sky130_fd_sc_hd__a31o_1 c581 (.A1(net567),
    .A2(clknet_1_1__leaf_net562),
    .A3(clknet_1_0__leaf_net564),
    .B1(net569),
    .X(net572));
 sky130_fd_sc_hd__xnor2_1 c582 (.A(clknet_1_1__leaf_net559),
    .B(clknet_1_1__leaf_net565),
    .Y(net573));
 sky130_fd_sc_hd__a21bo_1 c583 (.A1(net536),
    .A2(net570),
    .B1_N(clknet_1_0__leaf_net573),
    .X(net574));
 sky130_fd_sc_hd__a31o_1 c584 (.A1(net574),
    .A2(net567),
    .A3(clknet_1_0__leaf_net571),
    .B1(clknet_1_0__leaf_net573),
    .X(net761));
 sky130_fd_sc_hd__a31o_1 c585 (.A1(clknet_1_1__leaf_net571),
    .A2(clknet_1_0__leaf_net565),
    .A3(clknet_1_0__leaf_net573),
    .B1(clknet_1_0__leaf_net562),
    .X(net575));
 sky130_fd_sc_hd__dfrbp_1 c586 (.CLK(clknet_4_9_0_clk),
    .D(net816),
    .RESET_B(net575),
    .Q(net576));
 sky130_fd_sc_hd__xnor2_1 c587 (.A(net572),
    .B(net576),
    .Y(net577));
 sky130_fd_sc_hd__buf_1 c588 (.A(clknet_1_1__leaf_net573),
    .X(net578));
 sky130_fd_sc_hd__clkbuf_2 c589 (.A(net478),
    .X(net579));
 sky130_fd_sc_hd__a21bo_1 c59 (.A1(net32),
    .A2(net30),
    .B1_N(net33),
    .X(net34));
 sky130_fd_sc_hd__buf_1 c590 (.A(clknet_1_0__leaf_net578),
    .X(net580));
 sky130_fd_sc_hd__xnor2_1 c591 (.A(net579),
    .B(clknet_1_1__leaf_net573),
    .Y(net581));
 sky130_fd_sc_hd__xnor2_1 c592 (.A(net579),
    .B(clknet_1_0__leaf_net581),
    .Y(net582));
 sky130_fd_sc_hd__xnor2_1 c593 (.A(clknet_1_0__leaf_net582),
    .B(clknet_1_0__leaf_net580),
    .Y(net583));
 sky130_fd_sc_hd__xnor2_1 c594 (.A(net551),
    .B(clknet_1_1__leaf_net580),
    .Y(net584));
 sky130_fd_sc_hd__xnor2_1 c595 (.A(clknet_1_0__leaf_net582),
    .B(clknet_1_1__leaf_net584),
    .Y(net585));
 sky130_fd_sc_hd__xnor2_1 c596 (.A(clknet_1_0__leaf_net584),
    .B(net579),
    .Y(net586));
 sky130_fd_sc_hd__sdfxbp_1 c597 (.CLK(clknet_4_15_0_clk),
    .D(net583),
    .SCD(clknet_1_0__leaf_net580),
    .SCE(clknet_1_0__leaf_net585),
    .Q(net588),
    .Q_N(net587));
 sky130_fd_sc_hd__dfrtn_1 c598 (.CLK_N(clknet_4_15_0_clk),
    .D(clknet_1_0__leaf_net585),
    .RESET_B(net588),
    .Q(net589));
 sky130_fd_sc_hd__xnor2_1 c599 (.A(net579),
    .B(clknet_1_1__leaf_net582),
    .Y(net756));
 sky130_fd_sc_hd__mux4_1 c60 (.A0(net30),
    .A1(net33),
    .A2(net28),
    .A3(net18),
    .S0(net27),
    .S1(net20),
    .X(net35));
 sky130_fd_sc_hd__dfrtp_1 c600 (.CLK(clknet_4_14_0_clk),
    .D(net586),
    .RESET_B(clknet_1_0__leaf_net578),
    .Q(net590));
 sky130_fd_sc_hd__sdfxbp_1 c601 (.CLK(clknet_4_15_0_clk),
    .D(clknet_1_1__leaf_net581),
    .SCD(clknet_1_1__leaf_net585),
    .SCE(net820),
    .Q(net592),
    .Q_N(net591));
 sky130_fd_sc_hd__a21bo_1 c602 (.A1(net588),
    .A2(net591),
    .B1_N(clknet_1_0__leaf_net756),
    .X(net593));
 sky130_fd_sc_hd__sdfxtp_1 c603 (.CLK(clknet_4_14_0_clk),
    .D(net589),
    .SCD(net593),
    .SCE(clknet_1_0__leaf_net756),
    .Q(net594));
 sky130_fd_sc_hd__a21bo_1 c604 (.A1(net590),
    .A2(net594),
    .B1_N(clknet_1_0__leaf_net756),
    .X(net595));
 sky130_fd_sc_hd__sdfxtp_1 c605 (.CLK(clknet_4_14_0_clk),
    .D(clknet_1_1__leaf_net580),
    .SCD(net595),
    .SCE(net814),
    .Q(net596));
 sky130_fd_sc_hd__mux4_1 c606 (.A0(net596),
    .A1(net589),
    .A2(net594),
    .A3(clknet_1_1__leaf_net582),
    .S0(clknet_1_1__leaf_net578),
    .S1(clknet_1_0__leaf_net756),
    .X(net597));
 sky130_fd_sc_hd__sdfbbn_1 c607 (.CLK_N(clknet_4_14_0_clk),
    .D(net597),
    .RESET_B(net592),
    .SCD(net587),
    .SCE(net594),
    .SET_B(clknet_1_0__leaf_net756),
    .Q(net598));
 sky130_fd_sc_hd__a31o_1 c608 (.A1(clknet_1_1__leaf_net578),
    .A2(net598),
    .A3(net590),
    .B1(clknet_1_0__leaf_net756),
    .X(net757));
 sky130_fd_sc_hd__a21bo_1 c61 (.A1(net27),
    .A2(net35),
    .B1_N(net29),
    .X(net36));
 sky130_fd_sc_hd__a41o_1 c62 (.A1(net36),
    .A2(net29),
    .A3(net28),
    .A4(net33),
    .B1(net20),
    .X(net37));
 sky130_fd_sc_hd__buf_1 c63 (.A(net40),
    .X(net38));
 sky130_fd_sc_hd__dfxtp_2 c630 (.CLK(clknet_4_2_0_clk),
    .D(net513),
    .Q(net599));
 sky130_fd_sc_hd__dfrtp_4 c631 (.CLK(clknet_4_2_0_clk),
    .D(net802),
    .RESET_B(net513),
    .Q(net600));
 sky130_fd_sc_hd__xnor2_4 c632 (.A(net599),
    .B(net600),
    .Y(net601));
 sky130_fd_sc_hd__dfrtp_2 c633 (.CLK(clknet_4_2_0_clk),
    .D(net601),
    .RESET_B(net513),
    .Q(net602));
 sky130_fd_sc_hd__xnor2_4 c634 (.A(net602),
    .B(net601),
    .Y(net603));
 sky130_fd_sc_hd__xnor2_1 c635 (.A(net601),
    .B(net600),
    .Y(net604));
 sky130_fd_sc_hd__xnor2_2 c636 (.A(net600),
    .B(net603),
    .Y(net605));
 sky130_fd_sc_hd__dfsbp_1 c637 (.CLK(clknet_4_2_0_clk),
    .D(net802),
    .SET_B(net513),
    .Q(net607),
    .Q_N(net606));
 sky130_fd_sc_hd__xnor2_2 c638 (.A(net772),
    .B(net600),
    .Y(net608));
 sky130_fd_sc_hd__xnor2_4 c639 (.A(net608),
    .B(net603),
    .Y(net609));
 sky130_fd_sc_hd__clkbuf_1 c64 (.A(net40),
    .X(net39));
 sky130_fd_sc_hd__a21bo_2 c640 (.A1(net605),
    .A2(net599),
    .B1_N(net609),
    .X(net610));
 sky130_fd_sc_hd__xnor2_4 c641 (.A(net610),
    .B(net609),
    .Y(net611));
 sky130_fd_sc_hd__a21bo_1 c642 (.A1(net603),
    .A2(net604),
    .B1_N(net611),
    .X(net612));
 sky130_fd_sc_hd__a21bo_1 c643 (.A1(net602),
    .A2(net605),
    .B1_N(net772),
    .X(net613));
 sky130_fd_sc_hd__sdfsbp_1 c644 (.CLK(clknet_4_2_0_clk),
    .D(net604),
    .SCD(net612),
    .SCE(net513),
    .SET_B(net611),
    .Q(net614));
 sky130_fd_sc_hd__sdfbbn_1 c645 (.CLK_N(clknet_4_2_0_clk),
    .D(net612),
    .RESET_B(net614),
    .SCD(net607),
    .SCE(net610),
    .SET_B(net605),
    .Q(net615));
 sky130_fd_sc_hd__a21bo_1 c646 (.A1(net600),
    .A2(net611),
    .B1_N(net610),
    .X(net616));
 sky130_fd_sc_hd__sdfxtp_1 c647 (.CLK(clknet_4_2_0_clk),
    .D(net616),
    .SCD(net612),
    .SCE(net610),
    .Q(net617));
 sky130_fd_sc_hd__dfbbn_1 c648 (.CLK_N(clknet_4_2_0_clk),
    .D(net613),
    .RESET_B(net617),
    .SET_B(net612),
    .Q(net618));
 sky130_fd_sc_hd__sdfbbp_1 c649 (.CLK(clknet_4_2_0_clk),
    .D(net618),
    .RESET_B(net615),
    .SCD(net798),
    .SCE(net616),
    .SET_B(net834),
    .Q(net619));
 sky130_fd_sc_hd__buf_1 c65 (.A(net34),
    .X(net40));
 sky130_fd_sc_hd__sdfbbn_2 c650 (.CLK_N(clknet_4_2_0_clk),
    .D(net619),
    .RESET_B(net609),
    .SCD(net616),
    .SCE(net617),
    .SET_B(net606),
    .Q(net621),
    .Q_N(net620));
 sky130_fd_sc_hd__xnor2_4 c651 (.A(net621),
    .B(net771),
    .Y(net622));
 sky130_fd_sc_hd__xnor2_4 c652 (.A(net622),
    .B(net771),
    .Y(net623));
 sky130_fd_sc_hd__xnor2_4 c653 (.A(net611),
    .B(net622),
    .Y(net624));
 sky130_fd_sc_hd__dfsbp_1 c654 (.CLK(clknet_4_2_0_clk),
    .D(net623),
    .SET_B(net624),
    .Q(net626),
    .Q_N(net625));
 sky130_fd_sc_hd__xnor2_1 c655 (.A(net623),
    .B(net621),
    .Y(net627));
 sky130_fd_sc_hd__dfstp_1 c656 (.CLK(clknet_4_8_0_clk),
    .D(net624),
    .SET_B(net622),
    .Q(net628));
 sky130_fd_sc_hd__xnor2_1 c657 (.A(net827),
    .B(net623),
    .Y(net629));
 sky130_fd_sc_hd__dfstp_1 c658 (.CLK(clknet_4_2_0_clk),
    .D(net798),
    .SET_B(net624),
    .Q(net630));
 sky130_fd_sc_hd__dfstp_1 c659 (.CLK(clknet_4_8_0_clk),
    .D(net808),
    .SET_B(net629),
    .Q(net631));
 sky130_fd_sc_hd__buf_1 c66 (.A(net40),
    .X(net41));
 sky130_fd_sc_hd__a21bo_1 c660 (.A1(net631),
    .A2(net804),
    .B1_N(net623),
    .X(net632));
 sky130_fd_sc_hd__dfbbn_1 c661 (.CLK_N(clknet_4_8_0_clk),
    .D(net528),
    .RESET_B(net631),
    .SET_B(net629),
    .Q(net633));
 sky130_fd_sc_hd__dfbbp_1 c662 (.CLK(clknet_4_8_0_clk),
    .D(net629),
    .RESET_B(net623),
    .SET_B(net632),
    .Q(net635),
    .Q_N(net634));
 sky130_fd_sc_hd__sdfxbp_1 c663 (.CLK(clknet_4_8_0_clk),
    .D(net627),
    .SCD(net635),
    .SCE(net831),
    .Q(net637),
    .Q_N(net636));
 sky130_fd_sc_hd__a21bo_1 c664 (.A1(net534),
    .A2(net635),
    .B1_N(net636),
    .X(net638));
 sky130_fd_sc_hd__sdfxbp_1 c665 (.CLK(clknet_4_8_0_clk),
    .D(net638),
    .SCD(net810),
    .SCE(net632),
    .Q(net640),
    .Q_N(net639));
 sky130_fd_sc_hd__a41o_1 c666 (.A1(net628),
    .A2(net638),
    .A3(net620),
    .A4(net639),
    .B1(net623),
    .X(net641));
 sky130_fd_sc_hd__a21bo_1 c667 (.A1(net607),
    .A2(net637),
    .B1_N(net638),
    .X(net642));
 sky130_fd_sc_hd__sdfxtp_1 c668 (.CLK(clknet_4_8_0_clk),
    .D(net632),
    .SCD(net641),
    .SCE(net630),
    .Q(net643));
 sky130_fd_sc_hd__sdfbbn_1 c669 (.CLK_N(clknet_4_8_0_clk),
    .D(net643),
    .RESET_B(net642),
    .SCD(net630),
    .SCE(net624),
    .SET_B(net623),
    .Q(net644));
 sky130_fd_sc_hd__buf_4 c67 (.A(net41),
    .X(net42));
 sky130_fd_sc_hd__mux4_1 c670 (.A0(net633),
    .A1(net640),
    .A2(net634),
    .A3(net628),
    .S0(net623),
    .S1(net638),
    .X(net645));
 sky130_fd_sc_hd__sdfbbp_1 c671 (.CLK(clknet_4_8_0_clk),
    .D(net644),
    .RESET_B(net645),
    .SCD(net823),
    .SCE(net807),
    .SET_B(net623),
    .Q(net646));
 sky130_fd_sc_hd__dlclkp_1 c672 (.CLK(clknet_4_8_0_clk),
    .GATE(net556),
    .GCLK(net647));
 sky130_fd_sc_hd__buf_1 c673 (.A(clknet_1_0__leaf_net647),
    .X(net648));
 sky130_fd_sc_hd__dlrbn_1 c674 (.D(net830),
    .GATE_N(clknet_4_8_0_clk),
    .RESET_B(net556),
    .Q(net649));
 sky130_fd_sc_hd__dlclkp_2 c675 (.CLK(clknet_4_8_0_clk),
    .GATE(net624),
    .GCLK(net650));
 sky130_fd_sc_hd__buf_1 c676 (.A(clknet_1_1__leaf_net650),
    .X(net651));
 sky130_fd_sc_hd__xnor2_1 c677 (.A(clknet_1_0__leaf_net648),
    .B(clknet_1_0__leaf_net650),
    .Y(net652));
 sky130_fd_sc_hd__xnor2_1 c678 (.A(net540),
    .B(clknet_1_1__leaf_net652),
    .Y(net653));
 sky130_fd_sc_hd__xnor2_1 c679 (.A(clknet_1_1__leaf_net651),
    .B(clknet_1_1__leaf_net652),
    .Y(net654));
 sky130_fd_sc_hd__clkbuf_1 c68 (.A(net42),
    .X(net43));
 sky130_fd_sc_hd__xnor2_1 c680 (.A(clknet_1_0__leaf_net651),
    .B(clknet_1_0__leaf_net652),
    .Y(net655));
 sky130_fd_sc_hd__a21bo_1 c681 (.A1(clknet_1_1__leaf_net651),
    .A2(clknet_1_1__leaf_net654),
    .B1_N(net726),
    .X(net656));
 sky130_fd_sc_hd__xnor2_1 c682 (.A(clknet_1_1__leaf_net652),
    .B(clknet_1_0__leaf_net656),
    .Y(net657));
 sky130_fd_sc_hd__xnor2_1 c683 (.A(clknet_1_1__leaf_net647),
    .B(clknet_1_0__leaf_net654),
    .Y(net658));
 sky130_fd_sc_hd__a21bo_1 c684 (.A1(clknet_1_0__leaf_net653),
    .A2(clknet_1_0__leaf_net652),
    .B1_N(clknet_1_0__leaf_net654),
    .X(net659));
 sky130_fd_sc_hd__a31o_1 c685 (.A1(net649),
    .A2(clknet_1_0__leaf_net651),
    .A3(clknet_1_0__leaf_net648),
    .B1(clknet_1_0__leaf_net653),
    .X(net660));
 sky130_fd_sc_hd__sdfxtp_1 c686 (.CLK(clknet_4_11_0_clk),
    .D(clknet_1_1__leaf_net655),
    .SCD(clknet_1_1__leaf_net660),
    .SCE(net556),
    .Q(net661));
 sky130_fd_sc_hd__a31o_1 c687 (.A1(clknet_1_0__leaf_net659),
    .A2(clknet_1_0__leaf_net653),
    .A3(clknet_1_0__leaf_net655),
    .B1(clknet_1_1__leaf_net648),
    .X(net662));
 sky130_fd_sc_hd__a21bo_1 c688 (.A1(clknet_1_1__leaf_net654),
    .A2(clknet_1_1__leaf_net662),
    .B1_N(clknet_1_1__leaf_net653),
    .X(net663));
 sky130_fd_sc_hd__xnor2_1 c689 (.A(clknet_1_0__leaf_net662),
    .B(clknet_1_0__leaf_net652),
    .Y(net664));
 sky130_fd_sc_hd__xnor2_1 c69 (.A(net37),
    .B(net42),
    .Y(net44));
 sky130_fd_sc_hd__a21bo_1 c690 (.A1(net658),
    .A2(clknet_1_0__leaf_net660),
    .B1_N(clknet_1_0__leaf_net664),
    .X(net665));
 sky130_fd_sc_hd__a41o_1 c691 (.A1(clknet_1_0__leaf_net663),
    .A2(clknet_1_1__leaf_net664),
    .A3(clknet_1_1__leaf_net659),
    .A4(clknet_1_1__leaf_net648),
    .B1(clknet_1_0__leaf_net652),
    .X(net666));
 sky130_fd_sc_hd__a31o_1 c692 (.A1(net657),
    .A2(net666),
    .A3(clknet_1_1__leaf_net653),
    .B1(clknet_1_1__leaf_net663),
    .X(net667));
 sky130_fd_sc_hd__xnor2_1 c693 (.A(net577),
    .B(clknet_1_1__leaf_net656),
    .Y(net668));
 sky130_fd_sc_hd__xnor2_1 c694 (.A(net452),
    .B(clknet_1_1__leaf_net573),
    .Y(net669));
 sky130_fd_sc_hd__dlrbn_1 c695 (.D(clknet_1_0__leaf_net761),
    .GATE_N(clknet_4_11_0_clk),
    .RESET_B(clknet_1_0__leaf_net668),
    .Q(net671),
    .Q_N(net670));
 sky130_fd_sc_hd__xnor2_1 c696 (.A(net665),
    .B(net815),
    .Y(net672));
 sky130_fd_sc_hd__xnor2_1 c697 (.A(clknet_1_1__leaf_net672),
    .B(clknet_1_0__leaf_net669),
    .Y(net673));
 sky130_fd_sc_hd__dlrbp_1 c698 (.D(clknet_1_1__leaf_net441),
    .GATE(clknet_4_11_0_clk),
    .RESET_B(net815),
    .Q(net675),
    .Q_N(net674));
 sky130_fd_sc_hd__xnor2_1 c699 (.A(clknet_1_0__leaf_net668),
    .B(net815),
    .Y(net676));
 sky130_fd_sc_hd__dfrbp_1 c70 (.CLK(clknet_4_4_0_clk),
    .D(net43),
    .RESET_B(net38),
    .Q(net46),
    .Q_N(net45));
 sky130_fd_sc_hd__a21bo_1 c700 (.A1(clknet_1_0__leaf_net673),
    .A2(net674),
    .B1_N(net815),
    .X(net677));
 sky130_fd_sc_hd__dlrbp_1 c701 (.D(clknet_1_0__leaf_net677),
    .GATE(clknet_4_11_0_clk),
    .RESET_B(clknet_1_1__leaf_net668),
    .Q(net679),
    .Q_N(net678));
 sky130_fd_sc_hd__xnor2_1 c702 (.A(clknet_1_0__leaf_net676),
    .B(net667),
    .Y(net680));
 sky130_fd_sc_hd__xnor2_1 c703 (.A(clknet_1_0__leaf_net656),
    .B(clknet_1_0__leaf_net680),
    .Y(net681));
 sky130_fd_sc_hd__sdfbbn_1 c704 (.CLK_N(clknet_4_11_0_clk),
    .D(clknet_1_0__leaf_net672),
    .RESET_B(clknet_1_1__leaf_net668),
    .SCD(net678),
    .SCE(clknet_1_0__leaf_net681),
    .SET_B(net670),
    .Q(net683),
    .Q_N(net682));
 sky130_fd_sc_hd__sdfxtp_1 c705 (.CLK(clknet_4_11_0_clk),
    .D(net671),
    .SCD(clknet_1_0__leaf_net681),
    .SCE(clknet_1_0__leaf_net680),
    .Q(net684));
 sky130_fd_sc_hd__mux4_1 c706 (.A0(net684),
    .A1(clknet_1_0__leaf_net681),
    .A2(clknet_1_0__leaf_net676),
    .A3(clknet_1_0__leaf_net673),
    .S0(net682),
    .S1(net670),
    .X(net685));
 sky130_fd_sc_hd__dfbbn_1 c707 (.CLK_N(clknet_4_10_0_clk),
    .D(net684),
    .RESET_B(clknet_1_1__leaf_net681),
    .SET_B(net727),
    .Q(net687),
    .Q_N(net686));
 sky130_fd_sc_hd__dfbbn_1 c708 (.CLK_N(clknet_4_11_0_clk),
    .D(clknet_1_1__leaf_net680),
    .RESET_B(clknet_1_0__leaf_net681),
    .SET_B(clknet_1_1__leaf_net677),
    .Q(net689),
    .Q_N(net688));
 sky130_fd_sc_hd__a21bo_1 c709 (.A1(net675),
    .A2(net679),
    .B1_N(net688),
    .X(net690));
 sky130_fd_sc_hd__a21bo_1 c71 (.A1(net803),
    .A2(net42),
    .B1_N(net41),
    .X(net47));
 sky130_fd_sc_hd__dfbbp_1 c710 (.CLK(clknet_4_10_0_clk),
    .D(net687),
    .RESET_B(net683),
    .SET_B(clknet_1_1__leaf_net681),
    .Q(net691));
 sky130_fd_sc_hd__mux4_1 c711 (.A0(net661),
    .A1(net691),
    .A2(net683),
    .A3(net684),
    .S0(net670),
    .S1(clknet_1_0__leaf_net673),
    .X(net692));
 sky130_fd_sc_hd__mux4_1 c712 (.A0(clknet_1_1__leaf_net669),
    .A1(net690),
    .A2(net686),
    .A3(clknet_1_0__leaf_net692),
    .S0(clknet_1_1__leaf_net676),
    .S1(net670),
    .X(net693));
 sky130_fd_sc_hd__sdfxbp_1 c713 (.CLK(clknet_4_11_0_clk),
    .D(net689),
    .SCD(clknet_1_1__leaf_net692),
    .SCE(net806),
    .Q(net695),
    .Q_N(net694));
 sky130_fd_sc_hd__sdfxbp_1 c714 (.CLK(clknet_4_10_0_clk),
    .D(clknet_1_0__leaf_net757),
    .SCD(net817),
    .SCE(clknet_1_0__leaf_net756),
    .Q(net697),
    .Q_N(net696));
 sky130_fd_sc_hd__xnor2_1 c715 (.A(net697),
    .B(clknet_1_1__leaf_net673),
    .Y(net698));
 sky130_fd_sc_hd__dlrtn_1 c716 (.D(clknet_1_0__leaf_net698),
    .GATE_N(clknet_4_10_0_clk),
    .RESET_B(net793),
    .Q(net699));
 sky130_fd_sc_hd__sdfxtp_1 c717 (.CLK(clknet_4_11_0_clk),
    .D(clknet_1_1__leaf_net681),
    .SCD(net813),
    .SCE(net699),
    .Q(net700));
 sky130_fd_sc_hd__xnor2_2 c718 (.A(net699),
    .B(net700),
    .Y(net701));
 sky130_fd_sc_hd__sdfxtp_1 c719 (.CLK(clknet_4_10_0_clk),
    .D(clknet_1_0__leaf_net698),
    .SCD(net701),
    .SCE(net699),
    .Q(net702));
 sky130_fd_sc_hd__dfbbn_1 c72 (.CLK_N(clknet_4_4_0_clk),
    .D(net47),
    .RESET_B(net45),
    .SET_B(net42),
    .Q(net49),
    .Q_N(net48));
 sky130_fd_sc_hd__a21bo_1 c720 (.A1(net813),
    .A2(net695),
    .B1_N(net702),
    .X(net703));
 sky130_fd_sc_hd__a21bo_1 c721 (.A1(clknet_1_1__leaf_net673),
    .A2(net702),
    .B1_N(net701),
    .X(net704));
 sky130_fd_sc_hd__a21bo_1 c722 (.A1(net702),
    .A2(net825),
    .B1_N(clknet_1_1__leaf_net756),
    .X(net705));
 sky130_fd_sc_hd__sdfxtp_1 c723 (.CLK(clknet_4_14_0_clk),
    .D(net825),
    .SCD(clknet_1_0__leaf_net705),
    .SCE(net824),
    .Q(net706));
 sky130_fd_sc_hd__mux4_1 c724 (.A0(clknet_1_1__leaf_net698),
    .A1(net704),
    .A2(net701),
    .A3(net696),
    .S0(net706),
    .S1(clknet_1_1__leaf_net681),
    .X(net707));
 sky130_fd_sc_hd__dfbbn_1 c725 (.CLK_N(clknet_4_14_0_clk),
    .D(net700),
    .RESET_B(clknet_1_0__leaf_net705),
    .SET_B(clknet_1_1__leaf_net756),
    .Q(net709),
    .Q_N(net708));
 sky130_fd_sc_hd__a21bo_1 c726 (.A1(net706),
    .A2(net701),
    .B1_N(net703),
    .X(net710));
 sky130_fd_sc_hd__a21bo_1 c727 (.A1(net829),
    .A2(net710),
    .B1_N(net729),
    .X(net711));
 sky130_fd_sc_hd__dfbbn_1 c728 (.CLK_N(clknet_4_14_0_clk),
    .D(clknet_1_1__leaf_net705),
    .RESET_B(net710),
    .SET_B(net711),
    .Q(net713),
    .Q_N(net712));
 sky130_fd_sc_hd__a21bo_1 c729 (.A1(net710),
    .A2(net711),
    .B1_N(net713),
    .X(net714));
 sky130_fd_sc_hd__dfrbp_1 c73 (.CLK(clknet_4_4_0_clk),
    .D(net39),
    .RESET_B(net44),
    .Q(net51),
    .Q_N(net50));
 sky130_fd_sc_hd__mux4_1 c730 (.A0(net701),
    .A1(net713),
    .A2(net708),
    .A3(clknet_1_1__leaf_net756),
    .S0(clknet_1_1__leaf_net705),
    .S1(net714),
    .X(net715));
 sky130_fd_sc_hd__mux4_1 c731 (.A0(net714),
    .A1(net711),
    .A2(net712),
    .A3(net706),
    .S0(clknet_1_1__leaf_net756),
    .S1(net730));
 sky130_fd_sc_hd__dfrtn_1 c74 (.CLK_N(clknet_4_4_0_clk),
    .D(net43),
    .RESET_B(net39),
    .Q(net52));
 sky130_fd_sc_hd__xnor2_1 c75 (.A(net52),
    .B(net48),
    .Y(net53));
 sky130_fd_sc_hd__a31o_1 c76 (.A1(net41),
    .A2(net52),
    .A3(net795),
    .B1(net42),
    .X(net54));
 sky130_fd_sc_hd__dfrtp_1 c77 (.CLK(clknet_4_4_0_clk),
    .D(net53),
    .RESET_B(net54),
    .Q(net55));
 sky130_fd_sc_hd__dfbbn_1 c78 (.CLK_N(clknet_4_5_0_clk),
    .D(net54),
    .RESET_B(net44),
    .SET_B(net45),
    .Q(net57),
    .Q_N(net56));
 sky130_fd_sc_hd__dfrtp_1 c79 (.CLK(clknet_4_5_0_clk),
    .D(net44),
    .RESET_B(net56),
    .Q(net58));
 sky130_fd_sc_hd__a21bo_1 c80 (.A1(net46),
    .A2(net58),
    .B1_N(net42),
    .X(net59));
 sky130_fd_sc_hd__dfbbp_1 c81 (.CLK(clknet_4_4_0_clk),
    .D(net800),
    .RESET_B(net49),
    .SET_B(net47),
    .Q(net61),
    .Q_N(net60));
 sky130_fd_sc_hd__mux4_1 c82 (.A0(net38),
    .A1(net58),
    .A2(net53),
    .A3(net60),
    .S0(net42),
    .S1(net26),
    .X(net62));
 sky130_fd_sc_hd__mux4_1 c83 (.A0(net55),
    .A1(net59),
    .A2(net61),
    .A3(net62),
    .S0(net42),
    .S1(net54),
    .X(net63));
 sky130_fd_sc_hd__buf_1 c84 (.A(clknet_1_0__leaf_net716),
    .X(net64));
 sky130_fd_sc_hd__buf_1 c85 (.A(clknet_1_0__leaf_net64),
    .X(net65));
 sky130_fd_sc_hd__buf_1 c86 (.A(clknet_1_0__leaf_net65),
    .X(net66));
 sky130_fd_sc_hd__buf_1 c87 (.A(clknet_1_1__leaf_net65),
    .X(net67));
 sky130_fd_sc_hd__xnor2_1 c88 (.A(clknet_1_0__leaf_net67),
    .B(clknet_1_0__leaf_net64),
    .Y(net68));
 sky130_fd_sc_hd__buf_1 c89 (.A(clknet_1_1__leaf_net66),
    .X(net69));
 sky130_fd_sc_hd__xnor2_1 c90 (.A(clknet_1_1__leaf_net65),
    .B(clknet_1_0__leaf_net69),
    .Y(net70));
 sky130_fd_sc_hd__xnor2_1 c91 (.A(clknet_1_0__leaf_net65),
    .B(clknet_1_0__leaf_net69),
    .Y(net71));
 sky130_fd_sc_hd__xnor2_1 c92 (.A(clknet_1_1__leaf_net68),
    .B(clknet_1_1__leaf_net69),
    .Y(net72));
 sky130_fd_sc_hd__a31o_1 c93 (.A1(clknet_1_0__leaf_net70),
    .A2(clknet_1_0__leaf_net68),
    .A3(clknet_1_0__leaf_net71),
    .B1(clknet_1_0__leaf_net69),
    .X(net73));
 sky130_fd_sc_hd__xnor2_1 c94 (.A(clknet_1_0__leaf_net66),
    .B(clknet_1_0__leaf_net71),
    .Y(net74));
 sky130_fd_sc_hd__xnor2_1 c95 (.A(net74),
    .B(clknet_1_1__leaf_net68),
    .Y(net75));
 sky130_fd_sc_hd__xnor2_1 c96 (.A(clknet_1_1__leaf_net71),
    .B(clknet_1_0__leaf_net72),
    .Y(net76));
 sky130_fd_sc_hd__a21bo_1 c97 (.A1(clknet_1_0__leaf_net69),
    .A2(clknet_1_1__leaf_net67),
    .B1_N(clknet_1_0__leaf_net71),
    .X(net77));
 sky130_fd_sc_hd__a21bo_1 c98 (.A1(clknet_1_0__leaf_net77),
    .A2(clknet_1_0__leaf_net76),
    .B1_N(clknet_1_1__leaf_net71),
    .X(net78));
 sky130_fd_sc_hd__a21bo_1 c99 (.A1(net73),
    .A2(clknet_1_0__leaf_net69),
    .B1_N(clknet_1_0__leaf_net68),
    .X(net79));
 sky130_fd_sc_hd__dlclkp_4 s732 (.CLK(clknet_4_5_0_clk),
    .GATE(net63),
    .GCLK(net716));
 sky130_fd_sc_hd__dlxbn_1 s733 (.D(net169),
    .GATE_N(clknet_4_4_0_clk),
    .Q(net717));
 sky130_fd_sc_hd__dlxbn_1 s734 (.D(net259),
    .GATE_N(clknet_4_0_0_clk),
    .Q(net718));
 sky130_fd_sc_hd__dlxbp_1 s735 (.D(net281),
    .GATE(clknet_4_1_0_clk),
    .Q(net720),
    .Q_N(net719));
 sky130_fd_sc_hd__dlxtn_1 s736 (.D(net326),
    .GATE_N(clknet_4_6_0_clk),
    .Q(net721));
 sky130_fd_sc_hd__dlxtn_1 s737 (.D(net327),
    .GATE_N(clknet_4_6_0_clk),
    .Q(net722));
 sky130_fd_sc_hd__dlxtn_1 s738 (.D(net370),
    .GATE_N(clknet_4_13_0_clk),
    .Q(net723));
 sky130_fd_sc_hd__dlxtp_1 s739 (.D(net420),
    .GATE(clknet_4_3_0_clk),
    .Q(net724));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s740 (.D(net459),
    .SLEEP_B(clknet_4_12_0_clk),
    .Q(net725));
 sky130_fd_sc_hd__dfxbp_1 s741 (.CLK(clknet_4_9_0_clk),
    .D(net547),
    .Q(net726));
 sky130_fd_sc_hd__dfxbp_1 s742 (.CLK(clknet_4_10_0_clk),
    .D(net685),
    .Q(net727));
 sky130_fd_sc_hd__dfxtp_1 s743 (.CLK(clknet_4_10_0_clk),
    .D(net693),
    .Q(net728));
 sky130_fd_sc_hd__dfxtp_1 s744 (.CLK(clknet_4_11_0_clk),
    .D(net707),
    .Q(net729));
 sky130_fd_sc_hd__dfxtp_1 s745 (.CLK(clknet_4_14_0_clk),
    .D(net715),
    .Q(net730));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Right_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Right_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Right_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Right_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Right_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Right_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Right_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Right_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Right_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Right_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Right_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Right_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Right_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Right_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Right_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Right_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Right_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Right_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Right_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Right_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Right_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_161 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_162 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_163 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_164 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_165 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_166 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_167 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_168 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_169 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_170 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_171 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_172 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_173 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_174 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_175 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_176 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_177 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_178 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_179 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_180 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_181 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_182 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Left_183 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Left_184 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Left_185 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Left_186 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Left_187 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Left_188 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Left_189 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Left_190 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Left_191 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Left_192 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Left_193 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Left_194 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Left_195 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Left_196 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Left_197 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Left_198 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Left_199 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Left_200 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Left_201 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Left_202 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Left_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1347 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(in0),
    .X(net731));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(in1),
    .X(net732));
 sky130_fd_sc_hd__buf_1 input3 (.A(in10),
    .X(net733));
 sky130_fd_sc_hd__clkbuf_2 input4 (.A(in11),
    .X(net734));
 sky130_fd_sc_hd__clkbuf_2 input5 (.A(in12),
    .X(net735));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(in13),
    .X(net736));
 sky130_fd_sc_hd__clkbuf_2 input7 (.A(in15),
    .X(net737));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(in16),
    .X(net738));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(in17),
    .X(net739));
 sky130_fd_sc_hd__clkbuf_2 input10 (.A(in18),
    .X(net740));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(in19),
    .X(net741));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(in2),
    .X(net742));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(in20),
    .X(net743));
 sky130_fd_sc_hd__buf_2 input14 (.A(in21),
    .X(net744));
 sky130_fd_sc_hd__buf_2 input15 (.A(in22),
    .X(net745));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(in23),
    .X(net746));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(in24),
    .X(net747));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(in3),
    .X(net748));
 sky130_fd_sc_hd__clkbuf_1 input19 (.A(in4),
    .X(net749));
 sky130_fd_sc_hd__clkbuf_1 input20 (.A(in5),
    .X(net750));
 sky130_fd_sc_hd__clkbuf_1 input21 (.A(in6),
    .X(net751));
 sky130_fd_sc_hd__clkbuf_1 input22 (.A(in7),
    .X(net752));
 sky130_fd_sc_hd__clkbuf_1 input23 (.A(in8),
    .X(net753));
 sky130_fd_sc_hd__clkbuf_1 input24 (.A(in9),
    .X(net754));
 sky130_fd_sc_hd__buf_2 output25 (.A(net755),
    .X(out1));
 sky130_fd_sc_hd__clkbuf_1 output26 (.A(clknet_1_1__leaf_net756),
    .X(out10));
 sky130_fd_sc_hd__clkbuf_1 output27 (.A(clknet_1_1__leaf_net757),
    .X(out11));
 sky130_fd_sc_hd__buf_2 output28 (.A(net758),
    .X(out16));
 sky130_fd_sc_hd__buf_2 output29 (.A(net759),
    .X(out17));
 sky130_fd_sc_hd__clkbuf_4 output30 (.A(net760),
    .X(out18));
 sky130_fd_sc_hd__clkbuf_1 output31 (.A(clknet_1_1__leaf_net761),
    .X(out19));
 sky130_fd_sc_hd__buf_2 output32 (.A(net762),
    .X(out2));
 sky130_fd_sc_hd__buf_2 output33 (.A(net763),
    .X(out20));
 sky130_fd_sc_hd__buf_2 output34 (.A(net764),
    .X(out21));
 sky130_fd_sc_hd__buf_2 output35 (.A(net765),
    .X(out22));
 sky130_fd_sc_hd__buf_2 output36 (.A(net766),
    .X(out23));
 sky130_fd_sc_hd__buf_2 output37 (.A(net767),
    .X(out24));
 sky130_fd_sc_hd__buf_2 output38 (.A(net768),
    .X(out4));
 sky130_fd_sc_hd__clkbuf_1 output39 (.A(net769),
    .X(out6));
 sky130_fd_sc_hd__clkbuf_1 output40 (.A(net770),
    .X(out8));
 sky130_fd_sc_hd__buf_4 max_cap41 (.A(net525),
    .X(net771));
 sky130_fd_sc_hd__buf_4 max_cap42 (.A(net496),
    .X(net772));
 sky130_fd_sc_hd__buf_4 max_cap43 (.A(net137),
    .X(net773));
 sky130_fd_sc_hd__buf_4 wire44 (.A(net494),
    .X(net774));
 sky130_fd_sc_hd__buf_4 max_cap45 (.A(net239),
    .X(net775));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net716 (.A(net716),
    .X(clknet_0_net716));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net716 (.A(clknet_0_net716),
    .X(clknet_1_0__leaf_net716));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net716 (.A(clknet_0_net716),
    .X(clknet_1_1__leaf_net716));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net64 (.A(net64),
    .X(clknet_0_net64));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net64 (.A(clknet_0_net64),
    .X(clknet_1_0__leaf_net64));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net64 (.A(clknet_0_net64),
    .X(clknet_1_1__leaf_net64));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net68 (.A(net68),
    .X(clknet_0_net68));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net68 (.A(clknet_0_net68),
    .X(clknet_1_0__leaf_net68));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net68 (.A(clknet_0_net68),
    .X(clknet_1_1__leaf_net68));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net79 (.A(net79),
    .X(clknet_0_net79));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net79 (.A(clknet_0_net79),
    .X(clknet_1_0__leaf_net79));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net79 (.A(clknet_0_net79),
    .X(clknet_1_1__leaf_net79));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net82 (.A(net82),
    .X(clknet_0_net82));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net82 (.A(clknet_0_net82),
    .X(clknet_1_0__leaf_net82));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net82 (.A(clknet_0_net82),
    .X(clknet_1_1__leaf_net82));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net84 (.A(net84),
    .X(clknet_0_net84));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net84 (.A(clknet_0_net84),
    .X(clknet_1_0__leaf_net84));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net84 (.A(clknet_0_net84),
    .X(clknet_1_1__leaf_net84));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net219 (.A(net219),
    .X(clknet_0_net219));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net219 (.A(clknet_0_net219),
    .X(clknet_1_0__leaf_net219));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net219 (.A(clknet_0_net219),
    .X(clknet_1_1__leaf_net219));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net85 (.A(net85),
    .X(clknet_0_net85));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net85 (.A(clknet_0_net85),
    .X(clknet_1_0__leaf_net85));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net85 (.A(clknet_0_net85),
    .X(clknet_1_1__leaf_net85));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net92 (.A(net92),
    .X(clknet_0_net92));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net92 (.A(clknet_0_net92),
    .X(clknet_1_0__leaf_net92));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net92 (.A(clknet_0_net92),
    .X(clknet_1_1__leaf_net92));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net102 (.A(net102),
    .X(clknet_0_net102));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net102 (.A(clknet_0_net102),
    .X(clknet_1_0__leaf_net102));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net102 (.A(clknet_0_net102),
    .X(clknet_1_1__leaf_net102));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net87 (.A(net87),
    .X(clknet_0_net87));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net87 (.A(clknet_0_net87),
    .X(clknet_1_0__leaf_net87));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net87 (.A(clknet_0_net87),
    .X(clknet_1_1__leaf_net87));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net91 (.A(net91),
    .X(clknet_0_net91));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net91 (.A(clknet_0_net91),
    .X(clknet_1_0__leaf_net91));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net91 (.A(clknet_0_net91),
    .X(clknet_1_1__leaf_net91));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net90 (.A(net90),
    .X(clknet_0_net90));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net90 (.A(clknet_0_net90),
    .X(clknet_1_0__leaf_net90));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net90 (.A(clknet_0_net90),
    .X(clknet_1_1__leaf_net90));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net89 (.A(net89),
    .X(clknet_0_net89));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net89 (.A(clknet_0_net89),
    .X(clknet_1_0__leaf_net89));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net89 (.A(clknet_0_net89),
    .X(clknet_1_1__leaf_net89));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net88 (.A(net88),
    .X(clknet_0_net88));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net88 (.A(clknet_0_net88),
    .X(clknet_1_0__leaf_net88));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net88 (.A(clknet_0_net88),
    .X(clknet_1_1__leaf_net88));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net72 (.A(net72),
    .X(clknet_0_net72));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net72 (.A(clknet_0_net72),
    .X(clknet_1_0__leaf_net72));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net72 (.A(clknet_0_net72),
    .X(clknet_1_1__leaf_net72));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net76 (.A(net76),
    .X(clknet_0_net76));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net76 (.A(clknet_0_net76),
    .X(clknet_1_0__leaf_net76));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net76 (.A(clknet_0_net76),
    .X(clknet_1_1__leaf_net76));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net78 (.A(net78),
    .X(clknet_0_net78));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net78 (.A(clknet_0_net78),
    .X(clknet_1_0__leaf_net78));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net78 (.A(clknet_0_net78),
    .X(clknet_1_1__leaf_net78));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net336 (.A(net336),
    .X(clknet_0_net336));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net336 (.A(clknet_0_net336),
    .X(clknet_1_0__leaf_net336));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net336 (.A(clknet_0_net336),
    .X(clknet_1_1__leaf_net336));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net337 (.A(net337),
    .X(clknet_0_net337));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net337 (.A(clknet_0_net337),
    .X(clknet_1_0__leaf_net337));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net337 (.A(clknet_0_net337),
    .X(clknet_1_1__leaf_net337));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net355 (.A(net355),
    .X(clknet_0_net355));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net355 (.A(clknet_0_net355),
    .X(clknet_1_0__leaf_net355));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net355 (.A(clknet_0_net355),
    .X(clknet_1_1__leaf_net355));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net361 (.A(net361),
    .X(clknet_0_net361));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net361 (.A(clknet_0_net361),
    .X(clknet_1_0__leaf_net361));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net361 (.A(clknet_0_net361),
    .X(clknet_1_1__leaf_net361));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net356 (.A(net356),
    .X(clknet_0_net356));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net356 (.A(clknet_0_net356),
    .X(clknet_1_0__leaf_net356));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net356 (.A(clknet_0_net356),
    .X(clknet_1_1__leaf_net356));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net340 (.A(net340),
    .X(clknet_0_net340));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net340 (.A(clknet_0_net340),
    .X(clknet_1_0__leaf_net340));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net340 (.A(clknet_0_net340),
    .X(clknet_1_1__leaf_net340));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net341 (.A(net341),
    .X(clknet_0_net341));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net341 (.A(clknet_0_net341),
    .X(clknet_1_0__leaf_net341));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net341 (.A(clknet_0_net341),
    .X(clknet_1_1__leaf_net341));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net215 (.A(net215),
    .X(clknet_0_net215));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net215 (.A(clknet_0_net215),
    .X(clknet_1_0__leaf_net215));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net215 (.A(clknet_0_net215),
    .X(clknet_1_1__leaf_net215));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net210 (.A(net210),
    .X(clknet_0_net210));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net210 (.A(clknet_0_net210),
    .X(clknet_1_0__leaf_net210));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net210 (.A(clknet_0_net210),
    .X(clknet_1_1__leaf_net210));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net216 (.A(net216),
    .X(clknet_0_net216));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net216 (.A(clknet_0_net216),
    .X(clknet_1_0__leaf_net216));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net216 (.A(clknet_0_net216),
    .X(clknet_1_1__leaf_net216));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net223 (.A(net223),
    .X(clknet_0_net223));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net223 (.A(clknet_0_net223),
    .X(clknet_1_0__leaf_net223));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net223 (.A(clknet_0_net223),
    .X(clknet_1_1__leaf_net223));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net218 (.A(net218),
    .X(clknet_0_net218));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net218 (.A(clknet_0_net218),
    .X(clknet_1_0__leaf_net218));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net218 (.A(clknet_0_net218),
    .X(clknet_1_1__leaf_net218));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net211 (.A(net211),
    .X(clknet_0_net211));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net211 (.A(clknet_0_net211),
    .X(clknet_1_0__leaf_net211));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net211 (.A(clknet_0_net211),
    .X(clknet_1_1__leaf_net211));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net195 (.A(net195),
    .X(clknet_0_net195));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net195 (.A(clknet_0_net195),
    .X(clknet_1_0__leaf_net195));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net195 (.A(clknet_0_net195),
    .X(clknet_1_1__leaf_net195));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net198 (.A(net198),
    .X(clknet_0_net198));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net198 (.A(clknet_0_net198),
    .X(clknet_1_0__leaf_net198));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net198 (.A(net784),
    .X(clknet_1_1__leaf_net198));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net202 (.A(net202),
    .X(clknet_0_net202));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net202 (.A(clknet_0_net202),
    .X(clknet_1_0__leaf_net202));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net202 (.A(clknet_0_net202),
    .X(clknet_1_1__leaf_net202));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net206 (.A(net206),
    .X(clknet_0_net206));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net206 (.A(clknet_0_net206),
    .X(clknet_1_0__leaf_net206));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net206 (.A(clknet_0_net206),
    .X(clknet_1_1__leaf_net206));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net205 (.A(net205),
    .X(clknet_0_net205));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net205 (.A(clknet_0_net205),
    .X(clknet_1_0__leaf_net205));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net205 (.A(clknet_0_net205),
    .X(clknet_1_1__leaf_net205));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net207 (.A(net207),
    .X(clknet_0_net207));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net207 (.A(clknet_0_net207),
    .X(clknet_1_0__leaf_net207));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net207 (.A(clknet_0_net207),
    .X(clknet_1_1__leaf_net207));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net200 (.A(net200),
    .X(clknet_0_net200));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net200 (.A(clknet_0_net200),
    .X(clknet_1_0__leaf_net200));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net200 (.A(clknet_0_net200),
    .X(clknet_1_1__leaf_net200));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net196 (.A(net196),
    .X(clknet_0_net196));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net196 (.A(clknet_0_net196),
    .X(clknet_1_0__leaf_net196));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net196 (.A(net783),
    .X(clknet_1_1__leaf_net196));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net65 (.A(net65),
    .X(clknet_0_net65));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net65 (.A(clknet_0_net65),
    .X(clknet_1_0__leaf_net65));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net65 (.A(clknet_0_net65),
    .X(clknet_1_1__leaf_net65));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net71 (.A(net71),
    .X(clknet_0_net71));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net71 (.A(clknet_0_net71),
    .X(clknet_1_0__leaf_net71));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net71 (.A(clknet_0_net71),
    .X(clknet_1_1__leaf_net71));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net77 (.A(net77),
    .X(clknet_0_net77));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net77 (.A(clknet_0_net77),
    .X(clknet_1_0__leaf_net77));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net77 (.A(clknet_0_net77),
    .X(clknet_1_1__leaf_net77));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net70 (.A(net70),
    .X(clknet_0_net70));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net70 (.A(clknet_0_net70),
    .X(clknet_1_0__leaf_net70));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net70 (.A(clknet_0_net70),
    .X(clknet_1_1__leaf_net70));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net67 (.A(net67),
    .X(clknet_0_net67));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net67 (.A(clknet_0_net67),
    .X(clknet_1_0__leaf_net67));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net67 (.A(clknet_0_net67),
    .X(clknet_1_1__leaf_net67));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net66 (.A(net66),
    .X(clknet_0_net66));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net66 (.A(clknet_0_net66),
    .X(clknet_1_0__leaf_net66));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net66 (.A(clknet_0_net66),
    .X(clknet_1_1__leaf_net66));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net69 (.A(net69),
    .X(clknet_0_net69));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net69 (.A(clknet_0_net69),
    .X(clknet_1_0__leaf_net69));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net69 (.A(clknet_0_net69),
    .X(clknet_1_1__leaf_net69));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net192 (.A(net192),
    .X(clknet_0_net192));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net192 (.A(clknet_0_net192),
    .X(clknet_1_0__leaf_net192));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net192 (.A(clknet_0_net192),
    .X(clknet_1_1__leaf_net192));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net650 (.A(net650),
    .X(clknet_0_net650));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net650 (.A(clknet_0_net650),
    .X(clknet_1_0__leaf_net650));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net650 (.A(clknet_0_net650),
    .X(clknet_1_1__leaf_net650));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net652 (.A(net652),
    .X(clknet_0_net652));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net652 (.A(clknet_0_net652),
    .X(clknet_1_0__leaf_net652));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net652 (.A(clknet_0_net652),
    .X(clknet_1_1__leaf_net652));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net680 (.A(net680),
    .X(clknet_0_net680));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net680 (.A(clknet_0_net680),
    .X(clknet_1_0__leaf_net680));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net680 (.A(clknet_0_net680),
    .X(clknet_1_1__leaf_net680));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net681 (.A(net681),
    .X(clknet_0_net681));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net681 (.A(clknet_0_net681),
    .X(clknet_1_0__leaf_net681));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net681 (.A(clknet_0_net681),
    .X(clknet_1_1__leaf_net681));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net664 (.A(net664),
    .X(clknet_0_net664));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net664 (.A(clknet_0_net664),
    .X(clknet_1_0__leaf_net664));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net664 (.A(clknet_0_net664),
    .X(clknet_1_1__leaf_net664));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net672 (.A(net672),
    .X(clknet_0_net672));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net672 (.A(clknet_0_net672),
    .X(clknet_1_0__leaf_net672));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net672 (.A(clknet_0_net672),
    .X(clknet_1_1__leaf_net672));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net673 (.A(net673),
    .X(clknet_0_net673));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net673 (.A(clknet_0_net673),
    .X(clknet_1_0__leaf_net673));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net673 (.A(clknet_0_net673),
    .X(clknet_1_1__leaf_net673));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net698 (.A(net698),
    .X(clknet_0_net698));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net698 (.A(clknet_0_net698),
    .X(clknet_1_0__leaf_net698));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net698 (.A(clknet_0_net698),
    .X(clknet_1_1__leaf_net698));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net692 (.A(net692),
    .X(clknet_0_net692));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net692 (.A(clknet_0_net692),
    .X(clknet_1_0__leaf_net692));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net692 (.A(clknet_0_net692),
    .X(clknet_1_1__leaf_net692));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net677 (.A(net677),
    .X(clknet_0_net677));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net677 (.A(clknet_0_net677),
    .X(clknet_1_0__leaf_net677));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net677 (.A(clknet_0_net677),
    .X(clknet_1_1__leaf_net677));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net659 (.A(net659),
    .X(clknet_0_net659));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net659 (.A(clknet_0_net659),
    .X(clknet_1_0__leaf_net659));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net659 (.A(clknet_0_net659),
    .X(clknet_1_1__leaf_net659));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net662 (.A(net662),
    .X(clknet_0_net662));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net662 (.A(clknet_0_net662),
    .X(clknet_1_0__leaf_net662));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net662 (.A(clknet_0_net662),
    .X(clknet_1_1__leaf_net662));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net663 (.A(net663),
    .X(clknet_0_net663));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net663 (.A(clknet_0_net663),
    .X(clknet_1_0__leaf_net663));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net663 (.A(clknet_0_net663),
    .X(clknet_1_1__leaf_net663));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net655 (.A(net655),
    .X(clknet_0_net655));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net655 (.A(clknet_0_net655),
    .X(clknet_1_0__leaf_net655));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net655 (.A(clknet_0_net655),
    .X(clknet_1_1__leaf_net655));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net654 (.A(net654),
    .X(clknet_0_net654));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net654 (.A(clknet_0_net654),
    .X(clknet_1_0__leaf_net654));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net654 (.A(clknet_0_net654),
    .X(clknet_1_1__leaf_net654));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net656 (.A(net656),
    .X(clknet_0_net656));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net656 (.A(clknet_0_net656),
    .X(clknet_1_0__leaf_net656));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net656 (.A(clknet_0_net656),
    .X(clknet_1_1__leaf_net656));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net668 (.A(net668),
    .X(clknet_0_net668));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net668 (.A(clknet_0_net668),
    .X(clknet_1_0__leaf_net668));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net668 (.A(clknet_0_net668),
    .X(clknet_1_1__leaf_net668));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net676 (.A(net676),
    .X(clknet_0_net676));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net676 (.A(clknet_0_net676),
    .X(clknet_1_0__leaf_net676));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net676 (.A(clknet_0_net676),
    .X(clknet_1_1__leaf_net676));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net653 (.A(net653),
    .X(clknet_0_net653));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net653 (.A(clknet_0_net653),
    .X(clknet_1_0__leaf_net653));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net653 (.A(clknet_0_net653),
    .X(clknet_1_1__leaf_net653));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net660 (.A(net660),
    .X(clknet_0_net660));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net660 (.A(clknet_0_net660),
    .X(clknet_1_0__leaf_net660));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net660 (.A(clknet_0_net660),
    .X(clknet_1_1__leaf_net660));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net651 (.A(net651),
    .X(clknet_0_net651));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net651 (.A(clknet_0_net651),
    .X(clknet_1_0__leaf_net651));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net651 (.A(clknet_0_net651),
    .X(clknet_1_1__leaf_net651));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net647 (.A(net647),
    .X(clknet_0_net647));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net647 (.A(clknet_0_net647),
    .X(clknet_1_0__leaf_net647));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net647 (.A(clknet_0_net647),
    .X(clknet_1_1__leaf_net647));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net648 (.A(net648),
    .X(clknet_0_net648));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net648 (.A(clknet_0_net648),
    .X(clknet_1_0__leaf_net648));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net648 (.A(clknet_0_net648),
    .X(clknet_1_1__leaf_net648));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net559 (.A(net559),
    .X(clknet_0_net559));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net559 (.A(clknet_0_net559),
    .X(clknet_1_0__leaf_net559));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net559 (.A(clknet_0_net559),
    .X(clknet_1_1__leaf_net559));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net573 (.A(net573),
    .X(clknet_0_net573));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net573 (.A(clknet_0_net573),
    .X(clknet_1_0__leaf_net573));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net573 (.A(clknet_0_net573),
    .X(clknet_1_1__leaf_net573));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net669 (.A(net669),
    .X(clknet_0_net669));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net669 (.A(clknet_0_net669),
    .X(clknet_1_0__leaf_net669));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net669 (.A(clknet_0_net669),
    .X(clknet_1_1__leaf_net669));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net581 (.A(net581),
    .X(clknet_0_net581));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net581 (.A(clknet_0_net581),
    .X(clknet_1_0__leaf_net581));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net581 (.A(clknet_0_net581),
    .X(clknet_1_1__leaf_net581));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net582 (.A(net582),
    .X(clknet_0_net582));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net582 (.A(clknet_0_net582),
    .X(clknet_1_0__leaf_net582));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net582 (.A(clknet_0_net582),
    .X(clknet_1_1__leaf_net582));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net756 (.A(net756),
    .X(clknet_0_net756));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net756 (.A(clknet_0_net756),
    .X(clknet_1_0__leaf_net756));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net756 (.A(clknet_0_net756),
    .X(clknet_1_1__leaf_net756));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net705 (.A(net705),
    .X(clknet_0_net705));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net705 (.A(clknet_0_net705),
    .X(clknet_1_0__leaf_net705));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net705 (.A(clknet_0_net705),
    .X(clknet_1_1__leaf_net705));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net757 (.A(net757),
    .X(clknet_0_net757));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net757 (.A(clknet_0_net757),
    .X(clknet_1_0__leaf_net757));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net757 (.A(clknet_0_net757),
    .X(clknet_1_1__leaf_net757));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net585 (.A(net585),
    .X(clknet_0_net585));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net585 (.A(clknet_0_net585),
    .X(clknet_1_0__leaf_net585));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net585 (.A(clknet_0_net585),
    .X(clknet_1_1__leaf_net585));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net578 (.A(net578),
    .X(clknet_0_net578));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net578 (.A(clknet_0_net578),
    .X(clknet_1_0__leaf_net578));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net578 (.A(clknet_0_net578),
    .X(clknet_1_1__leaf_net578));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net580 (.A(net580),
    .X(clknet_0_net580));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net580 (.A(clknet_0_net580),
    .X(clknet_1_0__leaf_net580));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net580 (.A(clknet_0_net580),
    .X(clknet_1_1__leaf_net580));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net584 (.A(net584),
    .X(clknet_0_net584));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net584 (.A(clknet_0_net584),
    .X(clknet_1_0__leaf_net584));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net584 (.A(clknet_0_net584),
    .X(clknet_1_1__leaf_net584));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net761 (.A(net761),
    .X(clknet_0_net761));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net761 (.A(clknet_0_net761),
    .X(clknet_1_0__leaf_net761));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net761 (.A(clknet_0_net761),
    .X(clknet_1_1__leaf_net761));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net564 (.A(net564),
    .X(clknet_0_net564));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net564 (.A(clknet_0_net564),
    .X(clknet_1_0__leaf_net564));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net564 (.A(clknet_0_net564),
    .X(clknet_1_1__leaf_net564));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net565 (.A(net565),
    .X(clknet_0_net565));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net565 (.A(clknet_0_net565),
    .X(clknet_1_0__leaf_net565));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net565 (.A(clknet_0_net565),
    .X(clknet_1_1__leaf_net565));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net558 (.A(net558),
    .X(clknet_0_net558));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net558 (.A(clknet_0_net558),
    .X(clknet_1_0__leaf_net558));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net558 (.A(clknet_0_net558),
    .X(clknet_1_1__leaf_net558));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net562 (.A(net562),
    .X(clknet_0_net562));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net562 (.A(clknet_0_net562),
    .X(clknet_1_0__leaf_net562));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net562 (.A(clknet_0_net562),
    .X(clknet_1_1__leaf_net562));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net280 (.A(net280),
    .X(clknet_0_net280));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net280 (.A(clknet_0_net280),
    .X(clknet_1_0__leaf_net280));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net280 (.A(clknet_0_net280),
    .X(clknet_1_1__leaf_net280));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net398 (.A(net398),
    .X(clknet_0_net398));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net398 (.A(clknet_0_net398),
    .X(clknet_1_0__leaf_net398));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net398 (.A(clknet_0_net398),
    .X(clknet_1_1__leaf_net398));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net404 (.A(net404),
    .X(clknet_0_net404));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net404 (.A(clknet_0_net404),
    .X(clknet_1_0__leaf_net404));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net404 (.A(clknet_0_net404),
    .X(clknet_1_1__leaf_net404));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net408 (.A(net408),
    .X(clknet_0_net408));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net408 (.A(clknet_0_net408),
    .X(clknet_1_0__leaf_net408));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net408 (.A(clknet_0_net408),
    .X(clknet_1_1__leaf_net408));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net413 (.A(net413),
    .X(clknet_0_net413));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net413 (.A(clknet_0_net413),
    .X(clknet_1_0__leaf_net413));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net413 (.A(clknet_0_net413),
    .X(clknet_1_1__leaf_net413));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net411 (.A(net411),
    .X(clknet_0_net411));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net411 (.A(clknet_0_net411),
    .X(clknet_1_0__leaf_net411));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net411 (.A(clknet_0_net411),
    .X(clknet_1_1__leaf_net411));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net409 (.A(net409),
    .X(clknet_0_net409));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net409 (.A(clknet_0_net409),
    .X(clknet_1_0__leaf_net409));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net409 (.A(clknet_0_net409),
    .X(clknet_1_1__leaf_net409));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net530 (.A(net530),
    .X(clknet_0_net530));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net530 (.A(clknet_0_net530),
    .X(clknet_1_0__leaf_net530));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net530 (.A(clknet_0_net530),
    .X(clknet_1_1__leaf_net530));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net426 (.A(net426),
    .X(clknet_0_net426));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net426 (.A(clknet_0_net426),
    .X(clknet_1_0__leaf_net426));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net426 (.A(clknet_0_net426),
    .X(clknet_1_1__leaf_net426));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net441 (.A(net441),
    .X(clknet_0_net441));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net441 (.A(clknet_0_net441),
    .X(clknet_1_0__leaf_net441));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net441 (.A(clknet_0_net441),
    .X(clknet_1_1__leaf_net441));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net410 (.A(net410),
    .X(clknet_0_net410));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net410 (.A(clknet_0_net410),
    .X(clknet_1_0__leaf_net410));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net410 (.A(clknet_0_net410),
    .X(clknet_1_1__leaf_net410));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net407 (.A(net407),
    .X(clknet_0_net407));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net407 (.A(clknet_0_net407),
    .X(clknet_1_0__leaf_net407));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net407 (.A(clknet_0_net407),
    .X(clknet_1_1__leaf_net407));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net401 (.A(net401),
    .X(clknet_0_net401));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net401 (.A(clknet_0_net401),
    .X(clknet_1_0__leaf_net401));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net401 (.A(clknet_0_net401),
    .X(clknet_1_1__leaf_net401));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net402 (.A(net402),
    .X(clknet_0_net402));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net402 (.A(clknet_0_net402),
    .X(clknet_1_0__leaf_net402));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net402 (.A(clknet_0_net402),
    .X(clknet_1_1__leaf_net402));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net406 (.A(net406),
    .X(clknet_0_net406));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net406 (.A(clknet_0_net406),
    .X(clknet_1_0__leaf_net406));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net406 (.A(clknet_0_net406),
    .X(clknet_1_1__leaf_net406));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net405 (.A(net405),
    .X(clknet_0_net405));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net405 (.A(clknet_0_net405),
    .X(clknet_1_0__leaf_net405));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net405 (.A(clknet_0_net405),
    .X(clknet_1_1__leaf_net405));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net403 (.A(net403),
    .X(clknet_0_net403));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net403 (.A(clknet_0_net403),
    .X(clknet_1_0__leaf_net403));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net403 (.A(clknet_0_net403),
    .X(clknet_1_1__leaf_net403));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net437 (.A(net437),
    .X(clknet_0_net437));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net437 (.A(clknet_0_net437),
    .X(clknet_1_0__leaf_net437));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net437 (.A(clknet_0_net437),
    .X(clknet_1_1__leaf_net437));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net439 (.A(net439),
    .X(clknet_0_net439));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net439 (.A(clknet_0_net439),
    .X(clknet_1_0__leaf_net439));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net439 (.A(clknet_0_net439),
    .X(clknet_1_1__leaf_net439));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net571 (.A(net571),
    .X(clknet_0_net571));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net571 (.A(clknet_0_net571),
    .X(clknet_1_0__leaf_net571));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net571 (.A(clknet_0_net571),
    .X(clknet_1_1__leaf_net571));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net440 (.A(net440),
    .X(clknet_0_net440));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net440 (.A(clknet_0_net440),
    .X(clknet_1_0__leaf_net440));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net440 (.A(clknet_0_net440),
    .X(clknet_1_1__leaf_net440));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net270 (.A(net270),
    .X(clknet_0_net270));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net270 (.A(clknet_0_net270),
    .X(clknet_1_0__leaf_net270));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net270 (.A(clknet_0_net270),
    .X(clknet_1_1__leaf_net270));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net272 (.A(net272),
    .X(clknet_0_net272));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net272 (.A(clknet_0_net272),
    .X(clknet_1_0__leaf_net272));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net272 (.A(clknet_0_net272),
    .X(clknet_1_1__leaf_net272));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net275 (.A(net275),
    .X(clknet_0_net275));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net275 (.A(clknet_0_net275),
    .X(clknet_1_0__leaf_net275));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net275 (.A(clknet_0_net275),
    .X(clknet_1_1__leaf_net275));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net273 (.A(net273),
    .X(clknet_0_net273));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net273 (.A(clknet_0_net273),
    .X(clknet_1_0__leaf_net273));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net273 (.A(clknet_0_net273),
    .X(clknet_1_1__leaf_net273));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net285 (.A(net285),
    .X(clknet_0_net285));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net285 (.A(clknet_0_net285),
    .X(clknet_1_0__leaf_net285));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net285 (.A(clknet_0_net285),
    .X(clknet_1_1__leaf_net285));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net300 (.A(net300),
    .X(clknet_0_net300));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net300 (.A(clknet_0_net300),
    .X(clknet_1_0__leaf_net300));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net300 (.A(clknet_0_net300),
    .X(clknet_1_1__leaf_net300));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net287 (.A(net287),
    .X(clknet_0_net287));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net287 (.A(clknet_0_net287),
    .X(clknet_1_0__leaf_net287));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net287 (.A(clknet_0_net287),
    .X(clknet_1_1__leaf_net287));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer1 (.A(net181),
    .X(net776));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer2 (.A(net776),
    .X(net777));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer3 (.A(net777),
    .X(net778));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer4 (.A(net778),
    .X(net779));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer5 (.A(net187),
    .X(net780));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer6 (.A(net780),
    .X(net781));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer7 (.A(net180),
    .X(net782));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer8 (.A(clknet_0_net196),
    .X(net783));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer9 (.A(clknet_0_net198),
    .X(net784));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer10 (.A(clknet_1_0__leaf_net196),
    .X(net785));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(net286),
    .X(net786));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(net165),
    .X(net787));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(net295),
    .X(net788));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(net299),
    .X(net789));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(net303),
    .X(net790));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(net512),
    .X(net791));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(net508),
    .X(net792));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(net696),
    .X(net793));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(net95),
    .X(net794));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(net50),
    .X(net795));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(net549),
    .X(net796));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(net232),
    .X(net797));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(net617),
    .X(net798));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(net301),
    .X(net799));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(net51),
    .X(net800));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(net365),
    .X(net801));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(net599),
    .X(net802));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(net46),
    .X(net803));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(net625),
    .X(net804));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(net421),
    .X(net805));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(net728),
    .X(net806));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(net643),
    .X(net807));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(net630),
    .X(net808));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(net360),
    .X(net809));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(net637),
    .X(net810));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(net725),
    .X(net811));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(net98),
    .X(net812));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(net697),
    .X(net813));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(net594),
    .X(net814));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(net671),
    .X(net815));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(net570),
    .X(net816));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(net694),
    .X(net817));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(net278),
    .X(net818));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(net416),
    .X(net819));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(net587),
    .X(net820));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(net233),
    .X(net821));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(net362),
    .X(net822));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(net636),
    .X(net823));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(net700),
    .X(net824));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(net703),
    .X(net825));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(net566),
    .X(net826));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(net626),
    .X(net827));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(net357),
    .X(net828));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(net709),
    .X(net829));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(net646),
    .X(net830));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(net631),
    .X(net831));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(net760),
    .X(net832));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(net97),
    .X(net833));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(net605),
    .X(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_A (.DIODE(clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(in0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(in1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(in10));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(in11));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(in12));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(in13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c42_A (.DIODE(in14));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(in15));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(in16));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(in17));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(in18));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(in19));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(in2));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(in20));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(in21));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(in22));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(in23));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(in24));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(in3));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(in4));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(in5));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(in6));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_A (.DIODE(in7));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_A (.DIODE(in8));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_A (.DIODE(in9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c83_S0 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_c82_S0 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_c80_B1_N (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_c76_B1 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_c72_SET_B (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_c71_A2 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_c69_B (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_c68_A (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_c67_X (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_A (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_c190_B (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap41_A (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_B (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA_c565_A1 (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA_c558_S0 (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA_c542_B1 (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA_c541_A2 (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA_c538_A2 (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA_c536_Y (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA_output25_A (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_SCE (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_X (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold57_A (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA_output30_A (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_A (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_X (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap43_X (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_A3 (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA_c527_B (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA_c277_A (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA_c273_DE (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_B (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_15_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_14_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_13_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_12_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_11_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_10_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_9_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_8_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_7_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_6_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_5_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_4_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_3_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_2_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_1_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_0_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_X (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c519_GATE (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c523_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c528_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c543_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c633_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c644_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c645_CLK_N (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c647_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c648_CLK_N (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c649_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c650_CLK_N (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c654_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c658_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_2_0_clk_X (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c416_CLK_N (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_CLK_N (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c427_GATE (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_CLK_N (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c506_GATE (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c533_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c539_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c545_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s739_GATE (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_3_0_clk_X (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c184_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_GATE_N (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c191_GATE_N (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_GATE (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c70_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c72_CLK_N (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c73_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c74_CLK_N (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c77_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c81_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s733_GATE_N (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_4_0_clk_X (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c115_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c117_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c118_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c119_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c122_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c123_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_GATE (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c78_CLK_N (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c79_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s732_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_5_0_clk_X (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c311_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c313_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c321_CLK_N (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c323_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_CLK_N (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s736_GATE_N (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s737_GATE_N (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_6_0_clk_X (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c228_CLK_N (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c232_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c236_GATE_N (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c237_GATE_N (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c238_GATE_N (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c240_GATE (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c241_CLK_N (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c242_CLK_N (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c246_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c247_GATE (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c248_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c249_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c250_GATE (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c340_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_7_0_clk_X (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c686_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c695_GATE_N (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c698_GATE (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c701_GATE (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_CLK_N (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_CLK_N (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s744_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_11_0_clk_X (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_GATE_N (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c577_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_CLK_N (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c723_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_CLK_N (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_CLK_N (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s745_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_14_0_clk_X (.DIODE(clknet_4_14_0_clk));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_243 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_299 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_5 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_422 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_163 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_255 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_441 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_25 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_133 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_260 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_484 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_143 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_186 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_226 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_525 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_168 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_331 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_497 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_107 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_115 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_224 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_140 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_311 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_581 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_50 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_623 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_17 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_199 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_20 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_479 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_20 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_396 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_490 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_413 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_512 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_555 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_36 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_50 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_581 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_50 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_523 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_328 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_272 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_227 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_339 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_288 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_135 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_338 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_256 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_310 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_155 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_452 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_564 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_580 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_422 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_329 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_227 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_617 ();
endmodule
