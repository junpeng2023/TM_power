module netlist_0 (clk,
    in0,
    in1,
    in10,
    in11,
    in12,
    in13,
    in14,
    in15,
    in16,
    in17,
    in18,
    in19,
    in2,
    in20,
    in21,
    in22,
    in23,
    in24,
    in25,
    in26,
    in27,
    in28,
    in29,
    in3,
    in30,
    in31,
    in32,
    in33,
    in34,
    in35,
    in36,
    in37,
    in38,
    in39,
    in4,
    in40,
    in41,
    in42,
    in43,
    in44,
    in45,
    in46,
    in47,
    in48,
    in49,
    in5,
    in50,
    in51,
    in52,
    in53,
    in54,
    in55,
    in56,
    in57,
    in58,
    in59,
    in6,
    in60,
    in61,
    in62,
    in63,
    in64,
    in65,
    in66,
    in67,
    in68,
    in69,
    in7,
    in70,
    in71,
    in72,
    in73,
    in74,
    in75,
    in76,
    in77,
    in78,
    in79,
    in8,
    in80,
    in81,
    in82,
    in83,
    in84,
    in85,
    in86,
    in87,
    in88,
    in89,
    in9,
    in90,
    in91,
    in92,
    in93,
    in94,
    in95,
    in96,
    in97,
    in98,
    in99,
    out0,
    out1,
    out10,
    out11,
    out12,
    out13,
    out14,
    out15,
    out16,
    out17,
    out18,
    out19,
    out2,
    out20,
    out21,
    out22,
    out23,
    out24,
    out25,
    out26,
    out27,
    out28,
    out29,
    out3,
    out30,
    out31,
    out32,
    out33,
    out34,
    out35,
    out36,
    out37,
    out38,
    out39,
    out4,
    out40,
    out41,
    out42,
    out43,
    out44,
    out45,
    out46,
    out47,
    out48,
    out49,
    out5,
    out50,
    out51,
    out52,
    out53,
    out54,
    out55,
    out56,
    out57,
    out58,
    out59,
    out6,
    out60,
    out61,
    out62,
    out63,
    out64,
    out65,
    out66,
    out67,
    out68,
    out69,
    out7,
    out70,
    out71,
    out72,
    out73,
    out74,
    out75,
    out76,
    out77,
    out78,
    out79,
    out8,
    out80,
    out81,
    out82,
    out83,
    out84,
    out85,
    out86,
    out87,
    out88,
    out89,
    out9,
    out90,
    out91,
    out92,
    out93,
    out94,
    out95,
    out96,
    out97,
    out98,
    out99,
    rst);
 input clk;
 input in0;
 input in1;
 input in10;
 input in11;
 input in12;
 input in13;
 input in14;
 input in15;
 input in16;
 input in17;
 input in18;
 input in19;
 input in2;
 input in20;
 input in21;
 input in22;
 input in23;
 input in24;
 input in25;
 input in26;
 input in27;
 input in28;
 input in29;
 input in3;
 input in30;
 input in31;
 input in32;
 input in33;
 input in34;
 input in35;
 input in36;
 input in37;
 input in38;
 input in39;
 input in4;
 input in40;
 input in41;
 input in42;
 input in43;
 input in44;
 input in45;
 input in46;
 input in47;
 input in48;
 input in49;
 input in5;
 input in50;
 input in51;
 input in52;
 input in53;
 input in54;
 input in55;
 input in56;
 input in57;
 input in58;
 input in59;
 input in6;
 input in60;
 input in61;
 input in62;
 input in63;
 input in64;
 input in65;
 input in66;
 input in67;
 input in68;
 input in69;
 input in7;
 input in70;
 input in71;
 input in72;
 input in73;
 input in74;
 input in75;
 input in76;
 input in77;
 input in78;
 input in79;
 input in8;
 input in80;
 input in81;
 input in82;
 input in83;
 input in84;
 input in85;
 input in86;
 input in87;
 input in88;
 input in89;
 input in9;
 input in90;
 input in91;
 input in92;
 input in93;
 input in94;
 input in95;
 input in96;
 input in97;
 input in98;
 input in99;
 output out0;
 output out1;
 output out10;
 output out11;
 output out12;
 output out13;
 output out14;
 output out15;
 output out16;
 output out17;
 output out18;
 output out19;
 output out2;
 output out20;
 output out21;
 output out22;
 output out23;
 output out24;
 output out25;
 output out26;
 output out27;
 output out28;
 output out29;
 output out3;
 output out30;
 output out31;
 output out32;
 output out33;
 output out34;
 output out35;
 output out36;
 output out37;
 output out38;
 output out39;
 output out4;
 output out40;
 output out41;
 output out42;
 output out43;
 output out44;
 output out45;
 output out46;
 output out47;
 output out48;
 output out49;
 output out5;
 output out50;
 output out51;
 output out52;
 output out53;
 output out54;
 output out55;
 output out56;
 output out57;
 output out58;
 output out59;
 output out6;
 output out60;
 output out61;
 output out62;
 output out63;
 output out64;
 output out65;
 output out66;
 output out67;
 output out68;
 output out69;
 output out7;
 output out70;
 output out71;
 output out72;
 output out73;
 output out74;
 output out75;
 output out76;
 output out77;
 output out78;
 output out79;
 output out8;
 output out80;
 output out81;
 output out82;
 output out83;
 output out84;
 output out85;
 output out86;
 output out87;
 output out88;
 output out89;
 output out9;
 output out90;
 output out91;
 output out92;
 output out93;
 output out94;
 output out95;
 output out96;
 output out97;
 output out98;
 output out99;
 input rst;

 wire net0;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net182;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire clknet_0_net615;
 wire clknet_1_0__leaf_net615;
 wire clknet_1_1__leaf_net615;
 wire clknet_0_net475;
 wire clknet_1_0__leaf_net475;
 wire clknet_1_1__leaf_net475;
 wire clknet_0_net799;
 wire clknet_1_0__leaf_net799;
 wire clknet_1_1__leaf_net799;
 wire clknet_0_net370;
 wire clknet_1_0__leaf_net370;
 wire clknet_1_1__leaf_net370;
 wire clknet_0_net512;
 wire clknet_1_0__leaf_net512;
 wire clknet_1_1__leaf_net512;
 wire clknet_0_net295;
 wire clknet_1_0__leaf_net295;
 wire clknet_1_1__leaf_net295;
 wire clknet_0_net400;
 wire clknet_1_0__leaf_net400;
 wire clknet_1_1__leaf_net400;
 wire clknet_0_net300;
 wire clknet_1_0__leaf_net300;
 wire clknet_1_1__leaf_net300;
 wire clknet_0_net289;
 wire clknet_1_0__leaf_net289;
 wire clknet_1_1__leaf_net289;
 wire clknet_0_net305;
 wire clknet_1_0__leaf_net305;
 wire clknet_1_1__leaf_net305;
 wire clknet_0_net301;
 wire clknet_1_0__leaf_net301;
 wire clknet_1_1__leaf_net301;
 wire clknet_0_net268;
 wire clknet_1_0__leaf_net268;
 wire clknet_1_1__leaf_net268;
 wire clknet_0_net255;
 wire clknet_1_0__leaf_net255;
 wire clknet_1_1__leaf_net255;
 wire clknet_0_net614;
 wire clknet_1_0__leaf_net614;
 wire clknet_1_1__leaf_net614;
 wire clknet_0_net473;
 wire clknet_1_0__leaf_net473;
 wire clknet_1_1__leaf_net473;
 wire clknet_0_net793;
 wire clknet_1_0__leaf_net793;
 wire clknet_1_1__leaf_net793;
 wire clknet_0_net367;
 wire clknet_1_0__leaf_net367;
 wire clknet_1_1__leaf_net367;
 wire clknet_0_net198;
 wire clknet_1_0__leaf_net198;
 wire clknet_1_1__leaf_net198;
 wire clknet_0_net199;
 wire clknet_1_0__leaf_net199;
 wire clknet_1_1__leaf_net199;
 wire clknet_0_net200;
 wire clknet_1_0__leaf_net200;
 wire clknet_1_1__leaf_net200;
 wire clknet_0_net179;
 wire clknet_1_0__leaf_net179;
 wire clknet_1_1__leaf_net179;
 wire clknet_0_net178;
 wire clknet_1_0__leaf_net178;
 wire clknet_1_1__leaf_net178;
 wire clknet_0_net375;
 wire clknet_1_0__leaf_net375;
 wire clknet_1_1__leaf_net375;
 wire clknet_0_net277;
 wire clknet_1_0__leaf_net277;
 wire clknet_1_1__leaf_net277;
 wire clknet_0_net281;
 wire clknet_1_0__leaf_net281;
 wire clknet_1_1__leaf_net281;
 wire clknet_0_net282;
 wire clknet_1_0__leaf_net282;
 wire clknet_1_1__leaf_net282;
 wire clknet_0_net276;
 wire clknet_1_0__leaf_net276;
 wire clknet_1_1__leaf_net276;
 wire clknet_0_net166;
 wire clknet_1_0__leaf_net166;
 wire clknet_1_1__leaf_net166;
 wire clknet_0_net769;
 wire clknet_1_0__leaf_net769;
 wire clknet_1_1__leaf_net769;
 wire clknet_0_net162;
 wire clknet_1_0__leaf_net162;
 wire clknet_1_1__leaf_net162;
 wire clknet_0_net161;
 wire clknet_1_0__leaf_net161;
 wire clknet_1_1__leaf_net161;
 wire clknet_0_net159;
 wire clknet_1_0__leaf_net159;
 wire clknet_1_1__leaf_net159;
 wire clknet_0_net766;
 wire clknet_1_0__leaf_net766;
 wire clknet_1_1__leaf_net766;
 wire clknet_0_net786;
 wire clknet_1_0__leaf_net786;
 wire clknet_1_1__leaf_net786;
 wire clknet_0_net742;
 wire clknet_1_0__leaf_net742;
 wire clknet_1_1__leaf_net742;
 wire clknet_0_net97;
 wire clknet_1_0__leaf_net97;
 wire clknet_1_1__leaf_net97;
 wire clknet_0_net800;
 wire clknet_1_0__leaf_net800;
 wire clknet_1_1__leaf_net800;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net959;
 wire net960;
 wire net958;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;

 sky130_fd_sc_hd__and3_1 c100 (.A(net695),
    .B(net715),
    .C(net717),
    .X(net0));
 sky130_fd_sc_hd__and3_1 c101 (.A(net714),
    .B(net702),
    .C(net663),
    .X(net1));
 sky130_fd_sc_hd__mux4_1 c102 (.A0(net632),
    .A1(net673),
    .A2(net720),
    .A3(net700),
    .S0(net703),
    .S1(net716),
    .X(net2));
 sky130_fd_sc_hd__or4bb_2 c103 (.A(net720),
    .B(net1),
    .C_N(net647),
    .D_N(net722),
    .X(net774));
 sky130_fd_sc_hd__and3_1 c104 (.A(net711),
    .B(net662),
    .C(net670),
    .X(net3));
 sky130_fd_sc_hd__or4bb_2 c105 (.A(net713),
    .B(net649),
    .C_N(net719),
    .D_N(net3),
    .X(net758));
 sky130_fd_sc_hd__and3_1 c106 (.A(net717),
    .B(net721),
    .C(net844),
    .X(net4));
 sky130_fd_sc_hd__a2111o_1 c107 (.A1(net716),
    .A2(net3),
    .B1(net691),
    .C1(net695),
    .D1(net676),
    .X(net5));
 sky130_fd_sc_hd__a2111o_1 c108 (.A1(net2),
    .A2(net720),
    .B1(net716),
    .C1(net758),
    .D1(net962),
    .X(net756));
 sky130_fd_sc_hd__mux4_1 c109 (.A0(net1),
    .A1(net756),
    .A2(net5),
    .A3(net710),
    .S0(net711),
    .S1(net719),
    .X(net6));
 sky130_fd_sc_hd__and2_0 c110 (.A(net891),
    .B(net628),
    .X(net7));
 sky130_fd_sc_hd__and2_1 c111 (.A(net636),
    .B(net629),
    .X(net789));
 sky130_fd_sc_hd__and2_2 c112 (.A(net703),
    .B(net704),
    .X(net791));
 sky130_fd_sc_hd__and2_1 c113 (.A(net647),
    .B(net835),
    .X(net784));
 sky130_fd_sc_hd__and2_0 c114 (.A(net719),
    .B(net835),
    .X(net792));
 sky130_fd_sc_hd__and2_1 c115 (.A(net646),
    .B(net0),
    .X(net8));
 sky130_fd_sc_hd__and2_1 c116 (.A(net675),
    .B(net714),
    .X(net9));
 sky130_fd_sc_hd__and3_2 c117 (.A(net676),
    .B(net684),
    .C(net636),
    .X(net10));
 sky130_fd_sc_hd__and3_1 c118 (.A(net2),
    .B(net680),
    .C(net835),
    .X(net798));
 sky130_fd_sc_hd__and3_1 c119 (.A(net8),
    .B(net6),
    .C(net835),
    .X(net788));
 sky130_fd_sc_hd__a2111o_1 c120 (.A1(net10),
    .A2(net718),
    .B1(net632),
    .C1(net962),
    .D1(net798),
    .X(net11));
 sky130_fd_sc_hd__mux4_1 c121 (.A0(net11),
    .A1(net699),
    .A2(net789),
    .A3(net835),
    .S0(net704),
    .S1(net10),
    .X(net12));
 sky130_fd_sc_hd__and3_2 c122 (.A(net638),
    .B(net704),
    .C(net0),
    .X(net13));
 sky130_fd_sc_hd__and3_1 c123 (.A(net13),
    .B(net835),
    .C(net10),
    .X(net794));
 sky130_fd_sc_hd__and3_1 c124 (.A(net12),
    .B(net962),
    .C(net835),
    .X(net802));
 sky130_fd_sc_hd__a2111o_2 c125 (.A1(net10),
    .A2(net802),
    .B1(net835),
    .C1(net13),
    .D1(net756),
    .X(net768));
 sky130_fd_sc_hd__and3_1 c126 (.A(net962),
    .B(net13),
    .C(net718),
    .X(net781));
 sky130_fd_sc_hd__mux4_2 c127 (.A0(net663),
    .A1(net13),
    .A2(net10),
    .A3(net788),
    .S0(net8),
    .S1(net835),
    .X(net775));
 sky130_fd_sc_hd__and3_1 c128 (.A(net0),
    .B(net781),
    .C(net7),
    .X(net795));
 sky130_fd_sc_hd__and3_1 c129 (.A(net631),
    .B(net835),
    .C(net775),
    .X(net772));
 sky130_fd_sc_hd__a2111o_1 c130 (.A1(net632),
    .A2(net647),
    .B1(net9),
    .C1(net756),
    .D1(net768),
    .X(net14));
 sky130_fd_sc_hd__and3_1 c131 (.A(net718),
    .B(net10),
    .C(net14),
    .X(net15));
 sky130_fd_sc_hd__and2_4 c132 (.A(net679),
    .B(net657),
    .X(net16));
 sky130_fd_sc_hd__and2_4 c133 (.A(net848),
    .B(net633),
    .X(net17));
 sky130_fd_sc_hd__and3_4 c134 (.A(net831),
    .B(net633),
    .C(net847),
    .X(net777));
 sky130_fd_sc_hd__and3_4 c135 (.A(net777),
    .B(net632),
    .C(net844),
    .X(net761));
 sky130_fd_sc_hd__and2_4 c136 (.A(net17),
    .B(net646),
    .X(net18));
 sky130_fd_sc_hd__and3_2 c137 (.A(net646),
    .B(net633),
    .C(net831),
    .X(net19));
 sky130_fd_sc_hd__and2_1 c138 (.A(net18),
    .B(net17),
    .X(net730));
 sky130_fd_sc_hd__and3_4 c139 (.A(net961),
    .B(net18),
    .C(net761),
    .X(net20));
 sky130_fd_sc_hd__and2_4 c140 (.A(net17),
    .B(net635),
    .X(net21));
 sky130_fd_sc_hd__and3_4 c141 (.A(net831),
    .B(net18),
    .C(net632),
    .X(net760));
 sky130_fd_sc_hd__and2_4 c142 (.A(net635),
    .B(net636),
    .X(net22));
 sky130_fd_sc_hd__and3_4 c143 (.A(net832),
    .B(net21),
    .C(net843),
    .X(net23));
 sky130_fd_sc_hd__mux4_2 c144 (.A0(net777),
    .A1(net630),
    .A2(net760),
    .A3(net18),
    .S0(net23),
    .S1(net831),
    .X(net24));
 sky130_fd_sc_hd__mux4_2 c145 (.A0(net760),
    .A1(net19),
    .A2(net690),
    .A3(net962),
    .S0(net961),
    .S1(net956),
    .X(net744));
 sky130_fd_sc_hd__and3_4 c146 (.A(net760),
    .B(net630),
    .C(net844),
    .X(net25));
 sky130_fd_sc_hd__mux4_2 c147 (.A0(net24),
    .A1(net20),
    .A2(net23),
    .A3(net760),
    .S0(net19),
    .S1(net831),
    .X(net26));
 sky130_fd_sc_hd__or4bb_4 c148 (.A(net18),
    .B(net24),
    .C_N(net19),
    .D_N(net956),
    .X(net783));
 sky130_fd_sc_hd__and2_4 c149 (.A(net25),
    .B(net17),
    .X(net27));
 sky130_fd_sc_hd__mux4_2 c150 (.A0(net20),
    .A1(net27),
    .A2(net962),
    .A3(net633),
    .S0(net961),
    .S1(net831),
    .X(net771));
 sky130_fd_sc_hd__mux4_2 c151 (.A0(net26),
    .A1(net23),
    .A2(net25),
    .A3(net22),
    .S0(net832),
    .S1(net961),
    .X(net740));
 sky130_fd_sc_hd__a2111o_1 c152 (.A1(net744),
    .A2(net20),
    .B1(net771),
    .C1(net832),
    .D1(net961),
    .X(net28));
 sky130_fd_sc_hd__mux4_2 c153 (.A0(net21),
    .A1(net28),
    .A2(net817),
    .A3(net744),
    .S0(net25),
    .S1(net969),
    .X(net29));
 sky130_fd_sc_hd__or4bb_4 c154 (.A(net655),
    .B(net642),
    .C_N(net651),
    .D_N(net644),
    .X(net30));
 sky130_fd_sc_hd__and3_2 c155 (.A(net652),
    .B(net646),
    .C(net848),
    .X(net31));
 sky130_fd_sc_hd__and3_4 c156 (.A(net637),
    .B(net962),
    .C(net653),
    .X(net731));
 sky130_fd_sc_hd__and3_1 c157 (.A(net731),
    .B(net648),
    .C(net826),
    .X(net32));
 sky130_fd_sc_hd__or4bb_2 c158 (.A(net633),
    .B(net630),
    .C_N(net826),
    .D_N(net956),
    .X(net33));
 sky130_fd_sc_hd__a2111o_4 c159 (.A1(net32),
    .A2(net826),
    .B1(net637),
    .C1(net24),
    .D1(net961),
    .X(net797));
 sky130_fd_sc_hd__a2111o_2 c160 (.A1(net24),
    .A2(net634),
    .B1(net731),
    .C1(net956),
    .D1(net826),
    .X(net34));
 sky130_fd_sc_hd__and3_4 c161 (.A(net771),
    .B(net650),
    .C(net652),
    .X(net35));
 sky130_fd_sc_hd__a2111o_2 c162 (.A1(net644),
    .A2(net661),
    .B1(net826),
    .C1(net650),
    .D1(net690),
    .X(net36));
 sky130_fd_sc_hd__or4bb_4 c163 (.A(net797),
    .B(net34),
    .C_N(net32),
    .D_N(net961),
    .X(net725));
 sky130_fd_sc_hd__and3_2 c164 (.A(net660),
    .B(net36),
    .C(net652),
    .X(net37));
 sky130_fd_sc_hd__mux4_2 c165 (.A0(net18),
    .A1(net37),
    .A2(net647),
    .A3(net731),
    .S0(net826),
    .S1(net832),
    .X(net38));
 sky130_fd_sc_hd__mux4_2 c166 (.A0(net630),
    .A1(net30),
    .A2(net654),
    .A3(net644),
    .S0(net35),
    .S1(net826),
    .X(net732));
 sky130_fd_sc_hd__and3_2 c167 (.A(net634),
    .B(net731),
    .C(net32),
    .X(net780));
 sky130_fd_sc_hd__a2111o_4 c168 (.A1(net38),
    .A2(net34),
    .B1(net826),
    .C1(net813),
    .D1(net797),
    .X(net39));
 sky130_fd_sc_hd__and3_2 c169 (.A(net36),
    .B(net33),
    .C(net813),
    .X(net40));
 sky130_fd_sc_hd__a2111o_2 c170 (.A1(net35),
    .A2(net633),
    .B1(net813),
    .C1(net33),
    .D1(net826),
    .X(net41));
 sky130_fd_sc_hd__and3_2 c171 (.A(net40),
    .B(net962),
    .C(net41),
    .X(net42));
 sky130_fd_sc_hd__and3_4 c172 (.A(net39),
    .B(net642),
    .C(net961),
    .X(net43));
 sky130_fd_sc_hd__mux4_2 c173 (.A0(net826),
    .A1(net35),
    .A2(net813),
    .A3(net36),
    .S0(net26),
    .S1(net648),
    .X(net44));
 sky130_fd_sc_hd__a2111o_4 c174 (.A1(net813),
    .A2(net26),
    .B1(net822),
    .C1(net827),
    .D1(net43),
    .X(net45));
 sky130_fd_sc_hd__mux4_2 c175 (.A0(net44),
    .A1(net45),
    .A2(net41),
    .A3(net43),
    .S0(net651),
    .S1(net639),
    .X(net803));
 sky130_fd_sc_hd__mux4_2 c176 (.A0(net648),
    .A1(net678),
    .A2(net813),
    .A3(net654),
    .S0(net653),
    .S1(net803),
    .X(net46));
 sky130_fd_sc_hd__and3_2 c177 (.A(net643),
    .B(net683),
    .C(net761),
    .X(net47));
 sky130_fd_sc_hd__and3_1 c178 (.A(net648),
    .B(net47),
    .C(net827),
    .X(net48));
 sky130_fd_sc_hd__and3_2 c179 (.A(net24),
    .B(net38),
    .C(net630),
    .X(net49));
 sky130_fd_sc_hd__and3_2 c180 (.A(net630),
    .B(net671),
    .C(net47),
    .X(net796));
 sky130_fd_sc_hd__and3_1 c181 (.A(net639),
    .B(net658),
    .C(net24),
    .X(net50));
 sky130_fd_sc_hd__and3_2 c182 (.A(net30),
    .B(net50),
    .C(net34),
    .X(net51));
 sky130_fd_sc_hd__and3_2 c183 (.A(net760),
    .B(net666),
    .C(net643),
    .X(net52));
 sky130_fd_sc_hd__mux4_2 c184 (.A0(net669),
    .A1(net50),
    .A2(net52),
    .A3(net667),
    .S0(net43),
    .S1(net46),
    .X(net53));
 sky130_fd_sc_hd__mux4_2 c185 (.A0(net656),
    .A1(net678),
    .A2(net51),
    .A3(net30),
    .S0(net38),
    .S1(net666),
    .X(net54));
 sky130_fd_sc_hd__or4bb_2 c186 (.A(net49),
    .B(net680),
    .C_N(net682),
    .D_N(net54),
    .X(net55));
 sky130_fd_sc_hd__and3_4 c187 (.A(net53),
    .B(net796),
    .C(net827),
    .X(net728));
 sky130_fd_sc_hd__and3_2 c188 (.A(net646),
    .B(net649),
    .C(net829),
    .X(net56));
 sky130_fd_sc_hd__mux4_2 c189 (.A0(net41),
    .A1(net56),
    .A2(net728),
    .A3(net669),
    .S0(net683),
    .S1(net639),
    .X(net57));
 sky130_fd_sc_hd__and3_4 c190 (.A(net57),
    .B(net682),
    .C(net674),
    .X(net58));
 sky130_fd_sc_hd__mux4_2 c191 (.A0(net632),
    .A1(net728),
    .A2(net58),
    .A3(net662),
    .S0(net52),
    .S1(net827),
    .X(net782));
 sky130_fd_sc_hd__and3_2 c192 (.A(net27),
    .B(net55),
    .C(net827),
    .X(net59));
 sky130_fd_sc_hd__mux4_2 c193 (.A0(net782),
    .A1(net796),
    .A2(net659),
    .A3(net653),
    .S0(net55),
    .S1(net662),
    .X(net60));
 sky130_fd_sc_hd__a2111o_2 c194 (.A1(net52),
    .A2(net58),
    .B1(net60),
    .C1(net59),
    .D1(net827),
    .X(net61));
 sky130_fd_sc_hd__or4bb_4 c195 (.A(net54),
    .B(net58),
    .C_N(net846),
    .D_N(net59),
    .X(net62));
 sky130_fd_sc_hd__mux4_2 c196 (.A0(net59),
    .A1(net648),
    .A2(net62),
    .A3(net796),
    .S0(net924),
    .S1(net58),
    .X(net63));
 sky130_fd_sc_hd__mux4_1 c197 (.A0(net46),
    .A1(net62),
    .A2(net60),
    .A3(net58),
    .S0(net54),
    .S1(net829),
    .X(net64));
 sky130_fd_sc_hd__and3_2 c198 (.A(net35),
    .B(net26),
    .C(net638),
    .X(net65));
 sky130_fd_sc_hd__and3_2 c199 (.A(net50),
    .B(net761),
    .C(net827),
    .X(net66));
 sky130_fd_sc_hd__a2111o_1 c200 (.A1(net962),
    .A2(net697),
    .B1(net685),
    .C1(net834),
    .D1(net830),
    .X(net67));
 sky130_fd_sc_hd__and3_4 c201 (.A(net689),
    .B(net803),
    .C(net777),
    .X(net68));
 sky130_fd_sc_hd__and3_2 c202 (.A(net65),
    .B(net691),
    .C(net704),
    .X(net69));
 sky130_fd_sc_hd__and3_1 c203 (.A(net66),
    .B(net698),
    .C(net47),
    .X(net70));
 sky130_fd_sc_hd__mux4_2 c204 (.A0(net678),
    .A1(net45),
    .A2(net66),
    .A3(net797),
    .S0(net846),
    .S1(net810),
    .X(net71));
 sky130_fd_sc_hd__and3_2 c205 (.A(net71),
    .B(net60),
    .C(net680),
    .X(net746));
 sky130_fd_sc_hd__and3_1 c206 (.A(net26),
    .B(net684),
    .C(net670),
    .X(net72));
 sky130_fd_sc_hd__and3_2 c207 (.A(net60),
    .B(net691),
    .C(net693),
    .X(net73));
 sky130_fd_sc_hd__mux4_2 c208 (.A0(net73),
    .A1(net680),
    .A2(net672),
    .A3(net66),
    .S0(net810),
    .S1(net51),
    .X(net74));
 sky130_fd_sc_hd__or4bb_1 c209 (.A(net52),
    .B(net680),
    .C_N(net816),
    .D_N(net74),
    .X(net75));
 sky130_fd_sc_hd__a2111o_1 c210 (.A1(net74),
    .A2(net632),
    .B1(net66),
    .C1(net810),
    .D1(net829),
    .X(net76));
 sky130_fd_sc_hd__a2111o_2 c211 (.A1(net70),
    .A2(net782),
    .B1(net73),
    .C1(net64),
    .D1(net858),
    .X(net77));
 sky130_fd_sc_hd__a2111o_1 c212 (.A1(net68),
    .A2(net708),
    .B1(net77),
    .C1(net810),
    .D1(net664),
    .X(net78));
 sky130_fd_sc_hd__and3_1 c213 (.A(net70),
    .B(net73),
    .C(net842),
    .X(net79));
 sky130_fd_sc_hd__a2111o_2 c214 (.A1(net72),
    .A2(net70),
    .B1(net71),
    .C1(net829),
    .D1(net842),
    .X(net733));
 sky130_fd_sc_hd__buf_1 c215 (.A(net840),
    .X(net80));
 sky130_fd_sc_hd__a2111o_2 c216 (.A1(net42),
    .A2(net808),
    .B1(net80),
    .C1(net709),
    .D1(net842),
    .X(net81));
 sky130_fd_sc_hd__mux4_1 c217 (.A0(net77),
    .A1(net808),
    .A2(net636),
    .A3(net673),
    .S0(net79),
    .S1(net842),
    .X(net82));
 sky130_fd_sc_hd__a2111o_1 c218 (.A1(net58),
    .A2(net81),
    .B1(net77),
    .C1(net808),
    .D1(net79),
    .X(net83));
 sky130_fd_sc_hd__or4bb_4 c219 (.A(net80),
    .B(net81),
    .C_N(net808),
    .D_N(net840),
    .X(net762));
 sky130_fd_sc_hd__and3_1 c220 (.A(net72),
    .B(net777),
    .C(net774),
    .X(net787));
 sky130_fd_sc_hd__a2111o_1 c221 (.A1(net641),
    .A2(net697),
    .B1(net625),
    .C1(net721),
    .D1(net722),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_1 c222 (.A(net836),
    .X(net85));
 sky130_fd_sc_hd__mux4_1 c223 (.A0(net949),
    .A1(net783),
    .A2(net808),
    .A3(net710),
    .S0(net72),
    .S1(net63),
    .X(net776));
 sky130_fd_sc_hd__and3_1 c224 (.A(net715),
    .B(net797),
    .C(net66),
    .X(net86));
 sky130_fd_sc_hd__and3_1 c225 (.A(net710),
    .B(net681),
    .C(net685),
    .X(net87));
 sky130_fd_sc_hd__and3_1 c226 (.A(net85),
    .B(net776),
    .C(net64),
    .X(net88));
 sky130_fd_sc_hd__and3_1 c227 (.A(net953),
    .B(net787),
    .C(net696),
    .X(net89));
 sky130_fd_sc_hd__and3_1 c228 (.A(net62),
    .B(net698),
    .C(net842),
    .X(net90));
 sky130_fd_sc_hd__and3_1 c229 (.A(net38),
    .B(net711),
    .C(net811),
    .X(net91));
 sky130_fd_sc_hd__and3_1 c230 (.A(net90),
    .B(net811),
    .C(net68),
    .X(net765));
 sky130_fd_sc_hd__and3_1 c231 (.A(net64),
    .B(net91),
    .C(net706),
    .X(net92));
 sky130_fd_sc_hd__a2111o_4 c232 (.A1(net62),
    .A2(net824),
    .B1(net829),
    .C1(net713),
    .D1(net811),
    .X(net93));
 sky130_fd_sc_hd__a2111o_1 c233 (.A1(net911),
    .A2(net74),
    .B1(net646),
    .C1(net811),
    .D1(net87),
    .X(net94));
 sky130_fd_sc_hd__buf_1 c234 (.A(net836),
    .X(net95));
 sky130_fd_sc_hd__a2111o_1 c235 (.A1(net811),
    .A2(net87),
    .B1(net808),
    .C1(net88),
    .D1(net810),
    .X(net96));
 sky130_fd_sc_hd__mux4_1 c236 (.A0(net670),
    .A1(net713),
    .A2(net87),
    .A3(net699),
    .S0(net54),
    .S1(clknet_1_1__leaf_net799),
    .X(net97));
 sky130_fd_sc_hd__a2111o_1 c237 (.A1(net962),
    .A2(net85),
    .B1(net911),
    .C1(net811),
    .D1(clknet_1_1__leaf_net799),
    .X(net786));
 sky130_fd_sc_hd__and3_1 c238 (.A(net91),
    .B(net810),
    .C(net947),
    .X(net98));
 sky130_fd_sc_hd__clkbuf_1 c239 (.A(net840),
    .X(net99));
 sky130_fd_sc_hd__and3_1 c240 (.A(net93),
    .B(net70),
    .C(clknet_1_0__leaf_net799),
    .X(net766));
 sky130_fd_sc_hd__a2111o_1 c241 (.A1(net99),
    .A2(clknet_1_0__leaf_net766),
    .B1(net697),
    .C1(net628),
    .D1(net811),
    .X(net100));
 sky130_fd_sc_hd__mux4_2 c256 (.A0(net9),
    .A1(net11),
    .A2(net673),
    .A3(net808),
    .S0(net768),
    .S1(net693),
    .X(net779));
 sky130_fd_sc_hd__mux4_1 c257 (.A0(net746),
    .A1(clknet_1_0__leaf_net97),
    .A2(net6),
    .A3(net10),
    .S0(net13),
    .S1(net842),
    .X(net800));
 sky130_fd_sc_hd__mux4_1 c258 (.A0(clknet_1_1__leaf_net97),
    .A1(net15),
    .A2(net774),
    .A3(clknet_1_0__leaf_net800),
    .S0(net852),
    .S1(net795),
    .X(net101));
 sky130_fd_sc_hd__mux4_1 c259 (.A0(net86),
    .A1(net10),
    .A2(net794),
    .A3(net861),
    .S0(clknet_1_0__leaf_net800),
    .S1(net664),
    .X(net102));
 sky130_fd_sc_hd__mux4_1 c260 (.A0(net7),
    .A1(net14),
    .A2(clknet_1_0__leaf_net786),
    .A3(net10),
    .S0(net638),
    .S1(net910),
    .X(net742));
 sky130_fd_sc_hd__mux4_1 c261 (.A0(net684),
    .A1(net13),
    .A2(net784),
    .A3(net779),
    .S0(net842),
    .S1(net836),
    .X(net790));
 sky130_fd_sc_hd__mux4_1 c262 (.A0(net6),
    .A1(net684),
    .A2(clknet_1_1__leaf_net800),
    .A3(net709),
    .S0(net791),
    .S1(net891),
    .X(net103));
 sky130_fd_sc_hd__mux4_1 c263 (.A0(net100),
    .A1(net779),
    .A2(net7),
    .A3(clknet_1_1__leaf_net742),
    .S0(net842),
    .S1(net836),
    .X(net104));
 sky130_fd_sc_hd__and2_1 c264 (.A(net969),
    .B(net27),
    .X(net105));
 sky130_fd_sc_hd__and2_4 c265 (.A(net625),
    .B(net783),
    .X(net106));
 sky130_fd_sc_hd__and3_1 c266 (.A(net19),
    .B(net635),
    .C(net17),
    .X(net107));
 sky130_fd_sc_hd__and2_2 c267 (.A(net657),
    .B(net20),
    .X(net108));
 sky130_fd_sc_hd__and2_1 c268 (.A(net635),
    .B(net106),
    .X(net109));
 sky130_fd_sc_hd__and2_4 c269 (.A(net106),
    .B(net777),
    .X(net110));
 sky130_fd_sc_hd__and2_2 c270 (.A(net631),
    .B(net961),
    .X(net111));
 sky130_fd_sc_hd__and3_4 c271 (.A(net821),
    .B(net20),
    .C(net17),
    .X(net112));
 sky130_fd_sc_hd__and3_4 c272 (.A(net690),
    .B(net109),
    .C(net821),
    .X(net113));
 sky130_fd_sc_hd__and2_4 c273 (.A(net113),
    .B(net818),
    .X(net114));
 sky130_fd_sc_hd__and2_2 c274 (.A(net28),
    .B(net634),
    .X(net115));
 sky130_fd_sc_hd__and3_4 c275 (.A(net105),
    .B(net113),
    .C(net844),
    .X(net116));
 sky130_fd_sc_hd__and2_2 c276 (.A(net818),
    .B(net635),
    .X(net117));
 sky130_fd_sc_hd__and2_0 c277 (.A(net818),
    .B(net116),
    .X(net118));
 sky130_fd_sc_hd__and2_2 c278 (.A(net118),
    .B(net116),
    .X(net119));
 sky130_fd_sc_hd__or4bb_4 c279 (.A(net109),
    .B(net113),
    .C_N(net112),
    .D_N(net744),
    .X(net120));
 sky130_fd_sc_hd__or4bb_4 c280 (.A(net23),
    .B(net111),
    .C_N(net668),
    .D_N(net112),
    .X(net121));
 sky130_fd_sc_hd__and3_2 c281 (.A(net114),
    .B(net115),
    .C(net116),
    .X(net122));
 sky130_fd_sc_hd__a2111o_4 c282 (.A1(net815),
    .A2(net120),
    .B1(net122),
    .C1(net637),
    .D1(net833),
    .X(net123));
 sky130_fd_sc_hd__and3_4 c283 (.A(net110),
    .B(net122),
    .C(net821),
    .X(net124));
 sky130_fd_sc_hd__mux4_2 c284 (.A0(net116),
    .A1(net122),
    .A2(net106),
    .A3(net23),
    .S0(net29),
    .S1(net833),
    .X(net125));
 sky130_fd_sc_hd__mux4_2 c285 (.A0(net122),
    .A1(net124),
    .A2(net634),
    .A3(net114),
    .S0(net111),
    .S1(net113),
    .X(net738));
 sky130_fd_sc_hd__and3_1 c286 (.A(net651),
    .B(net118),
    .C(net843),
    .X(net126));
 sky130_fd_sc_hd__and2_1 c287 (.A(net39),
    .B(net661),
    .X(net127));
 sky130_fd_sc_hd__and2_1 c288 (.A(net625),
    .B(net36),
    .X(net128));
 sky130_fd_sc_hd__and3_2 c289 (.A(net34),
    .B(net643),
    .C(net823),
    .X(net129));
 sky130_fd_sc_hd__or4bb_2 c290 (.A(net626),
    .B(net114),
    .C_N(net113),
    .D_N(net655),
    .X(net130));
 sky130_fd_sc_hd__and3_1 c291 (.A(net129),
    .B(net121),
    .C(net823),
    .X(net763));
 sky130_fd_sc_hd__or4bb_4 c292 (.A(net654),
    .B(net780),
    .C_N(net814),
    .D_N(net848),
    .X(net131));
 sky130_fd_sc_hd__and2_2 c293 (.A(net131),
    .B(net814),
    .X(net132));
 sky130_fd_sc_hd__mux4_2 c294 (.A0(net125),
    .A1(net626),
    .A2(net847),
    .A3(net843),
    .S0(net777),
    .S1(net129),
    .X(net133));
 sky130_fd_sc_hd__or4bb_4 c295 (.A(net638),
    .B(net129),
    .C_N(net133),
    .D_N(net131),
    .X(net134));
 sky130_fd_sc_hd__and3_4 c296 (.A(net629),
    .B(net134),
    .C(net818),
    .X(net135));
 sky130_fd_sc_hd__mux4_2 c297 (.A0(net637),
    .A1(net119),
    .A2(net33),
    .A3(net135),
    .S0(net133),
    .S1(net821),
    .X(net136));
 sky130_fd_sc_hd__mux4_2 c298 (.A0(net127),
    .A1(net23),
    .A2(net132),
    .A3(net818),
    .S0(net44),
    .S1(net828),
    .X(net137));
 sky130_fd_sc_hd__and3_4 c299 (.A(net136),
    .B(net640),
    .C(net134),
    .X(net138));
 sky130_fd_sc_hd__and3_4 c300 (.A(net136),
    .B(net131),
    .C(net642),
    .X(net139));
 sky130_fd_sc_hd__and3_1 c301 (.A(net118),
    .B(net129),
    .C(net139),
    .X(net140));
 sky130_fd_sc_hd__and3_1 c302 (.A(net139),
    .B(net133),
    .C(net138),
    .X(net141));
 sky130_fd_sc_hd__mux4_2 c303 (.A0(net900),
    .A1(net639),
    .A2(net140),
    .A3(net119),
    .S0(net690),
    .S1(net761),
    .X(net142));
 sky130_fd_sc_hd__a2111o_4 c304 (.A1(net653),
    .A2(net135),
    .B1(net823),
    .C1(net814),
    .D1(net138),
    .X(net735));
 sky130_fd_sc_hd__mux4_1 c305 (.A0(net141),
    .A1(net128),
    .A2(net113),
    .A3(net122),
    .S0(net130),
    .S1(net814),
    .X(net143));
 sky130_fd_sc_hd__and3_4 c306 (.A(net127),
    .B(net121),
    .C(net140),
    .X(net757));
 sky130_fd_sc_hd__and3_1 c307 (.A(net143),
    .B(net636),
    .C(net757),
    .X(net144));
 sky130_fd_sc_hd__and3_2 c308 (.A(net675),
    .B(net658),
    .C(net827),
    .X(net145));
 sky130_fd_sc_hd__and3_4 c309 (.A(net23),
    .B(net780),
    .C(net804),
    .X(net146));
 sky130_fd_sc_hd__and3_4 c310 (.A(net48),
    .B(net33),
    .C(net814),
    .X(net770));
 sky130_fd_sc_hd__or4bb_2 c311 (.A(net34),
    .B(net126),
    .C_N(net51),
    .D_N(net25),
    .X(net147));
 sky130_fd_sc_hd__and3_4 c312 (.A(net146),
    .B(net48),
    .C(net54),
    .X(net148));
 sky130_fd_sc_hd__or4bb_1 c313 (.A(net128),
    .B(net875),
    .C_N(net112),
    .D_N(net126),
    .X(net149));
 sky130_fd_sc_hd__and3_1 c314 (.A(net666),
    .B(net846),
    .C(net832),
    .X(net150));
 sky130_fd_sc_hd__and3_4 c315 (.A(net844),
    .B(net873),
    .C(net56),
    .X(net151));
 sky130_fd_sc_hd__and3_1 c316 (.A(net33),
    .B(net63),
    .C(net27),
    .X(net152));
 sky130_fd_sc_hd__a2111o_2 c317 (.A1(net36),
    .A2(net145),
    .B1(net770),
    .C1(net832),
    .D1(net150),
    .X(net153));
 sky130_fd_sc_hd__a2111o_1 c318 (.A1(net669),
    .A2(net112),
    .B1(net153),
    .C1(net138),
    .D1(net151),
    .X(net154));
 sky130_fd_sc_hd__mux4_2 c319 (.A0(net122),
    .A1(net643),
    .A2(net152),
    .A3(net145),
    .S0(net41),
    .S1(net153),
    .X(net155));
 sky130_fd_sc_hd__and3_1 c320 (.A(net154),
    .B(net48),
    .C(net128),
    .X(net156));
 sky130_fd_sc_hd__a2111o_1 c321 (.A1(net146),
    .A2(net155),
    .B1(net815),
    .C1(net128),
    .D1(net151),
    .X(net157));
 sky130_fd_sc_hd__mux4_1 c322 (.A0(net148),
    .A1(net51),
    .A2(net153),
    .A3(net821),
    .S0(net650),
    .S1(net827),
    .X(net158));
 sky130_fd_sc_hd__mux4_1 c323 (.A0(net903),
    .A1(net152),
    .A2(net149),
    .A3(net61),
    .S0(net827),
    .S1(clknet_1_0__leaf_net799),
    .X(net159));
 sky130_fd_sc_hd__a2111o_1 c324 (.A1(net41),
    .A2(clknet_1_0__leaf_net159),
    .B1(net156),
    .C1(net674),
    .D1(net814),
    .X(net160));
 sky130_fd_sc_hd__a2111o_1 c325 (.A1(net154),
    .A2(net61),
    .B1(net782),
    .C1(net770),
    .D1(clknet_1_0__leaf_net799),
    .X(net161));
 sky130_fd_sc_hd__or4bb_4 c326 (.A(net158),
    .B(net153),
    .C_N(net780),
    .D_N(clknet_1_0__leaf_net799),
    .X(net162));
 sky130_fd_sc_hd__buf_2 c327 (.A(net842),
    .X(net749));
 sky130_fd_sc_hd__mux4_1 c328 (.A0(net126),
    .A1(clknet_1_0__leaf_net161),
    .A2(net158),
    .A3(net642),
    .S0(clknet_1_0__leaf_net162),
    .S1(net770),
    .X(net163));
 sky130_fd_sc_hd__mux4_1 c329 (.A0(clknet_1_0__leaf_net159),
    .A1(net858),
    .A2(net57),
    .A3(clknet_1_0__leaf_net162),
    .S0(clknet_1_0__leaf_net161),
    .S1(net129),
    .X(net164));
 sky130_fd_sc_hd__a2111o_1 c330 (.A1(net79),
    .A2(clknet_1_1__leaf_net159),
    .B1(net804),
    .C1(net829),
    .D1(net808),
    .X(net165));
 sky130_fd_sc_hd__and3_1 c331 (.A(net682),
    .B(net819),
    .C(clknet_1_0__leaf_net799),
    .X(net166));
 sky130_fd_sc_hd__and3_1 c332 (.A(net80),
    .B(net66),
    .C(net819),
    .X(net167));
 sky130_fd_sc_hd__and3_1 c333 (.A(clknet_1_0__leaf_net166),
    .B(net770),
    .C(net757),
    .X(net769));
 sky130_fd_sc_hd__or4bb_1 c334 (.A(net687),
    .B(net141),
    .C_N(net673),
    .D_N(net819),
    .X(net168));
 sky130_fd_sc_hd__a2111o_2 c335 (.A1(net780),
    .A2(net813),
    .B1(net679),
    .C1(net891),
    .D1(net572),
    .X(net169));
 sky130_fd_sc_hd__a2111o_4 c336 (.A1(net658),
    .A2(net61),
    .B1(net640),
    .C1(net816),
    .D1(net49),
    .X(net755));
 sky130_fd_sc_hd__and3_1 c337 (.A(net686),
    .B(net636),
    .C(net654),
    .X(net170));
 sky130_fd_sc_hd__buf_1 c338 (.A(net840),
    .X(net171));
 sky130_fd_sc_hd__and3_1 c339 (.A(net635),
    .B(net668),
    .C(net71),
    .X(net773));
 sky130_fd_sc_hd__buf_1 c340 (.A(net840),
    .X(net172));
 sky130_fd_sc_hd__or4bb_4 c341 (.A(net171),
    .B(net115),
    .C_N(net167),
    .D_N(net824),
    .X(net173));
 sky130_fd_sc_hd__mux4_1 c342 (.A0(net168),
    .A1(clknet_1_0__leaf_net769),
    .A2(net155),
    .A3(clknet_1_1__leaf_net166),
    .S0(net858),
    .S1(net572),
    .X(net174));
 sky130_fd_sc_hd__clkbuf_2 c343 (.A(net842),
    .X(net754));
 sky130_fd_sc_hd__a2111o_1 c344 (.A1(net172),
    .A2(net168),
    .B1(net679),
    .C1(net45),
    .D1(net687),
    .X(net175));
 sky130_fd_sc_hd__mux4_1 c345 (.A0(net182),
    .A1(net693),
    .A2(net145),
    .A3(net946),
    .S0(net824),
    .S1(net840),
    .X(net176));
 sky130_fd_sc_hd__and3_1 c346 (.A(net176),
    .B(net172),
    .C(net175),
    .X(net177));
 sky130_fd_sc_hd__mux4_1 c347 (.A0(net754),
    .A1(net172),
    .A2(net173),
    .A3(net921),
    .S0(net841),
    .S1(clknet_1_1__leaf_net799),
    .X(net178));
 sky130_fd_sc_hd__or4bb_1 c348 (.A(net175),
    .B(net177),
    .C_N(net840),
    .D_N(clknet_1_0__leaf_net799),
    .X(net179));
 sky130_fd_sc_hd__a2111o_2 c349 (.A1(net177),
    .A2(net773),
    .B1(net176),
    .C1(net172),
    .D1(net819),
    .X(net180));
 sky130_fd_sc_hd__a2111o_1 c350 (.A1(clknet_1_1__leaf_net179),
    .A2(clknet_1_0__leaf_net178),
    .B1(net696),
    .C1(net180),
    .D1(net840),
    .X(net181));
 sky130_fd_sc_hd__a2111o_4 c351 (.A1(clknet_1_0__leaf_net179),
    .A2(net760),
    .B1(net171),
    .C1(net572),
    .X(net748));
 sky130_fd_sc_hd__and3_1 c352 (.A(net706),
    .B(net690),
    .C(net819),
    .X(net778));
 sky130_fd_sc_hd__clkbuf_1 c353 (.A(net604),
    .X(net183));
 sky130_fd_sc_hd__a2111o_1 c354 (.A1(net647),
    .A2(net717),
    .B1(net180),
    .C1(net706),
    .D1(net948),
    .X(net184));
 sky130_fd_sc_hd__mux4_1 c355 (.A0(net115),
    .A1(net692),
    .A2(net812),
    .A3(net778),
    .S0(net708),
    .S1(net734),
    .X(net185));
 sky130_fd_sc_hd__a2111o_1 c356 (.A1(net180),
    .A2(net673),
    .B1(net858),
    .C1(net721),
    .D1(net744),
    .X(net186));
 sky130_fd_sc_hd__mux4_2 c357 (.A0(net87),
    .A1(net770),
    .A2(net762),
    .A3(net185),
    .S0(net153),
    .S1(net681),
    .X(net187));
 sky130_fd_sc_hd__a2111o_1 c358 (.A1(net662),
    .A2(net185),
    .B1(net844),
    .C1(net151),
    .D1(net814),
    .X(net188));
 sky130_fd_sc_hd__a2111o_1 c359 (.A1(net173),
    .A2(net810),
    .B1(net188),
    .C1(net713),
    .D1(net651),
    .X(net189));
 sky130_fd_sc_hd__a2111o_1 c360 (.A1(net5),
    .A2(net690),
    .B1(net47),
    .C1(net641),
    .D1(net947),
    .X(net190));
 sky130_fd_sc_hd__or4bb_2 c361 (.A(net654),
    .B(net702),
    .C_N(net699),
    .D_N(net844),
    .X(net191));
 sky130_fd_sc_hd__or4bb_1 c362 (.A(net113),
    .B(net811),
    .C_N(net185),
    .D_N(net706),
    .X(net192));
 sky130_fd_sc_hd__and3_1 c363 (.A(net696),
    .B(net141),
    .C(net191),
    .X(net193));
 sky130_fd_sc_hd__or4bb_4 c364 (.A(net61),
    .B(net947),
    .C_N(net190),
    .D_N(net87),
    .X(net194));
 sky130_fd_sc_hd__and3_1 c365 (.A(net3),
    .B(net112),
    .C(net170),
    .X(net195));
 sky130_fd_sc_hd__mux4_1 c366 (.A0(net188),
    .A1(net115),
    .A2(net783),
    .A3(net173),
    .S0(net4),
    .S1(net913),
    .X(net196));
 sky130_fd_sc_hd__mux4_2 c367 (.A0(net190),
    .A1(net147),
    .A2(net196),
    .A3(net631),
    .S0(net193),
    .S1(net713),
    .X(net197));
 sky130_fd_sc_hd__and3_1 c368 (.A(net193),
    .B(net696),
    .C(clknet_1_1__leaf_net799),
    .X(net198));
 sky130_fd_sc_hd__or4bb_2 c369 (.A(net63),
    .B(net713),
    .C_N(net814),
    .D_N(net638),
    .X(net750));
 sky130_fd_sc_hd__and3_1 c370 (.A(net697),
    .B(net45),
    .C(clknet_1_0__leaf_net198),
    .X(net199));
 sky130_fd_sc_hd__or4bb_1 c371 (.A(net153),
    .B(clknet_1_0__leaf_net199),
    .C_N(net68),
    .D_N(net840),
    .X(net200));
 sky130_fd_sc_hd__or4bb_4 c372 (.A(net170),
    .B(net4),
    .C_N(net3),
    .D_N(net195),
    .X(net201));
 sky130_fd_sc_hd__a2111o_1 c373 (.A1(net195),
    .A2(net816),
    .B1(clknet_1_1__leaf_net199),
    .C1(clknet_1_0__leaf_net200),
    .D1(net201),
    .X(net202));
 sky130_fd_sc_hd__and2_4 c396 (.A(net29),
    .B(net815),
    .X(net203));
 sky130_fd_sc_hd__and2_4 c397 (.A(net628),
    .B(net120),
    .X(net204));
 sky130_fd_sc_hd__and3_1 c398 (.A(net19),
    .B(net958),
    .C(net125),
    .X(net205));
 sky130_fd_sc_hd__and2_1 c399 (.A(net821),
    .B(net116),
    .X(net206));
 sky130_fd_sc_hd__and3_1 c400 (.A(net204),
    .B(net105),
    .C(net120),
    .X(net207));
 sky130_fd_sc_hd__and2_1 c401 (.A(net27),
    .B(net631),
    .X(net208));
 sky130_fd_sc_hd__a2111o_4 c402 (.A1(net817),
    .A2(net116),
    .B1(net204),
    .C1(net626),
    .D1(net29),
    .X(net767));
 sky130_fd_sc_hd__and2_1 c403 (.A(net783),
    .B(net17),
    .X(net209));
 sky130_fd_sc_hd__and2_1 c404 (.A(net112),
    .B(net28),
    .X(net210));
 sky130_fd_sc_hd__a2111o_4 c405 (.A1(net28),
    .A2(net208),
    .B1(net105),
    .C1(net958),
    .D1(net124),
    .X(net211));
 sky130_fd_sc_hd__and3_2 c406 (.A(net207),
    .B(net206),
    .C(net958),
    .X(net212));
 sky130_fd_sc_hd__and3_4 c407 (.A(net767),
    .B(net111),
    .C(net209),
    .X(net213));
 sky130_fd_sc_hd__and3_1 c408 (.A(net212),
    .B(net637),
    .C(net213),
    .X(net214));
 sky130_fd_sc_hd__and2_2 c409 (.A(net886),
    .B(net958),
    .X(net215));
 sky130_fd_sc_hd__mux4_2 c410 (.A0(net109),
    .A1(net628),
    .A2(net112),
    .A3(net211),
    .S0(net833),
    .S1(net958),
    .X(net216));
 sky130_fd_sc_hd__mux4_2 c411 (.A0(net631),
    .A1(net27),
    .A2(net206),
    .A3(net213),
    .S0(net821),
    .S1(net116),
    .X(net217));
 sky130_fd_sc_hd__mux4_2 c412 (.A0(net210),
    .A1(net679),
    .A2(net213),
    .A3(net958),
    .S0(net123),
    .S1(net114),
    .X(net727));
 sky130_fd_sc_hd__and3_1 c413 (.A(net120),
    .B(net958),
    .C(net213),
    .X(net218));
 sky130_fd_sc_hd__and3_1 c414 (.A(net217),
    .B(net19),
    .C(net211),
    .X(net219));
 sky130_fd_sc_hd__and3_4 c415 (.A(net213),
    .B(net210),
    .C(net214),
    .X(net220));
 sky130_fd_sc_hd__and3_1 c416 (.A(net219),
    .B(net220),
    .C(net106),
    .X(net221));
 sky130_fd_sc_hd__mux4_2 c417 (.A0(net214),
    .A1(net109),
    .A2(net958),
    .A3(net221),
    .S0(net220),
    .S1(net211),
    .X(net222));
 sky130_fd_sc_hd__and3_1 c418 (.A(net134),
    .B(net135),
    .C(net823),
    .X(net223));
 sky130_fd_sc_hd__or4bb_4 c419 (.A(net988),
    .B(net137),
    .C_N(net44),
    .D_N(net124),
    .X(net224));
 sky130_fd_sc_hd__mux4_2 c420 (.A0(net628),
    .A1(net123),
    .A2(net144),
    .A3(net27),
    .S0(net807),
    .S1(net951),
    .X(net225));
 sky130_fd_sc_hd__or4bb_1 c421 (.A(net636),
    .B(net127),
    .C_N(net668),
    .D_N(net828),
    .X(net226));
 sky130_fd_sc_hd__and3_2 c422 (.A(net226),
    .B(net205),
    .C(net828),
    .X(net227));
 sky130_fd_sc_hd__and3_2 c423 (.A(net143),
    .B(net203),
    .C(net131),
    .X(net228));
 sky130_fd_sc_hd__or4bb_4 c424 (.A(net144),
    .B(net44),
    .C_N(net656),
    .D_N(net223),
    .X(net229));
 sky130_fd_sc_hd__and3_1 c425 (.A(net223),
    .B(net222),
    .C(net208),
    .X(net230));
 sky130_fd_sc_hd__and3_1 c426 (.A(net44),
    .B(net651),
    .C(net127),
    .X(net231));
 sky130_fd_sc_hd__and3_2 c427 (.A(net690),
    .B(net230),
    .C(net229),
    .X(net232));
 sky130_fd_sc_hd__and3_1 c428 (.A(net656),
    .B(net821),
    .C(net215),
    .X(net233));
 sky130_fd_sc_hd__buf_1 c429 (.A(net569),
    .X(net234));
 sky130_fd_sc_hd__or4bb_1 c430 (.A(net232),
    .B(net135),
    .C_N(net123),
    .D_N(net233),
    .X(net235));
 sky130_fd_sc_hd__and3_4 c431 (.A(net234),
    .B(net230),
    .C(net130),
    .X(net236));
 sky130_fd_sc_hd__and3_2 c432 (.A(net659),
    .B(net125),
    .C(net227),
    .X(net237));
 sky130_fd_sc_hd__and3_1 c433 (.A(net32),
    .B(net228),
    .C(net886),
    .X(net238));
 sky130_fd_sc_hd__and3_1 c434 (.A(net20),
    .B(net134),
    .C(net626),
    .X(net239));
 sky130_fd_sc_hd__mux4_1 c435 (.A0(net227),
    .A1(net212),
    .A2(net220),
    .A3(net229),
    .S0(net234),
    .S1(net237),
    .X(net240));
 sky130_fd_sc_hd__or4bb_1 c436 (.A(net130),
    .B(net637),
    .C_N(net240),
    .D_N(net238),
    .X(net241));
 sky130_fd_sc_hd__or4bb_2 c437 (.A(net231),
    .B(net205),
    .C_N(net958),
    .D_N(net42),
    .X(net242));
 sky130_fd_sc_hd__and3_2 c438 (.A(net144),
    .B(net731),
    .C(net839),
    .X(net243));
 sky130_fd_sc_hd__or4bb_1 c439 (.A(net140),
    .B(net243),
    .C_N(net809),
    .D_N(net838),
    .X(net244));
 sky130_fd_sc_hd__a2111o_1 c440 (.A1(net231),
    .A2(net656),
    .B1(net828),
    .C1(net119),
    .D1(net242),
    .X(net245));
 sky130_fd_sc_hd__and3_1 c441 (.A(net641),
    .B(net42),
    .C(net763),
    .X(net246));
 sky130_fd_sc_hd__and3_2 c442 (.A(net154),
    .B(net150),
    .C(net59),
    .X(net247));
 sky130_fd_sc_hd__buf_1 c443 (.A(net839),
    .X(net248));
 sky130_fd_sc_hd__a2111o_2 c444 (.A1(net226),
    .A2(net671),
    .B1(net248),
    .C1(net142),
    .D1(net42),
    .X(net249));
 sky130_fd_sc_hd__clkbuf_1 c445 (.A(net839),
    .X(net250));
 sky130_fd_sc_hd__and3_2 c446 (.A(net925),
    .B(net123),
    .C(net767),
    .X(net737));
 sky130_fd_sc_hd__and3_1 c447 (.A(net685),
    .B(net672),
    .C(net683),
    .X(net251));
 sky130_fd_sc_hd__and3_1 c448 (.A(net45),
    .B(net236),
    .C(net874),
    .X(net252));
 sky130_fd_sc_hd__mux4_1 c449 (.A0(net240),
    .A1(net239),
    .A2(net150),
    .A3(net59),
    .S0(net151),
    .S1(clknet_1_0__leaf_net799),
    .X(net253));
 sky130_fd_sc_hd__and3_1 c450 (.A(net246),
    .B(net149),
    .C(net220),
    .X(net254));
 sky130_fd_sc_hd__a2111o_1 c451 (.A1(net248),
    .A2(net247),
    .B1(net683),
    .C1(net252),
    .D1(clknet_1_0__leaf_net799),
    .X(net255));
 sky130_fd_sc_hd__a2111o_1 c452 (.A1(net659),
    .A2(net248),
    .B1(net814),
    .C1(net874),
    .D1(clknet_1_0__leaf_net162),
    .X(net256));
 sky130_fd_sc_hd__and3_1 c453 (.A(net249),
    .B(net976),
    .C(net132),
    .X(net257));
 sky130_fd_sc_hd__mux4_1 c454 (.A0(net251),
    .A1(net247),
    .A2(net257),
    .A3(net245),
    .S0(net151),
    .S1(net603),
    .X(net258));
 sky130_fd_sc_hd__mux4_2 c455 (.A0(net245),
    .A1(net56),
    .A2(net151),
    .A3(net668),
    .S0(net139),
    .S1(net838),
    .X(net259));
 sky130_fd_sc_hd__or4bb_2 c456 (.A(net257),
    .B(net251),
    .C_N(net259),
    .D_N(net878),
    .X(net260));
 sky130_fd_sc_hd__mux4_2 c457 (.A0(net147),
    .A1(net40),
    .A2(net47),
    .A3(net757),
    .S0(net259),
    .S1(net603),
    .X(net261));
 sky130_fd_sc_hd__buf_1 c458 (.A(net604),
    .X(net262));
 sky130_fd_sc_hd__and3_1 c459 (.A(net262),
    .B(net664),
    .C(net237),
    .X(net263));
 sky130_fd_sc_hd__mux4_1 c460 (.A0(net259),
    .A1(net260),
    .A2(net246),
    .A3(net263),
    .S0(net261),
    .S1(net770),
    .X(net264));
 sky130_fd_sc_hd__mux4_2 c461 (.A0(net263),
    .A1(net805),
    .A2(net156),
    .A3(net261),
    .S0(net249),
    .S1(net248),
    .X(net265));
 sky130_fd_sc_hd__or4bb_2 c462 (.A(net239),
    .B(net245),
    .C_N(net254),
    .D_N(net829),
    .X(net266));
 sky130_fd_sc_hd__a2111o_1 c463 (.A1(net979),
    .A2(net262),
    .B1(net770),
    .C1(net681),
    .D1(net603),
    .X(net267));
 sky130_fd_sc_hd__a2111o_1 c464 (.A1(net650),
    .A2(net705),
    .B1(net67),
    .C1(net734),
    .D1(clknet_1_0__leaf_net799),
    .X(net268));
 sky130_fd_sc_hd__a2111o_1 c465 (.A1(net51),
    .A2(net220),
    .B1(clknet_1_0__leaf_net162),
    .C1(clknet_1_0__leaf_net268),
    .D1(net232),
    .X(net269));
 sky130_fd_sc_hd__a2111o_2 c466 (.A1(net167),
    .A2(net262),
    .B1(net921),
    .C1(net145),
    .D1(net734),
    .X(net270));
 sky130_fd_sc_hd__a2111o_2 c467 (.A1(net267),
    .A2(net805),
    .B1(net65),
    .C1(net707),
    .D1(net603),
    .X(net271));
 sky130_fd_sc_hd__mux4_1 c468 (.A0(net67),
    .A1(net250),
    .A2(net770),
    .A3(net810),
    .S0(net843),
    .S1(net829),
    .X(net272));
 sky130_fd_sc_hd__mux4_1 c469 (.A0(net149),
    .A1(net110),
    .A2(net683),
    .A3(net229),
    .S0(net239),
    .S1(net270),
    .X(net273));
 sky130_fd_sc_hd__or4bb_1 c470 (.A(net150),
    .B(net271),
    .C_N(net262),
    .D_N(net68),
    .X(net274));
 sky130_fd_sc_hd__mux4_1 c471 (.A0(net208),
    .A1(net762),
    .A2(net749),
    .A3(net150),
    .S0(net847),
    .S1(net828),
    .X(net275));
 sky130_fd_sc_hd__a2111o_1 c472 (.A1(net229),
    .A2(net271),
    .B1(net254),
    .C1(net677),
    .D1(clknet_1_0__leaf_net178),
    .X(net276));
 sky130_fd_sc_hd__mux4_1 c473 (.A0(net156),
    .A1(net51),
    .A2(net67),
    .A3(clknet_1_1__leaf_net178),
    .S0(net805),
    .S1(net169),
    .X(net277));
 sky130_fd_sc_hd__mux4_1 c474 (.A0(net254),
    .A1(net628),
    .A2(net54),
    .A3(net810),
    .S0(net151),
    .S1(net679),
    .X(net278));
 sky130_fd_sc_hd__mux4_1 c475 (.A0(net119),
    .A1(net808),
    .A2(net757),
    .A3(net272),
    .S0(net229),
    .S1(net839),
    .X(net279));
 sky130_fd_sc_hd__a2111o_1 c476 (.A1(net279),
    .A2(net49),
    .B1(net273),
    .C1(net757),
    .D1(net265),
    .X(net280));
 sky130_fd_sc_hd__a2111o_1 c477 (.A1(net707),
    .A2(net229),
    .B1(net642),
    .C1(net840),
    .D1(net839),
    .X(net736));
 sky130_fd_sc_hd__a2111o_1 c478 (.A1(net688),
    .A2(net677),
    .B1(net707),
    .C1(clknet_1_1__leaf_net277),
    .D1(net829),
    .X(net281));
 sky130_fd_sc_hd__mux4_1 c479 (.A0(clknet_1_0__leaf_net281),
    .A1(net112),
    .A2(net42),
    .A3(net239),
    .S0(net66),
    .S1(net271),
    .X(net282));
 sky130_fd_sc_hd__mux4_1 c480 (.A0(net705),
    .A1(net274),
    .A2(net271),
    .A3(net81),
    .S0(clknet_1_1__leaf_net281),
    .S1(net839),
    .X(net283));
 sky130_fd_sc_hd__mux4_1 c481 (.A0(clknet_1_0__leaf_net277),
    .A1(net278),
    .A2(net252),
    .A3(net274),
    .S0(net271),
    .S1(clknet_1_0__leaf_net281),
    .X(net284));
 sky130_fd_sc_hd__mux4_1 c482 (.A0(net691),
    .A1(net736),
    .A2(clknet_1_1__leaf_net282),
    .A3(net709),
    .S0(net592),
    .S1(net603),
    .X(net285));
 sky130_fd_sc_hd__mux4_1 c483 (.A0(net250),
    .A1(net37),
    .A2(net882),
    .A3(net77),
    .S0(net279),
    .S1(net819),
    .X(net286));
 sky130_fd_sc_hd__a2111o_1 c484 (.A1(net270),
    .A2(clknet_1_1__leaf_net200),
    .B1(net47),
    .C1(net685),
    .D1(net804),
    .X(net287));
 sky130_fd_sc_hd__mux4_1 c485 (.A0(net4),
    .A1(net713),
    .A2(net755),
    .A3(net722),
    .S0(net738),
    .S1(net629),
    .X(net288));
 sky130_fd_sc_hd__mux4_2 c486 (.A0(net700),
    .A1(net642),
    .A2(net816),
    .A3(net639),
    .S0(net804),
    .S1(net603),
    .X(net764));
 sky130_fd_sc_hd__mux4_1 c487 (.A0(net220),
    .A1(net877),
    .A2(net699),
    .A3(net763),
    .S0(net817),
    .S1(clknet_1_1__leaf_net799),
    .X(net289));
 sky130_fd_sc_hd__mux4_1 c488 (.A0(net95),
    .A1(net90),
    .A2(net189),
    .A3(net220),
    .S0(net693),
    .S1(net811),
    .X(net290));
 sky130_fd_sc_hd__mux4_1 c489 (.A0(net151),
    .A1(net260),
    .A2(net201),
    .A3(net749),
    .S0(net816),
    .S1(net649),
    .X(net291));
 sky130_fd_sc_hd__mux4_1 c490 (.A0(net721),
    .A1(net631),
    .A2(net247),
    .A3(clknet_1_0__leaf_net289),
    .S0(net811),
    .S1(net819),
    .X(net292));
 sky130_fd_sc_hd__mux4_2 c491 (.A0(net147),
    .A1(net66),
    .A2(net758),
    .A3(net65),
    .S0(net677),
    .S1(clknet_1_1__leaf_net766),
    .X(net293));
 sky130_fd_sc_hd__mux4_1 c492 (.A0(net47),
    .A1(net65),
    .A2(net674),
    .A3(net754),
    .S0(net762),
    .S1(net66),
    .X(net745));
 sky130_fd_sc_hd__mux4_1 c493 (.A0(clknet_1_0__leaf_net282),
    .A1(net764),
    .A2(net765),
    .A3(net690),
    .S0(net757),
    .S1(net746),
    .X(net294));
 sky130_fd_sc_hd__mux4_1 c494 (.A0(clknet_1_0__leaf_net289),
    .A1(net183),
    .A2(net270),
    .A3(net114),
    .S0(net151),
    .S1(clknet_1_1__leaf_net799),
    .X(net295));
 sky130_fd_sc_hd__mux4_1 c495 (.A0(net876),
    .A1(net49),
    .A2(net270),
    .A3(net824),
    .S0(net592),
    .S1(net612),
    .X(net296));
 sky130_fd_sc_hd__a2111o_1 c496 (.A1(net649),
    .A2(net746),
    .B1(clknet_1_0__leaf_net276),
    .C1(clknet_1_0__leaf_net769),
    .D1(net613),
    .X(net297));
 sky130_fd_sc_hd__mux4_1 c497 (.A0(net639),
    .A1(net888),
    .A2(net224),
    .A3(net201),
    .S0(net853),
    .S1(net804),
    .X(net298));
 sky130_fd_sc_hd__mux4_1 c498 (.A0(net290),
    .A1(net653),
    .A2(net192),
    .A3(net270),
    .S0(net734),
    .S1(net819),
    .X(net299));
 sky130_fd_sc_hd__mux4_1 c499 (.A0(net677),
    .A1(net298),
    .A2(net270),
    .A3(net750),
    .S0(clknet_1_0__leaf_net295),
    .S1(net829),
    .X(net300));
 sky130_fd_sc_hd__mux4_1 c500 (.A0(net292),
    .A1(net764),
    .A2(net98),
    .A3(net744),
    .S0(net201),
    .S1(net836),
    .X(net301));
 sky130_fd_sc_hd__mux4_2 c501 (.A0(net119),
    .A1(net296),
    .A2(net755),
    .A3(net812),
    .S0(net847),
    .S1(net877),
    .X(net302));
 sky130_fd_sc_hd__mux4_1 c502 (.A0(net56),
    .A1(net754),
    .A2(clknet_1_0__leaf_net300),
    .A3(clknet_1_0__leaf_net198),
    .S0(net173),
    .S1(net600),
    .X(net303));
 sky130_fd_sc_hd__a2111o_1 c503 (.A1(net183),
    .A2(clknet_1_1__leaf_net300),
    .B1(clknet_1_0__leaf_net301),
    .C1(net194),
    .D1(net819),
    .X(net304));
 sky130_fd_sc_hd__mux4_1 c504 (.A0(net674),
    .A1(net626),
    .A2(clknet_1_0__leaf_net301),
    .A3(net672),
    .S0(net649),
    .S1(clknet_1_0__leaf_net289),
    .X(net305));
 sky130_fd_sc_hd__mux4_1 c505 (.A0(net299),
    .A1(net717),
    .A2(clknet_1_0__leaf_net305),
    .A3(net816),
    .S0(clknet_1_0__leaf_net198),
    .S1(net600),
    .X(net306));
 sky130_fd_sc_hd__and3_4 c528 (.A(net211),
    .B(net111),
    .C(net634),
    .X(net307));
 sky130_fd_sc_hd__and2_1 c529 (.A(net121),
    .B(net111),
    .X(net308));
 sky130_fd_sc_hd__and2_4 c530 (.A(net848),
    .B(net307),
    .X(net309));
 sky130_fd_sc_hd__and2_2 c531 (.A(net17),
    .B(net637),
    .X(net310));
 sky130_fd_sc_hd__or4bb_4 c532 (.A(net211),
    .B(net848),
    .C_N(net210),
    .D_N(net310),
    .X(net311));
 sky130_fd_sc_hd__mux4_2 c533 (.A0(net213),
    .A1(net309),
    .A2(net307),
    .A3(net121),
    .S0(net634),
    .S1(net806),
    .X(net312));
 sky130_fd_sc_hd__and2_1 c534 (.A(net309),
    .B(net218),
    .X(net313));
 sky130_fd_sc_hd__and2_4 c535 (.A(net896),
    .B(net310),
    .X(net314));
 sky130_fd_sc_hd__and2_1 c536 (.A(net204),
    .B(net897),
    .X(net315));
 sky130_fd_sc_hd__or4bb_4 c537 (.A(net221),
    .B(net761),
    .C_N(net21),
    .D_N(net823),
    .X(net316));
 sky130_fd_sc_hd__or4bb_4 c538 (.A(net206),
    .B(net21),
    .C_N(net313),
    .D_N(net312),
    .X(net317));
 sky130_fd_sc_hd__and2_2 c539 (.A(net833),
    .B(net309),
    .X(net318));
 sky130_fd_sc_hd__and2_2 c540 (.A(net898),
    .B(net315),
    .X(net726));
 sky130_fd_sc_hd__and3_4 c541 (.A(net316),
    .B(net207),
    .C(net206),
    .X(net319));
 sky130_fd_sc_hd__and2_0 c542 (.A(net105),
    .B(net124),
    .X(net320));
 sky130_fd_sc_hd__and3_1 c543 (.A(net317),
    .B(net314),
    .C(net806),
    .X(net321));
 sky130_fd_sc_hd__mux4_2 c544 (.A0(net319),
    .A1(net307),
    .A2(net318),
    .A3(net815),
    .S0(net311),
    .S1(net668),
    .X(net322));
 sky130_fd_sc_hd__or4bb_1 c545 (.A(net314),
    .B(net896),
    .C_N(net123),
    .D_N(net964),
    .X(net323));
 sky130_fd_sc_hd__or4bb_2 c546 (.A(net207),
    .B(net679),
    .C_N(net320),
    .D_N(net313),
    .X(net324));
 sky130_fd_sc_hd__mux4_2 c547 (.A0(net321),
    .A1(net313),
    .A2(net324),
    .A3(net209),
    .S0(net316),
    .S1(net806),
    .X(net325));
 sky130_fd_sc_hd__a2111o_2 c548 (.A1(net111),
    .A2(net323),
    .B1(net894),
    .C1(net215),
    .D1(net314),
    .X(net326));
 sky130_fd_sc_hd__or4bb_1 c549 (.A(net326),
    .B(net316),
    .C_N(net213),
    .D_N(net325),
    .X(net327));
 sky130_fd_sc_hd__a2111o_4 c550 (.A1(net315),
    .A2(net884),
    .B1(net314),
    .C1(net625),
    .D1(net838),
    .X(net723));
 sky130_fd_sc_hd__a2111o_4 c551 (.A1(net325),
    .A2(net950),
    .B1(net900),
    .C1(net723),
    .D1(net322),
    .X(net752));
 sky130_fd_sc_hd__or4bb_4 c552 (.A(net661),
    .B(net30),
    .C_N(net886),
    .D_N(net862),
    .X(net328));
 sky130_fd_sc_hd__and3_4 c553 (.A(net328),
    .B(net815),
    .C(net891),
    .X(net329));
 sky130_fd_sc_hd__and3_1 c554 (.A(net238),
    .B(net43),
    .C(net818),
    .X(net330));
 sky130_fd_sc_hd__or4bb_1 c555 (.A(net321),
    .B(net723),
    .C_N(net327),
    .D_N(net901),
    .X(net331));
 sky130_fd_sc_hd__a2111o_1 c556 (.A1(net135),
    .A2(net232),
    .B1(net121),
    .C1(net952),
    .D1(net227),
    .X(net332));
 sky130_fd_sc_hd__buf_1 c557 (.A(net562),
    .X(net333));
 sky130_fd_sc_hd__or4bb_4 c558 (.A(net333),
    .B(net137),
    .C_N(net225),
    .D_N(net823),
    .X(net334));
 sky130_fd_sc_hd__clkbuf_1 c559 (.A(net562),
    .X(net335));
 sky130_fd_sc_hd__or4bb_4 c560 (.A(net230),
    .B(net752),
    .C_N(net807),
    .D_N(net823),
    .X(net336));
 sky130_fd_sc_hd__or4bb_1 c561 (.A(net335),
    .B(net25),
    .C_N(net806),
    .D_N(net573),
    .X(net337));
 sky130_fd_sc_hd__or4bb_4 c562 (.A(net221),
    .B(net336),
    .C_N(net328),
    .D_N(net839),
    .X(net338));
 sky130_fd_sc_hd__buf_1 c563 (.A(net569),
    .X(net339));
 sky130_fd_sc_hd__or4bb_1 c564 (.A(net339),
    .B(net318),
    .C_N(net43),
    .D_N(net107),
    .X(net340));
 sky130_fd_sc_hd__mux4_2 c565 (.A0(net337),
    .A1(net314),
    .A2(net131),
    .A3(net340),
    .S0(net339),
    .S1(net660),
    .X(net341));
 sky130_fd_sc_hd__mux4_2 c566 (.A0(net203),
    .A1(net950),
    .A2(net228),
    .A3(net25),
    .S0(net818),
    .S1(net333),
    .X(net747));
 sky130_fd_sc_hd__sdfbbn_1 c567 (.CLK_N(clknet_2_2__leaf_clk),
    .D(net313),
    .RESET_B(net338),
    .SCD(net747),
    .SCE(net341),
    .SET_B(net657),
    .Q(net343),
    .Q_N(net342));
 sky130_fd_sc_hd__or4bb_1 c568 (.A(net915),
    .B(net336),
    .C_N(net804),
    .D_N(net857),
    .X(net344));
 sky130_fd_sc_hd__mux4_1 c569 (.A0(net655),
    .A1(net747),
    .A2(net330),
    .A3(net752),
    .S0(net236),
    .S1(net574),
    .X(net345));
 sky130_fd_sc_hd__a2111o_4 c570 (.A1(net329),
    .A2(net804),
    .B1(net337),
    .C1(net342),
    .D1(net574),
    .X(net346));
 sky130_fd_sc_hd__mux4_2 c571 (.A0(net205),
    .A1(net338),
    .A2(net342),
    .A3(net330),
    .S0(net747),
    .S1(net574),
    .X(net347));
 sky130_fd_sc_hd__and3_1 c572 (.A(net340),
    .B(net860),
    .C(net645),
    .X(net348));
 sky130_fd_sc_hd__a2111o_1 c573 (.A1(net260),
    .A2(net844),
    .B1(net908),
    .C1(net927),
    .D1(net31),
    .X(net349));
 sky130_fd_sc_hd__a2111o_1 c574 (.A1(net25),
    .A2(net859),
    .B1(clknet_1_0__leaf_net162),
    .C1(net807),
    .D1(net833),
    .X(net350));
 sky130_fd_sc_hd__and3_1 c575 (.A(net857),
    .B(net672),
    .C(net671),
    .X(net351));
 sky130_fd_sc_hd__mux4_1 c576 (.A0(net236),
    .A1(net146),
    .A2(net737),
    .A3(net42),
    .S0(net265),
    .S1(clknet_1_1__leaf_net161),
    .X(net352));
 sky130_fd_sc_hd__and3_2 c577 (.A(net251),
    .B(net569),
    .C(net743),
    .X(net353));
 sky130_fd_sc_hd__and3_2 c578 (.A(net944),
    .B(net846),
    .C(net807),
    .X(net354));
 sky130_fd_sc_hd__mux4_1 c579 (.A0(net330),
    .A1(net341),
    .A2(net846),
    .A3(net679),
    .S0(net971),
    .S1(net569),
    .X(net355));
 sky130_fd_sc_hd__and3_1 c580 (.A(net261),
    .B(net955),
    .C(net236),
    .X(net356));
 sky130_fd_sc_hd__a2111o_1 c581 (.A1(net335),
    .A2(net25),
    .B1(net833),
    .C1(net242),
    .D1(net353),
    .X(net357));
 sky130_fd_sc_hd__or4bb_1 c582 (.A(net237),
    .B(net357),
    .C_N(net807),
    .D_N(net43),
    .X(net358));
 sky130_fd_sc_hd__and3_1 c583 (.A(net139),
    .B(net341),
    .C(net743),
    .X(net359));
 sky130_fd_sc_hd__mux4_1 c584 (.A0(net679),
    .A1(net660),
    .A2(net830),
    .A3(net341),
    .S0(net815),
    .S1(net353),
    .X(net360));
 sky130_fd_sc_hd__or4bb_1 c585 (.A(net132),
    .B(net637),
    .C_N(net915),
    .D_N(net327),
    .X(net361));
 sky130_fd_sc_hd__a2111o_1 c586 (.A1(net356),
    .A2(net358),
    .B1(net334),
    .C1(net131),
    .D1(net357),
    .X(net362));
 sky130_fd_sc_hd__mux4_1 c587 (.A0(net360),
    .A1(net915),
    .A2(net343),
    .A3(net356),
    .S0(net650),
    .S1(net846),
    .X(net363));
 sky130_fd_sc_hd__a2111o_1 c588 (.A1(net327),
    .A2(net353),
    .B1(net237),
    .C1(net943),
    .D1(clknet_1_0__leaf_net162),
    .X(net364));
 sky130_fd_sc_hd__mux4_1 c589 (.A0(clknet_1_1__leaf_net161),
    .A1(net353),
    .A2(net341),
    .A3(net354),
    .S0(net807),
    .S1(net618),
    .X(net365));
 sky130_fd_sc_hd__and3_1 c590 (.A(net359),
    .B(net318),
    .C(clknet_1_1__leaf_net614),
    .X(net366));
 sky130_fd_sc_hd__and3_1 c591 (.A(net366),
    .B(net257),
    .C(net359),
    .X(net367));
 sky130_fd_sc_hd__mux4_2 c592 (.A0(net324),
    .A1(net353),
    .A2(net227),
    .A3(net236),
    .S0(net597),
    .S1(net836),
    .X(net368));
 sky130_fd_sc_hd__a2111o_1 c593 (.A1(net152),
    .A2(net353),
    .B1(clknet_1_0__leaf_net367),
    .C1(net849),
    .D1(net836),
    .X(net369));
 sky130_fd_sc_hd__mux4_1 c594 (.A0(net81),
    .A1(net692),
    .A2(net902),
    .A3(net341),
    .S0(net954),
    .S1(clknet_1_0__leaf_net799),
    .X(net370));
 sky130_fd_sc_hd__mux4_2 c595 (.A0(net650),
    .A1(net902),
    .A2(net737),
    .A3(net890),
    .S0(net22),
    .S1(net888),
    .X(net751));
 sky130_fd_sc_hd__mux4_1 c596 (.A0(net169),
    .A1(net129),
    .A2(net847),
    .A3(net844),
    .S0(net734),
    .S1(net604),
    .X(net371));
 sky130_fd_sc_hd__a2111o_1 c597 (.A1(net645),
    .A2(net42),
    .B1(net224),
    .C1(net139),
    .D1(net820),
    .X(net372));
 sky130_fd_sc_hd__a2111o_1 c598 (.A1(net271),
    .A2(net267),
    .B1(net818),
    .C1(net850),
    .D1(net945),
    .X(net373));
 sky130_fd_sc_hd__a2111o_1 c599 (.A1(clknet_1_1__leaf_net268),
    .A2(net916),
    .B1(net749),
    .C1(net271),
    .D1(net667),
    .X(net374));
 sky130_fd_sc_hd__mux4_1 c600 (.A0(clknet_1_1__leaf_net178),
    .A1(net169),
    .A2(net59),
    .A3(net341),
    .S0(net597),
    .S1(net616),
    .X(net375));
 sky130_fd_sc_hd__a2111o_1 c601 (.A1(clknet_1_1__leaf_net375),
    .A2(net77),
    .B1(net373),
    .C1(net351),
    .D1(net838),
    .X(net376));
 sky130_fd_sc_hd__mux4_1 c602 (.A0(net30),
    .A1(net232),
    .A2(net907),
    .A3(net888),
    .S0(net733),
    .S1(net743),
    .X(net377));
 sky130_fd_sc_hd__a2111o_1 c603 (.A1(net371),
    .A2(net326),
    .B1(net22),
    .C1(net909),
    .D1(net859),
    .X(net378));
 sky130_fd_sc_hd__mux4_1 c604 (.A0(net679),
    .A1(net232),
    .A2(net906),
    .A3(net851),
    .S0(net372),
    .S1(net972),
    .X(net379));
 sky130_fd_sc_hd__mux4_1 c605 (.A0(net374),
    .A1(net334),
    .A2(net698),
    .A3(net351),
    .S0(net326),
    .S1(clknet_1_0__leaf_net799),
    .X(net380));
 sky130_fd_sc_hd__mux4_1 c606 (.A0(net252),
    .A1(net846),
    .A2(net110),
    .A3(net709),
    .S0(net681),
    .S1(net841),
    .X(net381));
 sky130_fd_sc_hd__mux4_1 c607 (.A0(net685),
    .A1(net353),
    .A2(net650),
    .A3(net824),
    .S0(net573),
    .S1(net759),
    .X(net382));
 sky130_fd_sc_hd__mux4_2 c608 (.A0(net341),
    .A1(net275),
    .A2(net751),
    .A3(net846),
    .S0(net905),
    .S1(net679),
    .X(net383));
 sky130_fd_sc_hd__mux4_1 c609 (.A0(net629),
    .A1(net382),
    .A2(net372),
    .A3(net849),
    .S0(net922),
    .S1(net743),
    .X(net384));
 sky130_fd_sc_hd__mux4_1 c610 (.A0(net895),
    .A1(net645),
    .A2(net275),
    .A3(net114),
    .S0(clknet_1_0__leaf_net255),
    .S1(net382),
    .X(net385));
 sky130_fd_sc_hd__mux4_1 c611 (.A0(net384),
    .A1(net311),
    .A2(net868),
    .A3(clknet_1_0__leaf_net375),
    .S0(clknet_1_1__leaf_net162),
    .S1(net602),
    .X(net386));
 sky130_fd_sc_hd__a2111o_4 c612 (.A1(net908),
    .A2(net683),
    .B1(net738),
    .C1(net692),
    .D1(net608),
    .X(net387));
 sky130_fd_sc_hd__mux4_1 c613 (.A0(net81),
    .A1(net709),
    .A2(net54),
    .A3(net691),
    .S0(net387),
    .S1(net608),
    .X(net388));
 sky130_fd_sc_hd__mux4_1 c614 (.A0(net385),
    .A1(net372),
    .A2(net224),
    .A3(net387),
    .S0(net625),
    .S1(net629),
    .X(net389));
 sky130_fd_sc_hd__mux4_1 c615 (.A0(net388),
    .A1(net387),
    .A2(net114),
    .A3(net726),
    .S0(net759),
    .S1(clknet_1_1__leaf_net614),
    .X(net793));
 sky130_fd_sc_hd__mux4_1 c616 (.A0(net387),
    .A1(net189),
    .A2(net813),
    .A3(net843),
    .S0(net749),
    .S1(net820),
    .X(net739));
 sky130_fd_sc_hd__mux4_1 c617 (.A0(net272),
    .A1(net804),
    .A2(net805),
    .A3(net629),
    .S0(net22),
    .S1(net836),
    .X(net390));
 sky130_fd_sc_hd__mux4_1 c618 (.A0(net247),
    .A1(clknet_1_1__leaf_net305),
    .A2(net685),
    .A3(net173),
    .S0(net836),
    .S1(clknet_1_1__leaf_net799),
    .X(net391));
 sky130_fd_sc_hd__mux4_1 c619 (.A0(clknet_1_0__leaf_net295),
    .A1(net191),
    .A2(net73),
    .A3(clknet_1_1__leaf_net301),
    .S0(net830),
    .S1(net592),
    .X(net392));
 sky130_fd_sc_hd__mux4_1 c620 (.A0(net351),
    .A1(net668),
    .A2(net699),
    .A3(clknet_1_1__leaf_net198),
    .S0(net722),
    .S1(net612),
    .X(net393));
 sky130_fd_sc_hd__mux4_1 c621 (.A0(net381),
    .A1(net348),
    .A2(net265),
    .A3(clknet_1_1__leaf_net289),
    .S0(net805),
    .S1(net841),
    .X(net394));
 sky130_fd_sc_hd__mux4_1 c622 (.A0(net672),
    .A1(net201),
    .A2(net702),
    .A3(net843),
    .S0(net759),
    .S1(net612),
    .X(net395));
 sky130_fd_sc_hd__mux4_1 c623 (.A0(net224),
    .A1(net394),
    .A2(net182),
    .A3(net953),
    .S0(net737),
    .S1(clknet_1_0__leaf_net793),
    .X(net396));
 sky130_fd_sc_hd__mux4_1 c624 (.A0(net196),
    .A1(net182),
    .A2(net260),
    .A3(net224),
    .S0(net608),
    .S1(net613),
    .X(net397));
 sky130_fd_sc_hd__mux4_1 c625 (.A0(net378),
    .A1(net643),
    .A2(clknet_1_1__leaf_net295),
    .A3(net667),
    .S0(net816),
    .S1(net593),
    .X(net398));
 sky130_fd_sc_hd__mux4_1 c626 (.A0(clknet_1_1__leaf_net276),
    .A1(net395),
    .A2(net651),
    .A3(net804),
    .S0(net191),
    .S1(net820),
    .X(net399));
 sky130_fd_sc_hd__mux4_1 c627 (.A0(net145),
    .A1(net54),
    .A2(clknet_1_0__leaf_net255),
    .A3(net625),
    .S0(net387),
    .S1(net620),
    .X(net741));
 sky130_fd_sc_hd__mux4_1 c628 (.A0(net685),
    .A1(net173),
    .A2(clknet_1_1__leaf_net295),
    .A3(net110),
    .S0(net847),
    .S1(net593),
    .X(net400));
 sky130_fd_sc_hd__a2111o_1 c629 (.A1(net201),
    .A2(net847),
    .B1(net354),
    .C1(net603),
    .D1(net621),
    .X(net401));
 sky130_fd_sc_hd__mux4_1 c630 (.A0(net390),
    .A1(net197),
    .A2(net804),
    .A3(net672),
    .S0(net812),
    .S1(net815),
    .X(net402));
 sky130_fd_sc_hd__mux4_1 c631 (.A0(net114),
    .A1(clknet_1_1__leaf_net289),
    .A2(net626),
    .A3(net593),
    .S0(net836),
    .S1(net620),
    .X(net403));
 sky130_fd_sc_hd__mux4_1 c632 (.A0(net651),
    .A1(net403),
    .A2(net197),
    .A3(net54),
    .S0(net387),
    .S1(clknet_1_0__leaf_net400),
    .X(net404));
 sky130_fd_sc_hd__mux4_2 c633 (.A0(net273),
    .A1(net395),
    .A2(net984),
    .A3(net351),
    .S0(net734),
    .S1(net612),
    .X(net405));
 sky130_fd_sc_hd__mux4_1 c634 (.A0(clknet_1_1__leaf_net198),
    .A1(net192),
    .A2(clknet_1_1__leaf_net289),
    .A3(net387),
    .S0(net837),
    .S1(net621),
    .X(net406));
 sky130_fd_sc_hd__mux4_1 c635 (.A0(net84),
    .A1(net683),
    .A2(net746),
    .A3(net759),
    .S0(net611),
    .S1(clknet_1_1__leaf_net615),
    .X(net407));
 sky130_fd_sc_hd__mux4_1 c636 (.A0(net98),
    .A1(clknet_1_1__leaf_net301),
    .A2(net668),
    .A3(net685),
    .S0(net844),
    .S1(net611),
    .X(net408));
 sky130_fd_sc_hd__mux4_2 c637 (.A0(net383),
    .A1(net408),
    .A2(net984),
    .A3(net593),
    .S0(clknet_1_1__leaf_net615),
    .S1(net621),
    .X(net409));
 sky130_fd_sc_hd__or4bb_4 c660 (.A(net309),
    .B(net311),
    .C_N(net825),
    .D_N(net879),
    .X(net410));
 sky130_fd_sc_hd__and3_1 c661 (.A(net854),
    .B(net308),
    .C(net218),
    .X(net411));
 sky130_fd_sc_hd__a2111o_2 c662 (.A1(net885),
    .A2(net898),
    .B1(net928),
    .C1(net817),
    .D1(net807),
    .X(net412));
 sky130_fd_sc_hd__and2_1 c663 (.A(net214),
    .B(net323),
    .X(net413));
 sky130_fd_sc_hd__and2_0 c664 (.A(net209),
    .B(net726),
    .X(net414));
 sky130_fd_sc_hd__and3_2 c665 (.A(net411),
    .B(net932),
    .C(net817),
    .X(net415));
 sky130_fd_sc_hd__or4bb_2 c666 (.A(net931),
    .B(net21),
    .C_N(net212),
    .D_N(net855),
    .X(net416));
 sky130_fd_sc_hd__and3_1 c667 (.A(net123),
    .B(net308),
    .C(net413),
    .X(net417));
 sky130_fd_sc_hd__a2111o_1 c668 (.A1(net417),
    .A2(net410),
    .B1(net307),
    .C1(net864),
    .D1(net124),
    .X(net418));
 sky130_fd_sc_hd__a2111o_1 c669 (.A1(net323),
    .A2(net413),
    .B1(net863),
    .C1(net807),
    .D1(net930),
    .X(net419));
 sky130_fd_sc_hd__and3_1 c670 (.A(net210),
    .B(net413),
    .C(net843),
    .X(net420));
 sky130_fd_sc_hd__and3_1 c671 (.A(net418),
    .B(net821),
    .C(net825),
    .X(net421));
 sky130_fd_sc_hd__or4bb_1 c672 (.A(net21),
    .B(net738),
    .C_N(net420),
    .D_N(net880),
    .X(net422));
 sky130_fd_sc_hd__and3_1 c673 (.A(net420),
    .B(net418),
    .C(net865),
    .X(net423));
 sky130_fd_sc_hd__and3_2 c674 (.A(net880),
    .B(net124),
    .C(net416),
    .X(net724));
 sky130_fd_sc_hd__and3_2 c675 (.A(net413),
    .B(net724),
    .C(net420),
    .X(net424));
 sky130_fd_sc_hd__a2111o_1 c676 (.A1(net419),
    .A2(net880),
    .B1(net424),
    .C1(net423),
    .D1(net116),
    .X(net425));
 sky130_fd_sc_hd__sdfbbn_1 c677 (.CLK_N(clknet_2_2__leaf_clk),
    .D(net414),
    .RESET_B(net929),
    .SCD(net124),
    .SCE(net424),
    .SET_B(net418),
    .Q(net427),
    .Q_N(net426));
 sky130_fd_sc_hd__sdfbbp_1 c678 (.CLK(clknet_2_2__leaf_clk),
    .D(net116),
    .RESET_B(net308),
    .SCD(net424),
    .SCE(net415),
    .SET_B(net744),
    .Q(net429),
    .Q_N(net428));
 sky130_fd_sc_hd__a2111o_1 c679 (.A1(net421),
    .A2(net960),
    .B1(net218),
    .C1(net424),
    .D1(net885),
    .X(net430));
 sky130_fd_sc_hd__a2111o_1 c680 (.A1(net422),
    .A2(net424),
    .B1(net427),
    .C1(net116),
    .D1(net856),
    .X(net431));
 sky130_fd_sc_hd__mux4_1 c681 (.A0(net424),
    .A1(net428),
    .A2(net881),
    .A3(net899),
    .S0(net543),
    .S1(net571),
    .X(net432));
 sky130_fd_sc_hd__mux4_1 c682 (.A0(net625),
    .A1(net243),
    .A2(net310),
    .A3(net657),
    .S0(net412),
    .S1(net839),
    .X(net433));
 sky130_fd_sc_hd__or4bb_1 c683 (.A(net315),
    .B(net29),
    .C_N(net139),
    .D_N(net838),
    .X(net434));
 sky130_fd_sc_hd__or4bb_1 c684 (.A(net243),
    .B(net626),
    .C_N(net215),
    .D_N(net346),
    .X(net435));
 sky130_fd_sc_hd__or4bb_2 c685 (.A(net212),
    .B(net315),
    .C_N(net847),
    .D_N(net830),
    .X(net436));
 sky130_fd_sc_hd__a2111o_1 c686 (.A1(net137),
    .A2(net215),
    .B1(net724),
    .C1(net225),
    .D1(net571),
    .X(net437));
 sky130_fd_sc_hd__a2111o_1 c687 (.A1(net124),
    .A2(net411),
    .B1(net815),
    .C1(net123),
    .D1(net346),
    .X(net438));
 sky130_fd_sc_hd__or4bb_2 c688 (.A(net856),
    .B(net434),
    .C_N(net562),
    .D_N(net838),
    .X(net439));
 sky130_fd_sc_hd__or4bb_1 c689 (.A(net435),
    .B(net343),
    .C_N(net242),
    .D_N(net830),
    .X(net440));
 sky130_fd_sc_hd__and3_1 c690 (.A(net434),
    .B(net863),
    .C(net549),
    .X(net441));
 sky130_fd_sc_hd__mux4_1 c691 (.A0(net985),
    .A1(net412),
    .A2(net845),
    .A3(net543),
    .S0(net839),
    .S1(net609),
    .X(net442));
 sky130_fd_sc_hd__or4bb_1 c692 (.A(net308),
    .B(net427),
    .C_N(net656),
    .D_N(net660),
    .X(net443));
 sky130_fd_sc_hd__or4bb_1 c693 (.A(net441),
    .B(net883),
    .C_N(net426),
    .D_N(net830),
    .X(net444));
 sky130_fd_sc_hd__or4bb_1 c694 (.A(net423),
    .B(net871),
    .C_N(net978),
    .D_N(net562),
    .X(net445));
 sky130_fd_sc_hd__and3_1 c695 (.A(net311),
    .B(net807),
    .C(net872),
    .X(net446));
 sky130_fd_sc_hd__or4bb_1 c696 (.A(net434),
    .B(net744),
    .C_N(net342),
    .D_N(net435),
    .X(net447));
 sky130_fd_sc_hd__mux4_1 c697 (.A0(net442),
    .A1(net334),
    .A2(net412),
    .A3(net227),
    .S0(net212),
    .S1(net549),
    .X(net448));
 sky130_fd_sc_hd__or4bb_1 c698 (.A(net871),
    .B(net437),
    .C_N(net311),
    .D_N(net571),
    .X(net449));
 sky130_fd_sc_hd__mux4_1 c699 (.A0(net446),
    .A1(net139),
    .A2(net441),
    .A3(net571),
    .S0(net607),
    .S1(net609),
    .X(net450));
 sky130_fd_sc_hd__or4bb_4 c700 (.A(net427),
    .B(net139),
    .C_N(net548),
    .D_N(net571),
    .X(net451));
 sky130_fd_sc_hd__mux4_1 c701 (.A0(net444),
    .A1(net660),
    .A2(net816),
    .A3(net426),
    .S0(net976),
    .S1(net609),
    .X(net452));
 sky130_fd_sc_hd__or4bb_2 c702 (.A(net215),
    .B(net228),
    .C_N(net917),
    .D_N(net543),
    .X(net453));
 sky130_fd_sc_hd__mux4_1 c703 (.A0(net443),
    .A1(net453),
    .A2(net436),
    .A3(net415),
    .S0(net243),
    .S1(net608),
    .X(net454));
 sky130_fd_sc_hd__a2111o_1 c704 (.A1(net310),
    .A2(net22),
    .B1(net981),
    .C1(net249),
    .D1(net816),
    .X(net455));
 sky130_fd_sc_hd__sdfbbn_1 c705 (.CLK_N(clknet_2_2__leaf_clk),
    .D(net416),
    .RESET_B(net660),
    .SCD(net453),
    .SCE(net843),
    .SET_B(net959),
    .Q(net457),
    .Q_N(net456));
 sky130_fd_sc_hd__mux4_1 c706 (.A0(net242),
    .A1(net976),
    .A2(net311),
    .A3(net724),
    .S0(net368),
    .S1(net622),
    .X(net458));
 sky130_fd_sc_hd__mux4_1 c707 (.A0(net671),
    .A1(net314),
    .A2(net265),
    .A3(net227),
    .S0(net982),
    .S1(net805),
    .X(net459));
 sky130_fd_sc_hd__mux4_2 c708 (.A0(net148),
    .A1(net123),
    .A2(net456),
    .A3(net816),
    .S0(net837),
    .S1(net622),
    .X(net460));
 sky130_fd_sc_hd__a2111o_1 c709 (.A1(net933),
    .A2(net458),
    .B1(net415),
    .C1(net889),
    .D1(net544),
    .X(net461));
 sky130_fd_sc_hd__mux4_2 c710 (.A0(net438),
    .A1(net249),
    .A2(net451),
    .A3(net415),
    .S0(net228),
    .S1(net607),
    .X(net462));
 sky130_fd_sc_hd__mux4_2 c711 (.A0(net228),
    .A1(net131),
    .A2(net436),
    .A3(net846),
    .S0(net889),
    .S1(net626),
    .X(net463));
 sky130_fd_sc_hd__mux4_1 c712 (.A0(net807),
    .A1(net334),
    .A2(net974),
    .A3(net805),
    .S0(net845),
    .S1(net837),
    .X(net464));
 sky130_fd_sc_hd__a2111o_1 c713 (.A1(net368),
    .A2(net428),
    .B1(net148),
    .C1(net548),
    .D1(net611),
    .X(net465));
 sky130_fd_sc_hd__mux4_1 c714 (.A0(net465),
    .A1(net410),
    .A2(net216),
    .A3(net813),
    .S0(net314),
    .S1(net412),
    .X(net466));
 sky130_fd_sc_hd__a2111o_1 c715 (.A1(net357),
    .A2(net123),
    .B1(net429),
    .C1(net416),
    .D1(clknet_1_0__leaf_net367),
    .X(net467));
 sky130_fd_sc_hd__mux4_1 c716 (.A0(clknet_1_1__leaf_net367),
    .A1(net429),
    .A2(net671),
    .A3(net660),
    .S0(net846),
    .S1(clknet_1_0__leaf_net614),
    .X(net468));
 sky130_fd_sc_hd__a2111o_1 c717 (.A1(net926),
    .A2(net460),
    .B1(net428),
    .C1(net726),
    .D1(clknet_1_0__leaf_net615),
    .X(net469));
 sky130_fd_sc_hd__sdfbbn_1 c718 (.CLK_N(clknet_2_2__leaf_clk),
    .D(net334),
    .RESET_B(net821),
    .SCD(clknet_1_1__leaf_net162),
    .SCE(net457),
    .SET_B(net830),
    .Q(net471),
    .Q_N(net470));
 sky130_fd_sc_hd__mux4_1 c719 (.A0(net986),
    .A1(net469),
    .A2(net444),
    .A3(net470),
    .S0(net847),
    .S1(net656),
    .X(net472));
 sky130_fd_sc_hd__mux4_2 c720 (.A0(net889),
    .A1(net933),
    .A2(net465),
    .A3(net818),
    .S0(net847),
    .S1(clknet_1_0__leaf_net614),
    .X(net473));
 sky130_fd_sc_hd__a2111o_1 c721 (.A1(net471),
    .A2(net462),
    .B1(net660),
    .C1(net671),
    .D1(clknet_1_0__leaf_net614),
    .X(net474));
 sky130_fd_sc_hd__mux4_1 c722 (.A0(net412),
    .A1(net470),
    .A2(net926),
    .A3(net139),
    .S0(net743),
    .S1(clknet_1_0__leaf_net615),
    .X(net475));
 sky130_fd_sc_hd__mux4_1 c723 (.A0(net453),
    .A1(net227),
    .A2(net460),
    .A3(net415),
    .S0(net867),
    .S1(net433),
    .X(net476));
 sky130_fd_sc_hd__a2111o_1 c724 (.A1(net437),
    .A2(net452),
    .B1(net888),
    .C1(clknet_1_0__leaf_net473),
    .D1(clknet_1_0__leaf_net614),
    .X(net477));
 sky130_fd_sc_hd__mux4_1 c725 (.A0(net436),
    .A1(net471),
    .A2(net410),
    .A3(net605),
    .S0(net611),
    .S1(clknet_1_0__leaf_net614),
    .X(net729));
 sky130_fd_sc_hd__mux4_1 c726 (.A0(net318),
    .A1(net439),
    .A2(net845),
    .A3(net353),
    .S0(net451),
    .S1(net838),
    .X(net478));
 sky130_fd_sc_hd__mux4_1 c727 (.A0(clknet_1_0__leaf_net473),
    .A1(net37),
    .A2(net843),
    .A3(clknet_1_1__leaf_net162),
    .S0(net456),
    .S1(clknet_1_0__leaf_net615),
    .X(net479));
 sky130_fd_sc_hd__mux4_1 c728 (.A0(net455),
    .A1(net450),
    .A2(net892),
    .A3(net22),
    .S0(net609),
    .S1(net622),
    .X(net480));
 sky130_fd_sc_hd__mux4_1 c729 (.A0(net860),
    .A1(clknet_1_1__leaf_net475),
    .A2(net731),
    .A3(net22),
    .S0(net702),
    .S1(net759),
    .X(net481));
 sky130_fd_sc_hd__mux4_1 c730 (.A0(net410),
    .A1(net738),
    .A2(net870),
    .A3(net605),
    .S0(net609),
    .S1(net759),
    .X(net482));
 sky130_fd_sc_hd__mux4_1 c731 (.A0(net354),
    .A1(net173),
    .A2(net629),
    .A3(net544),
    .S0(net619),
    .S1(net622),
    .X(net483));
 sky130_fd_sc_hd__mux4_1 c732 (.A0(net139),
    .A1(net457),
    .A2(net59),
    .A3(net683),
    .S0(net667),
    .S1(net616),
    .X(net484));
 sky130_fd_sc_hd__mux4_1 c733 (.A0(net668),
    .A1(net805),
    .A2(net68),
    .A3(net845),
    .S0(net820),
    .S1(net623),
    .X(net785));
 sky130_fd_sc_hd__mux4_1 c734 (.A0(net484),
    .A1(net805),
    .A2(net641),
    .A3(net605),
    .S0(net618),
    .S1(net623),
    .X(net485));
 sky130_fd_sc_hd__mux4_1 c735 (.A0(net629),
    .A1(net40),
    .A2(net805),
    .A3(net738),
    .S0(net608),
    .S1(net623),
    .X(net486));
 sky130_fd_sc_hd__mux4_1 c736 (.A0(net665),
    .A1(net466),
    .A2(net460),
    .A3(net982),
    .S0(net544),
    .S1(net623),
    .X(net487));
 sky130_fd_sc_hd__mux4_1 c737 (.A0(net906),
    .A1(net457),
    .A2(clknet_1_1__leaf_net370),
    .A3(net815),
    .S0(net702),
    .S1(net838),
    .X(net488));
 sky130_fd_sc_hd__mux4_1 c738 (.A0(net668),
    .A1(net71),
    .A2(net667),
    .A3(net977),
    .S0(net485),
    .S1(net110),
    .X(net489));
 sky130_fd_sc_hd__mux4_1 c739 (.A0(net433),
    .A1(net59),
    .A2(net37),
    .A3(net439),
    .S0(net110),
    .S1(net460),
    .X(net490));
 sky130_fd_sc_hd__mux4_1 c740 (.A0(net415),
    .A1(net353),
    .A2(net478),
    .A3(net665),
    .S0(net456),
    .S1(net623),
    .X(net491));
 sky130_fd_sc_hd__mux4_1 c741 (.A0(net451),
    .A1(net486),
    .A2(net624),
    .A3(net71),
    .S0(net982),
    .S1(net606),
    .X(net492));
 sky130_fd_sc_hd__mux4_1 c742 (.A0(net129),
    .A1(net415),
    .A2(net410),
    .A3(net839),
    .S0(net607),
    .S1(net623),
    .X(net493));
 sky130_fd_sc_hd__mux4_1 c743 (.A0(net491),
    .A1(clknet_1_1__leaf_net162),
    .A2(net692),
    .A3(net439),
    .S0(net785),
    .S1(net451),
    .X(net494));
 sky130_fd_sc_hd__mux4_1 c744 (.A0(clknet_1_0__leaf_net475),
    .A1(net459),
    .A2(net173),
    .A3(clknet_1_1__leaf_net473),
    .S0(net40),
    .S1(net606),
    .X(net495));
 sky130_fd_sc_hd__mux4_1 c745 (.A0(clknet_1_1__leaf_net162),
    .A1(net266),
    .A2(net463),
    .A3(net656),
    .S0(net611),
    .S1(net617),
    .X(net496));
 sky130_fd_sc_hd__mux4_1 c746 (.A0(net866),
    .A1(net701),
    .A2(net439),
    .A3(clknet_1_0__leaf_net615),
    .S0(net617),
    .S1(net623),
    .X(net497));
 sky130_fd_sc_hd__mux4_1 c747 (.A0(net849),
    .A1(net497),
    .A2(net626),
    .A3(net616),
    .S0(net622),
    .S1(net623),
    .X(net498));
 sky130_fd_sc_hd__mux4_1 c748 (.A0(net373),
    .A1(net266),
    .A2(net393),
    .A3(net645),
    .S0(net641),
    .S1(net815),
    .X(net499));
 sky130_fd_sc_hd__mux4_2 c749 (.A0(net69),
    .A1(net406),
    .A2(net812),
    .A3(net629),
    .S0(net463),
    .S1(net613),
    .X(net500));
 sky130_fd_sc_hd__mux4_2 c750 (.A0(net489),
    .A1(net293),
    .A2(net482),
    .A3(net681),
    .S0(net602),
    .S1(net608),
    .X(net501));
 sky130_fd_sc_hd__mux4_1 c751 (.A0(net37),
    .A1(net701),
    .A2(net498),
    .A3(net500),
    .S0(net22),
    .S1(net731),
    .X(net502));
 sky130_fd_sc_hd__mux4_1 c752 (.A0(net424),
    .A1(net354),
    .A2(net973),
    .A3(net887),
    .S0(net893),
    .S1(net838),
    .X(net503));
 sky130_fd_sc_hd__mux4_1 c753 (.A0(net84),
    .A1(net110),
    .A2(net493),
    .A3(net972),
    .S0(net841),
    .S1(net743),
    .X(net504));
 sky130_fd_sc_hd__mux4_1 c754 (.A0(net667),
    .A1(net681),
    .A2(net738),
    .A3(net600),
    .S0(net743),
    .S1(net617),
    .X(net505));
 sky130_fd_sc_hd__mux4_1 c755 (.A0(net624),
    .A1(net187),
    .A2(net668),
    .A3(net923),
    .S0(net744),
    .S1(net613),
    .X(net506));
 sky130_fd_sc_hd__mux4_1 c756 (.A0(net506),
    .A1(net31),
    .A2(net392),
    .A3(net629),
    .S0(net845),
    .S1(net611),
    .X(net507));
 sky130_fd_sc_hd__mux4_1 c757 (.A0(net818),
    .A1(net460),
    .A2(net480),
    .A3(net667),
    .S0(net194),
    .S1(net753),
    .X(net508));
 sky130_fd_sc_hd__mux4_1 c758 (.A0(net22),
    .A1(net40),
    .A2(net398),
    .A3(net173),
    .S0(net600),
    .S1(net820),
    .X(net509));
 sky130_fd_sc_hd__mux4_1 c759 (.A0(net722),
    .A1(net407),
    .A2(net641),
    .A3(net923),
    .S0(net597),
    .S1(net841),
    .X(net510));
 sky130_fd_sc_hd__mux4_1 c760 (.A0(net265),
    .A1(net187),
    .A2(net645),
    .A3(net600),
    .S0(net606),
    .S1(net611),
    .X(net511));
 sky130_fd_sc_hd__mux4_1 c761 (.A0(net343),
    .A1(clknet_1_0__leaf_net370),
    .A2(net22),
    .A3(net722),
    .S0(net724),
    .S1(net616),
    .X(net512));
 sky130_fd_sc_hd__mux4_1 c762 (.A0(net505),
    .A1(net656),
    .A2(net110),
    .A3(net609),
    .S0(net611),
    .S1(net613),
    .X(net513));
 sky130_fd_sc_hd__mux4_1 c763 (.A0(clknet_1_1__leaf_net255),
    .A1(net194),
    .A2(net485),
    .A3(clknet_1_0__leaf_net512),
    .S0(net511),
    .S1(net744),
    .X(net514));
 sky130_fd_sc_hd__mux4_1 c764 (.A0(net692),
    .A1(net68),
    .A2(net108),
    .A3(net838),
    .S0(net759),
    .S1(clknet_1_1__leaf_net615),
    .X(net515));
 sky130_fd_sc_hd__mux4_1 c765 (.A0(net681),
    .A1(net624),
    .A2(net511),
    .A3(net738),
    .S0(clknet_1_1__leaf_net512),
    .S1(net600),
    .X(net516));
 sky130_fd_sc_hd__mux4_1 c766 (.A0(net702),
    .A1(clknet_1_1__leaf_net400),
    .A2(net492),
    .A3(net488),
    .S0(net597),
    .S1(net619),
    .X(net517));
 sky130_fd_sc_hd__mux4_1 c767 (.A0(net683),
    .A1(net698),
    .A2(net463),
    .A3(net515),
    .S0(net725),
    .S1(net609),
    .X(net518));
 sky130_fd_sc_hd__mux4_1 c768 (.A0(net513),
    .A1(net117),
    .A2(net667),
    .A3(net517),
    .S0(net957),
    .S1(net617),
    .X(net519));
 sky130_fd_sc_hd__mux4_1 c769 (.A0(net429),
    .A1(net519),
    .A2(net518),
    .A3(net625),
    .S0(clknet_1_1__leaf_net615),
    .S1(net619),
    .X(net520));
 sky130_fd_sc_hd__mux4_1 merge790 (.A0(net169),
    .A1(clknet_1_0__leaf_net162),
    .A2(net694),
    .A3(net171),
    .S0(net755),
    .S1(net819),
    .X(net521));
 sky130_fd_sc_hd__a2111o_1 merge791 (.A1(net244),
    .A2(clknet_1_1__leaf_net161),
    .B1(net625),
    .C1(net121),
    .D1(net246),
    .X(net522));
 sky130_fd_sc_hd__mux4_1 merge792 (.A0(net55),
    .A1(net74),
    .A2(net810),
    .A3(net92),
    .S0(net86),
    .S1(net912),
    .X(net523));
 sky130_fd_sc_hd__mux4_1 merge793 (.A0(net320),
    .A1(net634),
    .A2(net330),
    .A3(net331),
    .S0(net843),
    .S1(net830),
    .X(net524));
 sky130_fd_sc_hd__mux4_1 merge794 (.A0(net258),
    .A1(net132),
    .A2(net761),
    .A3(net708),
    .S0(net914),
    .S1(net180),
    .X(net525));
 sky130_fd_sc_hd__mux4_1 merge795 (.A0(net330),
    .A1(net870),
    .A2(net311),
    .A3(net233),
    .S0(net232),
    .S1(net767),
    .X(net526));
 sky130_fd_sc_hd__mux4_1 merge796 (.A0(net74),
    .A1(net77),
    .A2(net79),
    .A3(net88),
    .S0(net95),
    .S1(net698),
    .X(net527));
 sky130_fd_sc_hd__mux4_1 merge797 (.A0(clknet_1_0__leaf_net162),
    .A1(net47),
    .A2(net158),
    .A3(net155),
    .S0(net757),
    .S1(net169),
    .X(net528));
 sky130_fd_sc_hd__and2_0 merge798 (.A(net164),
    .B(net528),
    .X(net529));
 sky130_fd_sc_hd__and2_0 merge799 (.A(net174),
    .B(net521),
    .X(net530));
 sky130_fd_sc_hd__and2_0 merge800 (.A(net285),
    .B(net269),
    .X(net531));
 sky130_fd_sc_hd__and2_0 merge801 (.A(net235),
    .B(net241),
    .X(net532));
 sky130_fd_sc_hd__and2_4 merge802 (.A(net467),
    .B(net474),
    .X(net533));
 sky130_fd_sc_hd__and2_0 merge803 (.A(net349),
    .B(net350),
    .X(net534));
 sky130_fd_sc_hd__and2_0 merge804 (.A(net94),
    .B(net523),
    .X(net535));
 sky130_fd_sc_hd__and2_0 merge805 (.A(net186),
    .B(net202),
    .X(net536));
 sky130_fd_sc_hd__and2_0 merge806 (.A(net391),
    .B(net396),
    .X(net537));
 sky130_fd_sc_hd__and2_0 merge807 (.A(net287),
    .B(net294),
    .X(net538));
 sky130_fd_sc_hd__and2_0 merge808 (.A(net102),
    .B(net104),
    .X(net539));
 sky130_fd_sc_hd__and2_0 merge809 (.A(net481),
    .B(net487),
    .X(net540));
 sky130_fd_sc_hd__and2_0 merge810 (.A(net520),
    .B(net499),
    .X(net541));
 sky130_fd_sc_hd__and2_0 merge811 (.A(net376),
    .B(net379),
    .X(net542));
 sky130_fd_sc_hd__dfrbp_2 merge812 (.CLK(clknet_2_2__leaf_clk),
    .D(net425),
    .RESET_B(net430),
    .Q(net544),
    .Q_N(net543));
 sky130_fd_sc_hd__and2_0 merge813 (.A(net345),
    .B(net332),
    .X(net545));
 sky130_fd_sc_hd__and2_0 merge814 (.A(net253),
    .B(net256),
    .X(net546));
 sky130_fd_sc_hd__and2_0 merge815 (.A(net75),
    .B(net527),
    .X(net547));
 sky130_fd_sc_hd__dfrbp_1 merge816 (.CLK(clknet_2_2__leaf_clk),
    .D(net440),
    .RESET_B(net447),
    .Q(net549),
    .Q_N(net548));
 sky130_fd_sc_hd__and2_0 merge817 (.A(net264),
    .B(net522),
    .X(net550));
 sky130_fd_sc_hd__and2_0 merge818 (.A(net157),
    .B(net163),
    .X(net551));
 sky130_fd_sc_hd__and2_0 merge819 (.A(net401),
    .B(net409),
    .X(net552));
 sky130_fd_sc_hd__and2_0 merge820 (.A(net541),
    .B(net516),
    .X(net553));
 sky130_fd_sc_hd__and2_0 merge821 (.A(net101),
    .B(net103),
    .X(net554));
 sky130_fd_sc_hd__and2_0 merge822 (.A(net380),
    .B(net306),
    .X(net555));
 sky130_fd_sc_hd__and2_0 merge823 (.A(net361),
    .B(net389),
    .X(net556));
 sky130_fd_sc_hd__and2_0 merge824 (.A(net304),
    .B(net404),
    .X(net557));
 sky130_fd_sc_hd__and2_0 merge825 (.A(net364),
    .B(net525),
    .X(net558));
 sky130_fd_sc_hd__and2_0 merge826 (.A(net76),
    .B(net78),
    .X(net559));
 sky130_fd_sc_hd__and2_0 merge827 (.A(net539),
    .B(net96),
    .X(net560));
 sky130_fd_sc_hd__and2_0 merge828 (.A(net288),
    .B(net297),
    .X(net561));
 sky130_fd_sc_hd__dfrtn_1 merge829 (.CLK_N(clknet_2_2__leaf_clk),
    .D(net347),
    .RESET_B(net524),
    .Q(net562));
 sky130_fd_sc_hd__and2_0 merge830 (.A(net494),
    .B(net514),
    .X(net563));
 sky130_fd_sc_hd__and2_0 merge831 (.A(net495),
    .B(net510),
    .X(net564));
 sky130_fd_sc_hd__and2_4 merge832 (.A(net501),
    .B(net502),
    .X(net565));
 sky130_fd_sc_hd__and2_0 merge833 (.A(net564),
    .B(net286),
    .X(net566));
 sky130_fd_sc_hd__and2_0 merge834 (.A(net83),
    .B(net529),
    .X(net567));
 sky130_fd_sc_hd__and2_1 merge835 (.A(net82),
    .B(net547),
    .X(net568));
 sky130_fd_sc_hd__dfrtp_1 merge836 (.CLK(clknet_2_0__leaf_clk),
    .D(net526),
    .RESET_B(net352),
    .Q(net569));
 sky130_fd_sc_hd__and2_0 merge837 (.A(net504),
    .B(net509),
    .X(net570));
 sky130_fd_sc_hd__dfrtp_1 merge838 (.CLK(clknet_2_2__leaf_clk),
    .D(net448),
    .RESET_B(net431),
    .Q(net571));
 sky130_fd_sc_hd__dfrtp_2 merge839 (.CLK(clknet_2_0__leaf_clk),
    .D(net559),
    .RESET_B(net567),
    .Q(net572));
 sky130_fd_sc_hd__dfsbp_1 merge840 (.CLK(clknet_2_2__leaf_clk),
    .D(net344),
    .SET_B(net545),
    .Q(net574),
    .Q_N(net573));
 sky130_fd_sc_hd__and2_0 merge841 (.A(net280),
    .B(net283),
    .X(net575));
 sky130_fd_sc_hd__and2_0 merge842 (.A(net531),
    .B(net546),
    .X(net576));
 sky130_fd_sc_hd__and2_0 merge843 (.A(net535),
    .B(net554),
    .X(net577));
 sky130_fd_sc_hd__and2_1 merge844 (.A(net461),
    .B(net477),
    .X(net578));
 sky130_fd_sc_hd__and2_0 merge845 (.A(net508),
    .B(net302),
    .X(net579));
 sky130_fd_sc_hd__and2_0 merge846 (.A(net303),
    .B(net538),
    .X(net580));
 sky130_fd_sc_hd__and2_0 merge847 (.A(net472),
    .B(net563),
    .X(net581));
 sky130_fd_sc_hd__and2_0 merge848 (.A(net184),
    .B(net530),
    .X(net582));
 sky130_fd_sc_hd__and2_0 merge849 (.A(net536),
    .B(net160),
    .X(net583));
 sky130_fd_sc_hd__and2_0 merge850 (.A(net557),
    .B(net291),
    .X(net584));
 sky130_fd_sc_hd__and2_0 merge851 (.A(net377),
    .B(net552),
    .X(net585));
 sky130_fd_sc_hd__and2_0 merge852 (.A(net468),
    .B(net405),
    .X(net586));
 sky130_fd_sc_hd__and2_0 merge853 (.A(net540),
    .B(net496),
    .X(net587));
 sky130_fd_sc_hd__and2_0 merge854 (.A(net555),
    .B(net542),
    .X(net588));
 sky130_fd_sc_hd__and2_0 merge855 (.A(net386),
    .B(net537),
    .X(net589));
 sky130_fd_sc_hd__and2_0 merge856 (.A(net402),
    .B(net570),
    .X(net590));
 sky130_fd_sc_hd__and2_0 merge857 (.A(net355),
    .B(net533),
    .X(net591));
 sky130_fd_sc_hd__dfsbp_1 merge858 (.CLK(clknet_2_1__leaf_clk),
    .D(net397),
    .SET_B(net284),
    .Q(net593),
    .Q_N(net592));
 sky130_fd_sc_hd__and2_0 merge859 (.A(net534),
    .B(net565),
    .X(net594));
 sky130_fd_sc_hd__and2_0 merge860 (.A(net476),
    .B(net556),
    .X(net595));
 sky130_fd_sc_hd__and2_0 merge861 (.A(net479),
    .B(net553),
    .X(net596));
 sky130_fd_sc_hd__dfstp_2 merge862 (.CLK(clknet_2_1__leaf_clk),
    .D(net362),
    .SET_B(net507),
    .Q(net597));
 sky130_fd_sc_hd__and2_0 merge863 (.A(net550),
    .B(net575),
    .X(net598));
 sky130_fd_sc_hd__and2_0 merge864 (.A(net560),
    .B(net551),
    .X(net599));
 sky130_fd_sc_hd__dfstp_2 merge865 (.CLK(clknet_2_3__leaf_clk),
    .D(net579),
    .SET_B(net503),
    .Q(net600));
 sky130_fd_sc_hd__dfstp_1 merge866 (.CLK(clknet_2_1__leaf_clk),
    .D(net582),
    .SET_B(net568),
    .Q(net601));
 sky130_fd_sc_hd__dlrbn_2 merge867 (.D(net598),
    .GATE_N(clknet_2_0__leaf_clk),
    .RESET_B(net532),
    .Q(net753),
    .Q_N(net602));
 sky130_fd_sc_hd__dlrbn_2 merge868 (.D(net576),
    .GATE_N(clknet_2_0__leaf_clk),
    .RESET_B(net181),
    .Q(net603),
    .Q_N(net734));
 sky130_fd_sc_hd__dlrbp_1 merge869 (.D(net369),
    .GATE(clknet_2_0__leaf_clk),
    .RESET_B(net558),
    .Q(net605),
    .Q_N(net604));
 sky130_fd_sc_hd__dlrbp_1 merge870 (.D(net445),
    .GATE(clknet_2_3__leaf_clk),
    .RESET_B(net490),
    .Q(net607),
    .Q_N(net606));
 sky130_fd_sc_hd__dlrtn_4 merge871 (.D(net449),
    .GATE_N(clknet_2_3__leaf_clk),
    .RESET_B(net589),
    .Q(net608));
 sky130_fd_sc_hd__dlrtn_2 merge872 (.D(net432),
    .GATE_N(clknet_2_2__leaf_clk),
    .RESET_B(net596),
    .Q(net609));
 sky130_fd_sc_hd__dlrtn_4 merge873 (.D(net585),
    .GATE_N(clknet_2_1__leaf_clk),
    .RESET_B(net588),
    .Q(net759));
 sky130_fd_sc_hd__and2_0 merge874 (.A(net561),
    .B(net365),
    .X(net610));
 sky130_fd_sc_hd__dlrtp_4 merge875 (.GATE(clknet_2_0__leaf_clk),
    .RESET_B(net165),
    .Q(net748));
 sky130_fd_sc_hd__dlrtp_4 merge876 (.D(net591),
    .GATE(clknet_2_2__leaf_clk),
    .RESET_B(net594),
    .Q(net743));
 sky130_fd_sc_hd__dlrtp_4 merge877 (.D(net578),
    .GATE(clknet_2_3__leaf_clk),
    .RESET_B(net590),
    .Q(net611));
 sky130_fd_sc_hd__edfxbp_1 merge878 (.CLK(clknet_2_1__leaf_clk),
    .D(net580),
    .DE(net584),
    .Q(net613),
    .Q_N(net612));
 sky130_fd_sc_hd__edfxtp_1 merge879 (.CLK(clknet_2_1__leaf_clk),
    .D(net577),
    .DE(net610),
    .Q(net801));
 sky130_fd_sc_hd__sdlclkp_1 merge880 (.CLK(clknet_2_3__leaf_clk),
    .GATE(net464),
    .SCE(net595),
    .GCLK(net614));
 sky130_fd_sc_hd__sdlclkp_2 merge881 (.CLK(clknet_2_0__leaf_clk),
    .GATE(net583),
    .SCE(net599),
    .GCLK(net799));
 sky130_fd_sc_hd__sdlclkp_4 merge882 (.CLK(clknet_2_3__leaf_clk),
    .GATE(net586),
    .SCE(net581),
    .GCLK(net615));
 sky130_fd_sc_hd__dfrbp_2 merge883 (.CLK(clknet_2_0__leaf_clk),
    .D(net587),
    .RESET_B(net566),
    .Q(net617),
    .Q_N(net616));
 sky130_fd_sc_hd__dfxbp_1 s884 (.CLK(clknet_2_3__leaf_clk),
    .D(net363),
    .Q(net619),
    .Q_N(net618));
 sky130_fd_sc_hd__dfxbp_1 s885 (.CLK(clknet_2_1__leaf_clk),
    .D(net399),
    .Q(net621),
    .Q_N(net620));
 sky130_fd_sc_hd__dfxtp_2 s886 (.CLK(clknet_2_2__leaf_clk),
    .D(net454),
    .Q(net622));
 sky130_fd_sc_hd__dfxtp_2 s887 (.CLK(clknet_2_3__leaf_clk),
    .D(net483),
    .Q(net623));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Right_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Right_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Right_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Right_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Right_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Right_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Right_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Right_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Right_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Right_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Right_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Right_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Right_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Right_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Right_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Right_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Right_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Right_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Right_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Right_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Right_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_161 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_162 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_163 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_164 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_165 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_166 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_167 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_168 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_169 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_170 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_171 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_172 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_173 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_174 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_175 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_176 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_177 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_178 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_179 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_180 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_181 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_182 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Left_183 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Left_184 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Left_185 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Left_186 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Left_187 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Left_188 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Left_189 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Left_190 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Left_191 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Left_192 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Left_193 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Left_194 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Left_195 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Left_196 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Left_197 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Left_198 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Left_199 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Left_200 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Left_201 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Left_202 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Left_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1347 ();
 sky130_fd_sc_hd__buf_6 input1 (.A(in0),
    .X(net182));
 sky130_fd_sc_hd__clkbuf_2 input2 (.A(in1),
    .X(net624));
 sky130_fd_sc_hd__buf_4 input3 (.A(in10),
    .X(net625));
 sky130_fd_sc_hd__buf_4 input4 (.A(in11),
    .X(net626));
 sky130_fd_sc_hd__clkbuf_2 input5 (.A(in12),
    .X(net627));
 sky130_fd_sc_hd__clkbuf_4 input6 (.A(in13),
    .X(net628));
 sky130_fd_sc_hd__buf_4 input7 (.A(in14),
    .X(net629));
 sky130_fd_sc_hd__clkbuf_2 input8 (.A(in15),
    .X(net630));
 sky130_fd_sc_hd__clkbuf_4 input9 (.A(in16),
    .X(net631));
 sky130_fd_sc_hd__clkbuf_4 input10 (.A(in17),
    .X(net632));
 sky130_fd_sc_hd__buf_2 input11 (.A(in18),
    .X(net633));
 sky130_fd_sc_hd__buf_2 input12 (.A(in19),
    .X(net634));
 sky130_fd_sc_hd__buf_2 input13 (.A(in2),
    .X(net635));
 sky130_fd_sc_hd__clkbuf_4 input14 (.A(in20),
    .X(net636));
 sky130_fd_sc_hd__clkbuf_4 input15 (.A(in21),
    .X(net637));
 sky130_fd_sc_hd__buf_2 input16 (.A(in22),
    .X(net638));
 sky130_fd_sc_hd__clkbuf_4 input17 (.A(in23),
    .X(net639));
 sky130_fd_sc_hd__clkbuf_2 input18 (.A(in24),
    .X(net640));
 sky130_fd_sc_hd__clkbuf_4 input19 (.A(in25),
    .X(net641));
 sky130_fd_sc_hd__clkbuf_4 input20 (.A(in26),
    .X(net642));
 sky130_fd_sc_hd__buf_2 input21 (.A(in27),
    .X(net643));
 sky130_fd_sc_hd__buf_1 input22 (.A(in28),
    .X(net644));
 sky130_fd_sc_hd__clkbuf_2 input23 (.A(in29),
    .X(net645));
 sky130_fd_sc_hd__clkbuf_4 input24 (.A(in3),
    .X(net646));
 sky130_fd_sc_hd__buf_2 input25 (.A(in30),
    .X(net647));
 sky130_fd_sc_hd__clkbuf_2 input26 (.A(in31),
    .X(net648));
 sky130_fd_sc_hd__clkbuf_2 input27 (.A(in32),
    .X(net649));
 sky130_fd_sc_hd__clkbuf_4 input28 (.A(in33),
    .X(net650));
 sky130_fd_sc_hd__clkbuf_4 input29 (.A(in34),
    .X(net651));
 sky130_fd_sc_hd__buf_1 input30 (.A(in35),
    .X(net652));
 sky130_fd_sc_hd__clkbuf_4 input31 (.A(in36),
    .X(net653));
 sky130_fd_sc_hd__clkbuf_4 input32 (.A(in37),
    .X(net654));
 sky130_fd_sc_hd__clkbuf_2 input33 (.A(in38),
    .X(net655));
 sky130_fd_sc_hd__clkbuf_4 input34 (.A(in39),
    .X(net656));
 sky130_fd_sc_hd__buf_12 input35 (.A(in4),
    .X(net657));
 sky130_fd_sc_hd__buf_1 input36 (.A(in40),
    .X(net658));
 sky130_fd_sc_hd__clkbuf_2 input37 (.A(in41),
    .X(net659));
 sky130_fd_sc_hd__clkbuf_4 input38 (.A(in42),
    .X(net660));
 sky130_fd_sc_hd__clkbuf_2 input39 (.A(in43),
    .X(net661));
 sky130_fd_sc_hd__buf_2 input40 (.A(in44),
    .X(net662));
 sky130_fd_sc_hd__buf_1 input41 (.A(in45),
    .X(net663));
 sky130_fd_sc_hd__clkbuf_2 input42 (.A(in46),
    .X(net664));
 sky130_fd_sc_hd__buf_1 input43 (.A(in47),
    .X(net665));
 sky130_fd_sc_hd__buf_1 input44 (.A(in48),
    .X(net666));
 sky130_fd_sc_hd__clkbuf_4 input45 (.A(in49),
    .X(net667));
 sky130_fd_sc_hd__clkbuf_8 input46 (.A(in5),
    .X(net668));
 sky130_fd_sc_hd__dlymetal6s2s_1 input47 (.A(in50),
    .X(net669));
 sky130_fd_sc_hd__buf_1 input48 (.A(in51),
    .X(net670));
 sky130_fd_sc_hd__buf_2 input49 (.A(in52),
    .X(net671));
 sky130_fd_sc_hd__clkbuf_4 input50 (.A(in53),
    .X(net672));
 sky130_fd_sc_hd__clkbuf_2 input51 (.A(in54),
    .X(net673));
 sky130_fd_sc_hd__clkbuf_2 input52 (.A(in55),
    .X(net674));
 sky130_fd_sc_hd__buf_1 input53 (.A(in56),
    .X(net675));
 sky130_fd_sc_hd__buf_1 input54 (.A(in57),
    .X(net676));
 sky130_fd_sc_hd__clkbuf_2 input55 (.A(in58),
    .X(net677));
 sky130_fd_sc_hd__dlymetal6s2s_1 input56 (.A(in59),
    .X(net678));
 sky130_fd_sc_hd__buf_12 input57 (.A(in6),
    .X(net679));
 sky130_fd_sc_hd__buf_1 input58 (.A(in60),
    .X(net680));
 sky130_fd_sc_hd__clkbuf_4 input59 (.A(in61),
    .X(net681));
 sky130_fd_sc_hd__buf_1 input60 (.A(in62),
    .X(net682));
 sky130_fd_sc_hd__buf_4 input61 (.A(in63),
    .X(net683));
 sky130_fd_sc_hd__buf_1 input62 (.A(in64),
    .X(net684));
 sky130_fd_sc_hd__clkbuf_4 input63 (.A(in65),
    .X(net685));
 sky130_fd_sc_hd__clkbuf_1 input64 (.A(in66),
    .X(net686));
 sky130_fd_sc_hd__buf_1 input65 (.A(in67),
    .X(net687));
 sky130_fd_sc_hd__buf_1 input66 (.A(in68),
    .X(net688));
 sky130_fd_sc_hd__clkbuf_1 input67 (.A(in69),
    .X(net689));
 sky130_fd_sc_hd__clkbuf_4 input68 (.A(in7),
    .X(net690));
 sky130_fd_sc_hd__clkbuf_2 input69 (.A(in70),
    .X(net691));
 sky130_fd_sc_hd__buf_2 input70 (.A(in71),
    .X(net692));
 sky130_fd_sc_hd__clkbuf_2 input71 (.A(in72),
    .X(net693));
 sky130_fd_sc_hd__buf_1 input72 (.A(in73),
    .X(net694));
 sky130_fd_sc_hd__clkbuf_1 input73 (.A(in74),
    .X(net695));
 sky130_fd_sc_hd__dlymetal6s2s_1 input74 (.A(in75),
    .X(net696));
 sky130_fd_sc_hd__clkbuf_2 input75 (.A(in76),
    .X(net697));
 sky130_fd_sc_hd__buf_2 input76 (.A(in77),
    .X(net698));
 sky130_fd_sc_hd__clkbuf_2 input77 (.A(in78),
    .X(net699));
 sky130_fd_sc_hd__buf_1 input78 (.A(in79),
    .X(net700));
 sky130_fd_sc_hd__dlymetal6s2s_1 input79 (.A(in8),
    .X(net701));
 sky130_fd_sc_hd__clkbuf_4 input80 (.A(in80),
    .X(net702));
 sky130_fd_sc_hd__buf_1 input81 (.A(in81),
    .X(net703));
 sky130_fd_sc_hd__clkbuf_2 input82 (.A(in82),
    .X(net704));
 sky130_fd_sc_hd__buf_1 input83 (.A(in83),
    .X(net705));
 sky130_fd_sc_hd__dlymetal6s2s_1 input84 (.A(in84),
    .X(net706));
 sky130_fd_sc_hd__dlymetal6s2s_1 input85 (.A(in85),
    .X(net707));
 sky130_fd_sc_hd__clkbuf_2 input86 (.A(in86),
    .X(net708));
 sky130_fd_sc_hd__buf_2 input87 (.A(in87),
    .X(net709));
 sky130_fd_sc_hd__buf_1 input88 (.A(in88),
    .X(net710));
 sky130_fd_sc_hd__buf_1 input89 (.A(in89),
    .X(net711));
 sky130_fd_sc_hd__buf_4 input90 (.A(in9),
    .X(net712));
 sky130_fd_sc_hd__buf_2 input91 (.A(in90),
    .X(net713));
 sky130_fd_sc_hd__buf_1 input92 (.A(in91),
    .X(net714));
 sky130_fd_sc_hd__buf_1 input93 (.A(in92),
    .X(net715));
 sky130_fd_sc_hd__buf_1 input94 (.A(in93),
    .X(net716));
 sky130_fd_sc_hd__clkbuf_2 input95 (.A(in94),
    .X(net717));
 sky130_fd_sc_hd__buf_1 input96 (.A(in95),
    .X(net718));
 sky130_fd_sc_hd__dlymetal6s2s_1 input97 (.A(in96),
    .X(net719));
 sky130_fd_sc_hd__clkbuf_1 input98 (.A(in97),
    .X(net720));
 sky130_fd_sc_hd__dlymetal6s2s_1 input99 (.A(in98),
    .X(net721));
 sky130_fd_sc_hd__buf_2 input100 (.A(in99),
    .X(net722));
 sky130_fd_sc_hd__clkbuf_4 output101 (.A(net983),
    .X(out0));
 sky130_fd_sc_hd__clkbuf_4 output102 (.A(net724),
    .X(out1));
 sky130_fd_sc_hd__clkbuf_4 output103 (.A(net725),
    .X(out10));
 sky130_fd_sc_hd__clkbuf_4 output104 (.A(net726),
    .X(out12));
 sky130_fd_sc_hd__clkbuf_4 output105 (.A(net892),
    .X(out13));
 sky130_fd_sc_hd__buf_2 output106 (.A(net922),
    .X(out14));
 sky130_fd_sc_hd__clkbuf_1 output107 (.A(net729),
    .X(out15));
 sky130_fd_sc_hd__clkbuf_4 output108 (.A(net973),
    .X(out16));
 sky130_fd_sc_hd__buf_2 output109 (.A(net731),
    .X(out18));
 sky130_fd_sc_hd__buf_2 output110 (.A(net813),
    .X(out19));
 sky130_fd_sc_hd__buf_2 output111 (.A(net808),
    .X(out2));
 sky130_fd_sc_hd__buf_2 output112 (.A(net734),
    .X(out20));
 sky130_fd_sc_hd__buf_2 output113 (.A(net735),
    .X(out21));
 sky130_fd_sc_hd__buf_2 output114 (.A(net736),
    .X(out22));
 sky130_fd_sc_hd__clkbuf_4 output115 (.A(net737),
    .X(out23));
 sky130_fd_sc_hd__clkbuf_4 output116 (.A(net738),
    .X(out24));
 sky130_fd_sc_hd__buf_2 output117 (.A(net739),
    .X(out25));
 sky130_fd_sc_hd__clkbuf_4 output118 (.A(net869),
    .X(out27));
 sky130_fd_sc_hd__clkbuf_1 output119 (.A(net741),
    .X(out28));
 sky130_fd_sc_hd__clkbuf_1 output120 (.A(clknet_1_0__leaf_net742),
    .X(out29));
 sky130_fd_sc_hd__clkbuf_4 output121 (.A(net743),
    .X(out3));
 sky130_fd_sc_hd__clkbuf_4 output122 (.A(net744),
    .X(out30));
 sky130_fd_sc_hd__buf_2 output123 (.A(net745),
    .X(out31));
 sky130_fd_sc_hd__buf_2 output124 (.A(net746),
    .X(out35));
 sky130_fd_sc_hd__buf_2 output125 (.A(net747),
    .X(out36));
 sky130_fd_sc_hd__clkbuf_4 output126 (.A(net820),
    .X(out37));
 sky130_fd_sc_hd__buf_2 output127 (.A(net749),
    .X(out38));
 sky130_fd_sc_hd__buf_2 output128 (.A(net750),
    .X(out39));
 sky130_fd_sc_hd__clkbuf_4 output129 (.A(net751),
    .X(out40));
 sky130_fd_sc_hd__buf_2 output130 (.A(net904),
    .X(out41));
 sky130_fd_sc_hd__clkbuf_4 output131 (.A(net753),
    .X(out42));
 sky130_fd_sc_hd__buf_2 output132 (.A(net754),
    .X(out44));
 sky130_fd_sc_hd__buf_2 output133 (.A(net755),
    .X(out45));
 sky130_fd_sc_hd__buf_2 output134 (.A(net756),
    .X(out46));
 sky130_fd_sc_hd__buf_2 output135 (.A(net757),
    .X(out48));
 sky130_fd_sc_hd__buf_2 output136 (.A(net758),
    .X(out49));
 sky130_fd_sc_hd__clkbuf_4 output137 (.A(net759),
    .X(out5));
 sky130_fd_sc_hd__buf_2 output138 (.A(net760),
    .X(out51));
 sky130_fd_sc_hd__buf_2 output139 (.A(net761),
    .X(out52));
 sky130_fd_sc_hd__buf_2 output140 (.A(net762),
    .X(out53));
 sky130_fd_sc_hd__buf_2 output141 (.A(net814),
    .X(out54));
 sky130_fd_sc_hd__buf_2 output142 (.A(net764),
    .X(out55));
 sky130_fd_sc_hd__buf_2 output143 (.A(net765),
    .X(out57));
 sky130_fd_sc_hd__clkbuf_1 output144 (.A(clknet_1_0__leaf_net766),
    .X(out58));
 sky130_fd_sc_hd__buf_2 output145 (.A(net767),
    .X(out59));
 sky130_fd_sc_hd__buf_2 output146 (.A(net768),
    .X(out60));
 sky130_fd_sc_hd__clkbuf_1 output147 (.A(clknet_1_1__leaf_net769),
    .X(out61));
 sky130_fd_sc_hd__buf_2 output148 (.A(net770),
    .X(out62));
 sky130_fd_sc_hd__buf_2 output149 (.A(net858),
    .X(out64));
 sky130_fd_sc_hd__buf_2 output150 (.A(net772),
    .X(out65));
 sky130_fd_sc_hd__buf_2 output151 (.A(net773),
    .X(out66));
 sky130_fd_sc_hd__buf_2 output152 (.A(net774),
    .X(out67));
 sky130_fd_sc_hd__buf_2 output153 (.A(net775),
    .X(out69));
 sky130_fd_sc_hd__buf_2 output154 (.A(net776),
    .X(out70));
 sky130_fd_sc_hd__buf_2 output155 (.A(net777),
    .X(out71));
 sky130_fd_sc_hd__buf_2 output156 (.A(net778),
    .X(out72));
 sky130_fd_sc_hd__buf_2 output157 (.A(net779),
    .X(out73));
 sky130_fd_sc_hd__buf_2 output158 (.A(net780),
    .X(out75));
 sky130_fd_sc_hd__buf_2 output159 (.A(net781),
    .X(out76));
 sky130_fd_sc_hd__buf_2 output160 (.A(net782),
    .X(out77));
 sky130_fd_sc_hd__buf_2 output161 (.A(net783),
    .X(out78));
 sky130_fd_sc_hd__buf_2 output162 (.A(net784),
    .X(out79));
 sky130_fd_sc_hd__clkbuf_4 output163 (.A(net785),
    .X(out8));
 sky130_fd_sc_hd__clkbuf_1 output164 (.A(clknet_1_1__leaf_net786),
    .X(out83));
 sky130_fd_sc_hd__buf_2 output165 (.A(net787),
    .X(out84));
 sky130_fd_sc_hd__buf_2 output166 (.A(net788),
    .X(out85));
 sky130_fd_sc_hd__buf_2 output167 (.A(net789),
    .X(out86));
 sky130_fd_sc_hd__buf_2 output168 (.A(net790),
    .X(out87));
 sky130_fd_sc_hd__buf_2 output169 (.A(net791),
    .X(out88));
 sky130_fd_sc_hd__buf_2 output170 (.A(net792),
    .X(out89));
 sky130_fd_sc_hd__clkbuf_1 output171 (.A(clknet_1_1__leaf_net793),
    .X(out9));
 sky130_fd_sc_hd__buf_2 output172 (.A(net794),
    .X(out90));
 sky130_fd_sc_hd__buf_2 output173 (.A(net795),
    .X(out91));
 sky130_fd_sc_hd__buf_2 output174 (.A(net796),
    .X(out92));
 sky130_fd_sc_hd__buf_2 output175 (.A(net797),
    .X(out93));
 sky130_fd_sc_hd__buf_2 output176 (.A(net798),
    .X(out94));
 sky130_fd_sc_hd__clkbuf_1 output177 (.A(clknet_1_1__leaf_net799),
    .X(out95));
 sky130_fd_sc_hd__clkbuf_1 output178 (.A(clknet_1_1__leaf_net800),
    .X(out96));
 sky130_fd_sc_hd__clkbuf_4 output179 (.A(net837),
    .X(out97));
 sky130_fd_sc_hd__buf_2 output180 (.A(net802),
    .X(out98));
 sky130_fd_sc_hd__buf_2 output181 (.A(net861),
    .X(out99));
 sky130_fd_sc_hd__buf_6 fanout182 (.A(net735),
    .X(net804));
 sky130_fd_sc_hd__clkbuf_4 fanout183 (.A(net919),
    .X(net805));
 sky130_fd_sc_hd__buf_8 fanout184 (.A(net727),
    .X(net806));
 sky130_fd_sc_hd__buf_4 fanout185 (.A(net216),
    .X(net807));
 sky130_fd_sc_hd__clkbuf_4 fanout186 (.A(net733),
    .X(net808));
 sky130_fd_sc_hd__clkbuf_4 fanout187 (.A(net203),
    .X(net809));
 sky130_fd_sc_hd__clkbuf_4 fanout188 (.A(net69),
    .X(net810));
 sky130_fd_sc_hd__clkbuf_4 fanout189 (.A(net812),
    .X(net811));
 sky130_fd_sc_hd__clkbuf_2 fanout190 (.A(net89),
    .X(net812));
 sky130_fd_sc_hd__buf_8 fanout191 (.A(net732),
    .X(net813));
 sky130_fd_sc_hd__buf_4 fanout192 (.A(net763),
    .X(net814));
 sky130_fd_sc_hd__buf_4 fanout193 (.A(net117),
    .X(net815));
 sky130_fd_sc_hd__buf_4 fanout194 (.A(net725),
    .X(net816));
 sky130_fd_sc_hd__buf_12 fanout195 (.A(net740),
    .X(net817));
 sky130_fd_sc_hd__buf_4 fanout196 (.A(net108),
    .X(net818));
 sky130_fd_sc_hd__clkbuf_4 fanout197 (.A(net820),
    .X(net819));
 sky130_fd_sc_hd__clkbuf_4 fanout198 (.A(net748),
    .X(net820));
 sky130_fd_sc_hd__buf_4 fanout199 (.A(net107),
    .X(net821));
 sky130_fd_sc_hd__buf_6 fanout200 (.A(net823),
    .X(net822));
 sky130_fd_sc_hd__buf_6 fanout201 (.A(net824),
    .X(net823));
 sky130_fd_sc_hd__buf_6 fanout202 (.A(net825),
    .X(net824));
 sky130_fd_sc_hd__buf_8 fanout203 (.A(net730),
    .X(net825));
 sky130_fd_sc_hd__clkbuf_4 fanout204 (.A(net828),
    .X(net826));
 sky130_fd_sc_hd__buf_2 fanout205 (.A(net828),
    .X(net827));
 sky130_fd_sc_hd__buf_2 fanout206 (.A(net830),
    .X(net828));
 sky130_fd_sc_hd__buf_4 fanout207 (.A(net830),
    .X(net829));
 sky130_fd_sc_hd__buf_4 fanout208 (.A(net31),
    .X(net830));
 sky130_fd_sc_hd__buf_8 fanout209 (.A(net832),
    .X(net831));
 sky130_fd_sc_hd__buf_12 fanout210 (.A(net833),
    .X(net832));
 sky130_fd_sc_hd__buf_12 fanout211 (.A(net834),
    .X(net833));
 sky130_fd_sc_hd__buf_8 fanout212 (.A(net16),
    .X(net834));
 sky130_fd_sc_hd__buf_2 fanout213 (.A(net791),
    .X(net835));
 sky130_fd_sc_hd__buf_4 fanout214 (.A(net801),
    .X(net836));
 sky130_fd_sc_hd__clkbuf_4 wire215 (.A(net801),
    .X(net837));
 sky130_fd_sc_hd__buf_4 fanout216 (.A(net602),
    .X(net838));
 sky130_fd_sc_hd__buf_4 fanout217 (.A(net753),
    .X(net839));
 sky130_fd_sc_hd__clkbuf_4 fanout218 (.A(net841),
    .X(net840));
 sky130_fd_sc_hd__clkbuf_4 fanout219 (.A(net601),
    .X(net841));
 sky130_fd_sc_hd__clkbuf_4 fanout220 (.A(net572),
    .X(net842));
 sky130_fd_sc_hd__buf_4 fanout221 (.A(net701),
    .X(net843));
 sky130_fd_sc_hd__buf_4 fanout222 (.A(net627),
    .X(net844));
 sky130_fd_sc_hd__buf_2 fanout223 (.A(net627),
    .X(net845));
 sky130_fd_sc_hd__buf_4 fanout224 (.A(net665),
    .X(net846));
 sky130_fd_sc_hd__buf_4 fanout225 (.A(net624),
    .X(net847));
 sky130_fd_sc_hd__buf_12 fanout226 (.A(net182),
    .X(net848));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net615 (.A(net615),
    .X(clknet_0_net615));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net615 (.A(clknet_0_net615),
    .X(clknet_1_0__leaf_net615));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net615 (.A(clknet_0_net615),
    .X(clknet_1_1__leaf_net615));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net475 (.A(net475),
    .X(clknet_0_net475));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net475 (.A(clknet_0_net475),
    .X(clknet_1_0__leaf_net475));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net475 (.A(clknet_0_net475),
    .X(clknet_1_1__leaf_net475));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net799 (.A(net799),
    .X(clknet_0_net799));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net799 (.A(clknet_0_net799),
    .X(clknet_1_0__leaf_net799));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net799 (.A(clknet_0_net799),
    .X(clknet_1_1__leaf_net799));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net370 (.A(net370),
    .X(clknet_0_net370));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net370 (.A(clknet_0_net370),
    .X(clknet_1_0__leaf_net370));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net370 (.A(clknet_0_net370),
    .X(clknet_1_1__leaf_net370));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net512 (.A(net512),
    .X(clknet_0_net512));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net512 (.A(clknet_0_net512),
    .X(clknet_1_0__leaf_net512));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net512 (.A(clknet_0_net512),
    .X(clknet_1_1__leaf_net512));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net295 (.A(net295),
    .X(clknet_0_net295));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net295 (.A(clknet_0_net295),
    .X(clknet_1_0__leaf_net295));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net295 (.A(clknet_0_net295),
    .X(clknet_1_1__leaf_net295));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net400 (.A(net400),
    .X(clknet_0_net400));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net400 (.A(clknet_0_net400),
    .X(clknet_1_0__leaf_net400));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net400 (.A(clknet_0_net400),
    .X(clknet_1_1__leaf_net400));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net300 (.A(net300),
    .X(clknet_0_net300));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net300 (.A(clknet_0_net300),
    .X(clknet_1_0__leaf_net300));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net300 (.A(clknet_0_net300),
    .X(clknet_1_1__leaf_net300));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net289 (.A(net289),
    .X(clknet_0_net289));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net289 (.A(clknet_0_net289),
    .X(clknet_1_0__leaf_net289));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net289 (.A(clknet_0_net289),
    .X(clknet_1_1__leaf_net289));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net305 (.A(net305),
    .X(clknet_0_net305));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net305 (.A(clknet_0_net305),
    .X(clknet_1_0__leaf_net305));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net305 (.A(clknet_0_net305),
    .X(clknet_1_1__leaf_net305));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net301 (.A(net301),
    .X(clknet_0_net301));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net301 (.A(clknet_0_net301),
    .X(clknet_1_0__leaf_net301));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net301 (.A(clknet_0_net301),
    .X(clknet_1_1__leaf_net301));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net268 (.A(net268),
    .X(clknet_0_net268));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net268 (.A(clknet_0_net268),
    .X(clknet_1_0__leaf_net268));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net268 (.A(clknet_0_net268),
    .X(clknet_1_1__leaf_net268));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net255 (.A(net255),
    .X(clknet_0_net255));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net255 (.A(clknet_0_net255),
    .X(clknet_1_0__leaf_net255));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net255 (.A(clknet_0_net255),
    .X(clknet_1_1__leaf_net255));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net614 (.A(net614),
    .X(clknet_0_net614));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net614 (.A(clknet_0_net614),
    .X(clknet_1_0__leaf_net614));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net614 (.A(clknet_0_net614),
    .X(clknet_1_1__leaf_net614));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net473 (.A(net473),
    .X(clknet_0_net473));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net473 (.A(clknet_0_net473),
    .X(clknet_1_0__leaf_net473));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net473 (.A(clknet_0_net473),
    .X(clknet_1_1__leaf_net473));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net793 (.A(net793),
    .X(clknet_0_net793));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net793 (.A(clknet_0_net793),
    .X(clknet_1_0__leaf_net793));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net793 (.A(clknet_0_net793),
    .X(clknet_1_1__leaf_net793));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net367 (.A(net367),
    .X(clknet_0_net367));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net367 (.A(clknet_0_net367),
    .X(clknet_1_0__leaf_net367));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net367 (.A(clknet_0_net367),
    .X(clknet_1_1__leaf_net367));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net198 (.A(net198),
    .X(clknet_0_net198));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net198 (.A(clknet_0_net198),
    .X(clknet_1_0__leaf_net198));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net198 (.A(clknet_0_net198),
    .X(clknet_1_1__leaf_net198));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net199 (.A(net199),
    .X(clknet_0_net199));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net199 (.A(clknet_0_net199),
    .X(clknet_1_0__leaf_net199));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net199 (.A(clknet_0_net199),
    .X(clknet_1_1__leaf_net199));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net200 (.A(net200),
    .X(clknet_0_net200));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net200 (.A(clknet_0_net200),
    .X(clknet_1_0__leaf_net200));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net200 (.A(clknet_0_net200),
    .X(clknet_1_1__leaf_net200));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net179 (.A(net179),
    .X(clknet_0_net179));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net179 (.A(clknet_0_net179),
    .X(clknet_1_0__leaf_net179));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net179 (.A(clknet_0_net179),
    .X(clknet_1_1__leaf_net179));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net178 (.A(net178),
    .X(clknet_0_net178));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net178 (.A(clknet_0_net178),
    .X(clknet_1_0__leaf_net178));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net178 (.A(clknet_0_net178),
    .X(clknet_1_1__leaf_net178));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net375 (.A(net375),
    .X(clknet_0_net375));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net375 (.A(clknet_0_net375),
    .X(clknet_1_0__leaf_net375));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net375 (.A(clknet_0_net375),
    .X(clknet_1_1__leaf_net375));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net277 (.A(net277),
    .X(clknet_0_net277));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net277 (.A(clknet_0_net277),
    .X(clknet_1_0__leaf_net277));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net277 (.A(clknet_0_net277),
    .X(clknet_1_1__leaf_net277));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net281 (.A(net281),
    .X(clknet_0_net281));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net281 (.A(clknet_0_net281),
    .X(clknet_1_0__leaf_net281));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net281 (.A(clknet_0_net281),
    .X(clknet_1_1__leaf_net281));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net282 (.A(net282),
    .X(clknet_0_net282));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net282 (.A(clknet_0_net282),
    .X(clknet_1_0__leaf_net282));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net282 (.A(clknet_0_net282),
    .X(clknet_1_1__leaf_net282));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net276 (.A(net276),
    .X(clknet_0_net276));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net276 (.A(clknet_0_net276),
    .X(clknet_1_0__leaf_net276));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net276 (.A(clknet_0_net276),
    .X(clknet_1_1__leaf_net276));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net166 (.A(net166),
    .X(clknet_0_net166));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net166 (.A(clknet_0_net166),
    .X(clknet_1_0__leaf_net166));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net166 (.A(clknet_0_net166),
    .X(clknet_1_1__leaf_net166));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net769 (.A(net769),
    .X(clknet_0_net769));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net769 (.A(clknet_0_net769),
    .X(clknet_1_0__leaf_net769));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net769 (.A(clknet_0_net769),
    .X(clknet_1_1__leaf_net769));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net162 (.A(net162),
    .X(clknet_0_net162));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net162 (.A(clknet_0_net162),
    .X(clknet_1_0__leaf_net162));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net162 (.A(clknet_0_net162),
    .X(clknet_1_1__leaf_net162));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net161 (.A(net161),
    .X(clknet_0_net161));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net161 (.A(clknet_0_net161),
    .X(clknet_1_0__leaf_net161));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net161 (.A(clknet_0_net161),
    .X(clknet_1_1__leaf_net161));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net159 (.A(net159),
    .X(clknet_0_net159));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net159 (.A(clknet_0_net159),
    .X(clknet_1_0__leaf_net159));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net159 (.A(clknet_0_net159),
    .X(clknet_1_1__leaf_net159));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net766 (.A(net766),
    .X(clknet_0_net766));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net766 (.A(clknet_0_net766),
    .X(clknet_1_0__leaf_net766));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net766 (.A(clknet_0_net766),
    .X(clknet_1_1__leaf_net766));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net786 (.A(net786),
    .X(clknet_0_net786));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net786 (.A(clknet_0_net786),
    .X(clknet_1_0__leaf_net786));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net786 (.A(clknet_0_net786),
    .X(clknet_1_1__leaf_net786));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net742 (.A(net742),
    .X(clknet_0_net742));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net742 (.A(clknet_0_net742),
    .X(clknet_1_0__leaf_net742));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net742 (.A(clknet_0_net742),
    .X(clknet_1_1__leaf_net742));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net97 (.A(net97),
    .X(clknet_0_net97));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net97 (.A(clknet_0_net97),
    .X(clknet_1_0__leaf_net97));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net97 (.A(clknet_0_net97),
    .X(clknet_1_1__leaf_net97));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net800 (.A(net800),
    .X(clknet_0_net800));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net800 (.A(clknet_0_net800),
    .X(clknet_1_0__leaf_net800));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net800 (.A(clknet_0_net800),
    .X(clknet_1_1__leaf_net800));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer1 (.A(net897),
    .X(net849));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer2 (.A(net849),
    .X(net850));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer3 (.A(net850),
    .X(net851));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer4 (.A(net783),
    .X(net852));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer5 (.A(net783),
    .X(net853));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer6 (.A(net322),
    .X(net854));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer7 (.A(net854),
    .X(net855));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer8 (.A(net855),
    .X(net856));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer9 (.A(net322),
    .X(net857));
 sky130_fd_sc_hd__mux4_1 clone10 (.A0(net20),
    .A1(net27),
    .A2(net712),
    .A3(net633),
    .S0(net961),
    .S1(net956),
    .X(net858));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer11 (.A(net46),
    .X(net859));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer12 (.A(net859),
    .X(net860));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer13 (.A(net803),
    .X(net861));
 sky130_fd_sc_hd__dlymetal6s4s_1 rebuffer14 (.A(net317),
    .X(net862));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer15 (.A(net317),
    .X(net863));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer16 (.A(net863),
    .X(net864));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer17 (.A(net863),
    .X(net865));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer18 (.A(net863),
    .X(net866));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer19 (.A(net866),
    .X(net867));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer20 (.A(net866),
    .X(net868));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer21 (.A(net740),
    .X(net869));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer22 (.A(net732),
    .X(net870));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer23 (.A(net29),
    .X(net871));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer24 (.A(net871),
    .X(net872));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer25 (.A(net53),
    .X(net873));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer26 (.A(net873),
    .X(net874));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer27 (.A(net874),
    .X(net875));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer28 (.A(net874),
    .X(net876));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer29 (.A(net57),
    .X(net877));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer30 (.A(net877),
    .X(net878));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer31 (.A(net125),
    .X(net879));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer32 (.A(net879),
    .X(net880));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer33 (.A(net880),
    .X(net881));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer34 (.A(net767),
    .X(net882));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer35 (.A(net886),
    .X(net883));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer36 (.A(net133),
    .X(net884));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer37 (.A(net217),
    .X(net885));
 sky130_fd_sc_hd__a2111o_1 clone38 (.A1(net28),
    .A2(net208),
    .B1(net105),
    .C1(net124),
    .D1(net958),
    .X(net886));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer39 (.A(net888),
    .X(net887));
 sky130_fd_sc_hd__clkbuf_1 clone40 (.A(net740),
    .X(net888));
 sky130_fd_sc_hd__clkbuf_2 rebuffer41 (.A(net346),
    .X(net889));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer42 (.A(net891),
    .X(net890));
 sky130_fd_sc_hd__clkbuf_1 clone43 (.A(net182),
    .X(net891));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer44 (.A(net806),
    .X(net892));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer45 (.A(net892),
    .X(net893));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer46 (.A(net325),
    .X(net894));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer47 (.A(net894),
    .X(net895));
 sky130_fd_sc_hd__buf_6 rebuffer48 (.A(net312),
    .X(net896));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer49 (.A(net896),
    .X(net897));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer50 (.A(net316),
    .X(net898));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer51 (.A(net898),
    .X(net899));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer52 (.A(net138),
    .X(net900));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer53 (.A(net900),
    .X(net901));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer54 (.A(net900),
    .X(net902));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer55 (.A(net138),
    .X(net903));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer56 (.A(net752),
    .X(net904));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer57 (.A(net934),
    .X(net905));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer58 (.A(net307),
    .X(net906));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer59 (.A(net906),
    .X(net907));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer60 (.A(net920),
    .X(net908));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer61 (.A(net908),
    .X(net909));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer62 (.A(net771),
    .X(net910));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer63 (.A(net93),
    .X(net911));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer64 (.A(net911),
    .X(net912));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer65 (.A(net93),
    .X(net913));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer66 (.A(net913),
    .X(net914));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer67 (.A(net338),
    .X(net915));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer68 (.A(net319),
    .X(net916));
 sky130_fd_sc_hd__dlymetal6s4s_1 rebuffer69 (.A(net918),
    .X(net917));
 sky130_fd_sc_hd__clkbuf_1 rebuffer70 (.A(net438),
    .X(net918));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer71 (.A(net806),
    .X(net919));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer72 (.A(net329),
    .X(net920));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer73 (.A(net728),
    .X(net921));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer74 (.A(net921),
    .X(net922));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer75 (.A(net922),
    .X(net923));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer76 (.A(net728),
    .X(net924));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer77 (.A(net222),
    .X(net925));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer78 (.A(net925),
    .X(net926));
 sky130_fd_sc_hd__clkbuf_1 rebuffer79 (.A(net925),
    .X(net927));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer80 (.A(net411),
    .X(net928));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer81 (.A(net928),
    .X(net929));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer82 (.A(net411),
    .X(net930));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer83 (.A(net219),
    .X(net931));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer84 (.A(net931),
    .X(net932));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer85 (.A(net43),
    .X(net933));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer86 (.A(net935),
    .X(net934));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer87 (.A(net936),
    .X(net935));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer88 (.A(net937),
    .X(net936));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer89 (.A(net938),
    .X(net937));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer90 (.A(net939),
    .X(net938));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer91 (.A(net940),
    .X(net939));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer92 (.A(net941),
    .X(net940));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer93 (.A(net942),
    .X(net941));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer94 (.A(net752),
    .X(net942));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer95 (.A(net336),
    .X(net943));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer96 (.A(net943),
    .X(net944));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer97 (.A(net834),
    .X(net945));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer98 (.A(net834),
    .X(net946));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer99 (.A(net946),
    .X(net947));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer100 (.A(net947),
    .X(net948));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer101 (.A(net946),
    .X(net949));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer102 (.A(net39),
    .X(net950));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer103 (.A(net950),
    .X(net951));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer104 (.A(net950),
    .X(net952));
 sky130_fd_sc_hd__buf_6 rebuffer105 (.A(net657),
    .X(net953));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer106 (.A(net953),
    .X(net954));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer107 (.A(net954),
    .X(net955));
 sky130_fd_sc_hd__clkbuf_1 clone108 (.A(net832),
    .X(net956));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer109 (.A(net657),
    .X(net957));
 sky130_fd_sc_hd__dlygate4sd3_1 hold111 (.A(net608),
    .X(net959));
 sky130_fd_sc_hd__dlygate4sd3_1 hold112 (.A(net429),
    .X(net960));
 sky130_fd_sc_hd__buf_4 fanout1 (.A(net809),
    .X(net958));
 sky130_fd_sc_hd__buf_8 fanout2 (.A(net822),
    .X(net961));
 sky130_fd_sc_hd__clkbuf_1 fanout3 (.A(net712),
    .X(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_A (.DIODE(clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(in0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(in1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(in10));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(in11));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(in12));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(in13));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(in14));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(in15));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(in16));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(in17));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(in18));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(in19));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(in2));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(in20));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(in21));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(in22));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(in23));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(in24));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(in25));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(in26));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(in27));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_A (.DIODE(in28));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_A (.DIODE(in29));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_A (.DIODE(in3));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_A (.DIODE(in30));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_A (.DIODE(in31));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_A (.DIODE(in32));
 sky130_fd_sc_hd__diode_2 ANTENNA_input28_A (.DIODE(in33));
 sky130_fd_sc_hd__diode_2 ANTENNA_input29_A (.DIODE(in34));
 sky130_fd_sc_hd__diode_2 ANTENNA_input30_A (.DIODE(in35));
 sky130_fd_sc_hd__diode_2 ANTENNA_input31_A (.DIODE(in36));
 sky130_fd_sc_hd__diode_2 ANTENNA_input32_A (.DIODE(in37));
 sky130_fd_sc_hd__diode_2 ANTENNA_input33_A (.DIODE(in38));
 sky130_fd_sc_hd__diode_2 ANTENNA_input34_A (.DIODE(in39));
 sky130_fd_sc_hd__diode_2 ANTENNA_input35_A (.DIODE(in4));
 sky130_fd_sc_hd__diode_2 ANTENNA_input36_A (.DIODE(in40));
 sky130_fd_sc_hd__diode_2 ANTENNA_input37_A (.DIODE(in41));
 sky130_fd_sc_hd__diode_2 ANTENNA_input38_A (.DIODE(in42));
 sky130_fd_sc_hd__diode_2 ANTENNA_input39_A (.DIODE(in43));
 sky130_fd_sc_hd__diode_2 ANTENNA_input40_A (.DIODE(in44));
 sky130_fd_sc_hd__diode_2 ANTENNA_input41_A (.DIODE(in45));
 sky130_fd_sc_hd__diode_2 ANTENNA_input42_A (.DIODE(in46));
 sky130_fd_sc_hd__diode_2 ANTENNA_input43_A (.DIODE(in47));
 sky130_fd_sc_hd__diode_2 ANTENNA_input44_A (.DIODE(in48));
 sky130_fd_sc_hd__diode_2 ANTENNA_input45_A (.DIODE(in49));
 sky130_fd_sc_hd__diode_2 ANTENNA_input46_A (.DIODE(in5));
 sky130_fd_sc_hd__diode_2 ANTENNA_input47_A (.DIODE(in50));
 sky130_fd_sc_hd__diode_2 ANTENNA_input48_A (.DIODE(in51));
 sky130_fd_sc_hd__diode_2 ANTENNA_input49_A (.DIODE(in52));
 sky130_fd_sc_hd__diode_2 ANTENNA_input50_A (.DIODE(in53));
 sky130_fd_sc_hd__diode_2 ANTENNA_input51_A (.DIODE(in54));
 sky130_fd_sc_hd__diode_2 ANTENNA_input52_A (.DIODE(in55));
 sky130_fd_sc_hd__diode_2 ANTENNA_input53_A (.DIODE(in56));
 sky130_fd_sc_hd__diode_2 ANTENNA_input54_A (.DIODE(in57));
 sky130_fd_sc_hd__diode_2 ANTENNA_input55_A (.DIODE(in58));
 sky130_fd_sc_hd__diode_2 ANTENNA_input56_A (.DIODE(in59));
 sky130_fd_sc_hd__diode_2 ANTENNA_input57_A (.DIODE(in6));
 sky130_fd_sc_hd__diode_2 ANTENNA_input58_A (.DIODE(in60));
 sky130_fd_sc_hd__diode_2 ANTENNA_input59_A (.DIODE(in61));
 sky130_fd_sc_hd__diode_2 ANTENNA_input60_A (.DIODE(in62));
 sky130_fd_sc_hd__diode_2 ANTENNA_input61_A (.DIODE(in63));
 sky130_fd_sc_hd__diode_2 ANTENNA_input62_A (.DIODE(in64));
 sky130_fd_sc_hd__diode_2 ANTENNA_input63_A (.DIODE(in65));
 sky130_fd_sc_hd__diode_2 ANTENNA_input64_A (.DIODE(in66));
 sky130_fd_sc_hd__diode_2 ANTENNA_input65_A (.DIODE(in67));
 sky130_fd_sc_hd__diode_2 ANTENNA_input66_A (.DIODE(in68));
 sky130_fd_sc_hd__diode_2 ANTENNA_input67_A (.DIODE(in69));
 sky130_fd_sc_hd__diode_2 ANTENNA_input68_A (.DIODE(in7));
 sky130_fd_sc_hd__diode_2 ANTENNA_input69_A (.DIODE(in70));
 sky130_fd_sc_hd__diode_2 ANTENNA_input70_A (.DIODE(in71));
 sky130_fd_sc_hd__diode_2 ANTENNA_input71_A (.DIODE(in72));
 sky130_fd_sc_hd__diode_2 ANTENNA_input72_A (.DIODE(in73));
 sky130_fd_sc_hd__diode_2 ANTENNA_input73_A (.DIODE(in74));
 sky130_fd_sc_hd__diode_2 ANTENNA_input74_A (.DIODE(in75));
 sky130_fd_sc_hd__diode_2 ANTENNA_input75_A (.DIODE(in76));
 sky130_fd_sc_hd__diode_2 ANTENNA_input76_A (.DIODE(in77));
 sky130_fd_sc_hd__diode_2 ANTENNA_input77_A (.DIODE(in78));
 sky130_fd_sc_hd__diode_2 ANTENNA_input78_A (.DIODE(in79));
 sky130_fd_sc_hd__diode_2 ANTENNA_input79_A (.DIODE(in8));
 sky130_fd_sc_hd__diode_2 ANTENNA_input80_A (.DIODE(in80));
 sky130_fd_sc_hd__diode_2 ANTENNA_input81_A (.DIODE(in81));
 sky130_fd_sc_hd__diode_2 ANTENNA_input82_A (.DIODE(in82));
 sky130_fd_sc_hd__diode_2 ANTENNA_input83_A (.DIODE(in83));
 sky130_fd_sc_hd__diode_2 ANTENNA_input84_A (.DIODE(in84));
 sky130_fd_sc_hd__diode_2 ANTENNA_input85_A (.DIODE(in85));
 sky130_fd_sc_hd__diode_2 ANTENNA_input86_A (.DIODE(in86));
 sky130_fd_sc_hd__diode_2 ANTENNA_input87_A (.DIODE(in87));
 sky130_fd_sc_hd__diode_2 ANTENNA_input88_A (.DIODE(in88));
 sky130_fd_sc_hd__diode_2 ANTENNA_input89_A (.DIODE(in89));
 sky130_fd_sc_hd__diode_2 ANTENNA_input90_A (.DIODE(in9));
 sky130_fd_sc_hd__diode_2 ANTENNA_input91_A (.DIODE(in90));
 sky130_fd_sc_hd__diode_2 ANTENNA_input92_A (.DIODE(in91));
 sky130_fd_sc_hd__diode_2 ANTENNA_input93_A (.DIODE(in92));
 sky130_fd_sc_hd__diode_2 ANTENNA_input94_A (.DIODE(in93));
 sky130_fd_sc_hd__diode_2 ANTENNA_input95_A (.DIODE(in94));
 sky130_fd_sc_hd__diode_2 ANTENNA_input96_A (.DIODE(in95));
 sky130_fd_sc_hd__diode_2 ANTENNA_input97_A (.DIODE(in96));
 sky130_fd_sc_hd__diode_2 ANTENNA_input98_A (.DIODE(in97));
 sky130_fd_sc_hd__diode_2 ANTENNA_input99_A (.DIODE(in98));
 sky130_fd_sc_hd__diode_2 ANTENNA_input100_A (.DIODE(in99));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone38_B1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c542_A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c405_B1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c400_B (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c275_A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c264_X (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout199_A (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c564_D_N (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c266_X (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout196_A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA_c764_A2 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA_c267_X (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA_c762_A2 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_A1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c739_S0 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_S1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_A3 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_A2 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_A1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c283_A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c269_X (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c548_A1 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_c529_B (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_c528_B (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_c407_B (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_S0 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_B (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_c270_X (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_A1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c410_A2 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c404_A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c365_B (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_A2 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c313_C_N (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_D_N (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c279_C_N (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c271_X (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_A2 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_C_N (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_S1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c279_B (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c275_B (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c273_A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c272_X (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_A0 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_c615_A2 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_c610_A3 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_c494_A3 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_c412_S1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_B (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_A3 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_A (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_c273_X (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_c366_A1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_A0 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_B (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_B (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c274_X (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c680_C1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c678_D (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c676_D1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c411_S1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c402_A2 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c399_B (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_A0 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_C (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c278_B (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c277_B (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c275_X (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout193_A (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c768_A1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c276_X (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_A0 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_A0 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_C1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_A3 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c297_A1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c278_X (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge791_C1 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c556_B1 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c533_A3 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c529_A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_B (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_B (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_X (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_A0 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_A3 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_A0 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_A1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c283_B (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_B1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_X (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c687_C1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_A2 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_A1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c667_A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c545_C_N (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c446_B (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c430_C_N (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_A1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c412_S0 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_X (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone38_C1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c405_C1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c687_A1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c677_SCD (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c674_B (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c668_D1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c542_B (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_D_N (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_A1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c283_X (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c742_A0 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_A1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_S1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_B (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_c295_B (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_S1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_A (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_X (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_A1 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA_c586_C1 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA_c565_A2 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_C (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_A (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA_c295_D_N (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_A (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_X (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge794_A1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_A (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_C (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_A2 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_X (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_c686_A1 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_c558_B (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_B (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_X (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_A0 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_A3 (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA_c700_B (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_A1 (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_C_N (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_C1 (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_A (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_S0 (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_A (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_C (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_X (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_B (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_B (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_A0 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_X (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_A3 (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_A1 (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_c701_S0 (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_C_N (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_A1 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_B (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_C1 (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_X (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_A0 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_C1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_A2 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_A3 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_A2 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_X (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_A0 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_A0 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_A1 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_c311_X (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_B1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_A0 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_A0 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_X (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_A3 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_A (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_A2 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_B (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_D1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_X (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_c494_S0 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_A0 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_S0 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_A2 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_S0 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_S0 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_C1 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA_c321_D1 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_D1 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_X (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_A1 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA_c323_A1 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_A2 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_X (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA_c371_A (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_S0 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_B (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_A2 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_S1 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_B1 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_X (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge797_S1 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge790_A0 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_A1 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_A0 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_S1 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_X (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_c531_A (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c403_B (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c271_C (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c266_C (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_B (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c140_A (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c138_B (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c136_A (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_X (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_A3 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA_c744_A2 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_A1 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_A1 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_A3 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA_c502_S0 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA_c366_A3 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_A1 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_A2 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_X (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net178_A (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_X (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA_c760_A1 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A1 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_X (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_A1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_A2 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_X (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_A1 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_A2 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_X (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_c763_A1 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA_c757_S0 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_C1 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA_c364_X (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_A2 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_A1 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_X (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone10_A0 (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c434_A (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c271_B (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c267_B (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_A2 (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_A0 (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_A1 (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_X (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_A1 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_A1 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_S0 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_A3 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_A2 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_c373_D1 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_c372_X (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone38_A2 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_A0 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_C (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA_c405_A2 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA_c401_X (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA_c407_C (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_c664_A (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_c547_A3 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_c403_X (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_c672_A (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c666_B (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c538_B (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c537_C_N (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_A0 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c143_B (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c140_X (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c670_A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA_c532_C_N (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA_c415_B (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA_c412_A0 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA_c404_X (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_S0 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA_c685_A (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA_c666_C_N (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_A1 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA_c408_A (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA_c406_X (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA_c702_A (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_c686_A2 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_C_N (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_c548_C1 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_c428_C (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_c409_X (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout185_A (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_A2 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA_c410_X (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA_c761_A2 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_A0 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_S0 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_A3 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_A3 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_A2 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_S0 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_B1 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_S0 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_A3 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_X (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_A3 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_A0 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_A2 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_C (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_A2 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_S0 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA_c416_B (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA_c415_X (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_A3 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_A0 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_c614_A2 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_B1 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_A2 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_X (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_A0 (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_c691_A0 (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c686_C1 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA_c558_C_N (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_X (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA_c723_A1 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_A3 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_A3 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_A2 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_c556_D1 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_A0 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_C (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_X (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_A0 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_S0 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA_c702_B (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA_c566_A2 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_B (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_X (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_A2 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_S0 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_A1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_A3 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_A3 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA_c427_C (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA_c424_X (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge795_S0 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_A1 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_A1 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c556_A2 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_D1 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c430_A (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c427_X (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_A3 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_C (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_A0 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_S0 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_B (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c431_X (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_B1 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA_c582_A (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_C (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_S1 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_X (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_A3 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_S0 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_A (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_A1 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_c434_X (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_A0 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_C_N (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_C1 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_D1 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_c437_X (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_c703_S0 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_A (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_A1 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_B (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_X (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_A0 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_A2 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_A1 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_A2 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_X (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_A1 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_C1 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_S0 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_A (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_X (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_A2 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_A1 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_c566_A3 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_c561_B (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_c311_D_N (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_S0 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_A2 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_A (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_X (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_c206_A (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c198_B (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_A2 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_S0 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_A0 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_X (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_A2 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_A1 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_A1 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_A1 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_X (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA_c760_A0 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_A2 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_A2 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_S0 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_D1 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_X (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_A1 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA_c745_A1 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_X (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone10_A1 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_A3 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_c411_A1 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_c401_A (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_C (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_c264_B (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_A (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_A1 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_X (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_c402_D1 (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer23_A (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_B (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c545_D_N (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_A (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_S0 (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_X (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_A1 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_X (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_A0 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_B (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_A3 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_c182_A (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_A1 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_X (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge845_B (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_X (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_A (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA_c678_RESET_B (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA_c667_B (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA_c661_B (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA_c529_X (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout208_A (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_A1 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_D1 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_X (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_A1 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_A2 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA_c535_B (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA_c532_D_N (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA_c531_X (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge795_A2 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_A2 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA_c698_C_N (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA_c695_A (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA_c660_B (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA_c611_A1 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA_c544_S0 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA_c532_X (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_S0 (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_A1 (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA_c565_A1 (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_B1 (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA_c548_D1 (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA_c545_A (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA_c543_B (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA_c535_X (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A0 (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_B (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA_c564_B (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA_c544_A2 (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA_c539_X (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_S0 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_A2 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA_c549_A (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA_c548_X (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_D (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_A1 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_A1 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_A1 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA_c586_B1 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA_c558_X (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_A0 (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_A3 (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_A3 (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_A2 (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_A3 (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_B (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_A1 (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_SCE (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA_c565_X (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA_c761_A0 (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_B (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA_c587_A2 (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_Q (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_A1 (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A3 (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_A1 (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_A2 (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_A1 (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_A1 (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_A2 (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_S1 (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_D1 (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA_c577_X (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_A1 (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_A0 (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_B1 (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_A3 (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_X (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge862_D (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA_c586_X (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge874_B (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_X (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_A0 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c739_A2 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_A1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_A1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_X (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c229_A (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_S0 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_B (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_A1 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_X (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_A3 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_S0 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_S0 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_A0 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA_c615_A1 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA_c614_A3 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA_c613_S0 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_X (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_A1 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_c744_S0 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_A1 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_A1 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_A (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_X (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge852_B (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA_c633_X (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_A1 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_S0 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_A0 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_A2 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_C (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_X (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_c742_A2 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_A0 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_A2 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_A1 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_c668_A2 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_c660_X (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_c742_A1 (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_A0 (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA_c723_A3 (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_A3 (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_B1 (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA_c703_A3 (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA_c678_SCE (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA_c665_X (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_C1 (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_D (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA_c674_C (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA_c666_X (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_A2 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_A3 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_A2 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_D1 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_B (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_c437_D_N (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_c216_A1 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_X (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_A0 (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA_c681_A0 (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA_c680_A2 (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA_c679_C1 (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA_c678_SCD (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA_c677_SCE (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA_c676_B1 (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA_c675_X (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold112_A (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA_c769_A0 (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_A1 (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_B1 (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA_c678_Q (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_D1 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer85_A (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_c582_D_N (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_c564_C_N (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_c554_B (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_c184_S0 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_A3 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_X (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_c746_A2 (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA_c743_A3 (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA_c739_A3 (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A1 (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_X (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_A (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_c370_B (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_c344_C1 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_A1 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_A1 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_X (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_c743_S1 (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_A0 (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_S0 (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_A2 (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA_c700_X (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_A1 (.DIODE(net457));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_A1 (.DIODE(net457));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_SCE (.DIODE(net457));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_Q (.DIODE(net457));
 sky130_fd_sc_hd__diode_2 ANTENNA_c767_A2 (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_S0 (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA_c745_A2 (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_X (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge797_A1 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_A0 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_B1 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_A2 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_B1 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA_c203_C (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA_c180_C (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_B (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_X (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_A1 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_A2 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_D1 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_X (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_A1 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_A1 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_A1 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_c311_C_N (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_c208_S1 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_A2 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_c182_X (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_A3 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_A1 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_c613_A2 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_A2 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_C (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_c236_S0 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_S0 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_A (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_D_N (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_X (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge812_Q (.DIODE(net544));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_S0 (.DIODE(net544));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_A3 (.DIODE(net544));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_D1 (.DIODE(net544));
 sky130_fd_sc_hd__diode_2 ANTENNA_c502_A0 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_A1 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_C (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_A1 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_X (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge877_D (.DIODE(net578));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge844_X (.DIODE(net578));
 sky130_fd_sc_hd__diode_2 ANTENNA_c739_A1 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_A2 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_A2 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_A3 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_C (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_A0 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_D_N (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA_c194_C1 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_X (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge862_Q (.DIODE(net597));
 sky130_fd_sc_hd__diode_2 ANTENNA_c766_S0 (.DIODE(net597));
 sky130_fd_sc_hd__diode_2 ANTENNA_c759_S0 (.DIODE(net597));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_S0 (.DIODE(net597));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_S0 (.DIODE(net597));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge865_Q (.DIODE(net600));
 sky130_fd_sc_hd__diode_2 ANTENNA_c765_S1 (.DIODE(net600));
 sky130_fd_sc_hd__diode_2 ANTENNA_c760_A3 (.DIODE(net600));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_S0 (.DIODE(net600));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A3 (.DIODE(net600));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_S1 (.DIODE(net600));
 sky130_fd_sc_hd__diode_2 ANTENNA_c502_S1 (.DIODE(net600));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout216_A (.DIODE(net602));
 sky130_fd_sc_hd__diode_2 ANTENNA_c611_S1 (.DIODE(net602));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_S0 (.DIODE(net602));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge867_Q_N (.DIODE(net602));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge868_Q (.DIODE(net603));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_C1 (.DIODE(net603));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_S1 (.DIODE(net603));
 sky130_fd_sc_hd__diode_2 ANTENNA_c482_S1 (.DIODE(net603));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_D1 (.DIODE(net603));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_D1 (.DIODE(net603));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_S1 (.DIODE(net603));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_S1 (.DIODE(net603));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge869_Q (.DIODE(net605));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_A3 (.DIODE(net605));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_A3 (.DIODE(net605));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_A3 (.DIODE(net605));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold111_A (.DIODE(net608));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge871_Q (.DIODE(net608));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_S1 (.DIODE(net608));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_S0 (.DIODE(net608));
 sky130_fd_sc_hd__diode_2 ANTENNA_c703_S1 (.DIODE(net608));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_S0 (.DIODE(net608));
 sky130_fd_sc_hd__diode_2 ANTENNA_c613_S1 (.DIODE(net608));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_D1 (.DIODE(net608));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge872_Q (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA_c767_S1 (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA_c762_A3 (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_S0 (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_S0 (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA_c701_S1 (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_S1 (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA_c691_S1 (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA_c364_A (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_A2 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_A2 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA_c323_A3 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA_c194_X (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge877_Q (.DIODE(net611));
 sky130_fd_sc_hd__diode_2 ANTENNA_c762_S0 (.DIODE(net611));
 sky130_fd_sc_hd__diode_2 ANTENNA_c760_S1 (.DIODE(net611));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_S1 (.DIODE(net611));
 sky130_fd_sc_hd__diode_2 ANTENNA_c745_S0 (.DIODE(net611));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_S0 (.DIODE(net611));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_D1 (.DIODE(net611));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_S1 (.DIODE(net611));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_S0 (.DIODE(net611));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge878_Q_N (.DIODE(net612));
 sky130_fd_sc_hd__diode_2 ANTENNA_c633_S1 (.DIODE(net612));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_S1 (.DIODE(net612));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_S1 (.DIODE(net612));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_S1 (.DIODE(net612));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge878_Q (.DIODE(net613));
 sky130_fd_sc_hd__diode_2 ANTENNA_c762_S1 (.DIODE(net613));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_S1 (.DIODE(net613));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_S1 (.DIODE(net613));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_S1 (.DIODE(net613));
 sky130_fd_sc_hd__diode_2 ANTENNA_c496_D1 (.DIODE(net613));
 sky130_fd_sc_hd__diode_2 ANTENNA_s886_Q (.DIODE(net622));
 sky130_fd_sc_hd__diode_2 ANTENNA_c747_S0 (.DIODE(net622));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_S1 (.DIODE(net622));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_S1 (.DIODE(net622));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_S1 (.DIODE(net622));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_S1 (.DIODE(net622));
 sky130_fd_sc_hd__diode_2 ANTENNA_s887_Q (.DIODE(net623));
 sky130_fd_sc_hd__diode_2 ANTENNA_c747_S1 (.DIODE(net623));
 sky130_fd_sc_hd__diode_2 ANTENNA_c746_S1 (.DIODE(net623));
 sky130_fd_sc_hd__diode_2 ANTENNA_c742_S1 (.DIODE(net623));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_S1 (.DIODE(net623));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_S1 (.DIODE(net623));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_S1 (.DIODE(net623));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_S1 (.DIODE(net623));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_S1 (.DIODE(net623));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_A1 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_A3 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_B1 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_A (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA_c198_X (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_S1 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_A1 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_S0 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_B (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_C (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_B1 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_c208_A3 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_A2 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_c203_A (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_X (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_c764_A1 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_A2 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_D_N (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c371_C_N (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c230_C (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c212_A1 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_X (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout188_A (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_A0 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_X (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_A3 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_A1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_C (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_B1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_c205_A (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_X (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_A2 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_B (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_B1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_c208_A0 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_X (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge796_A1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_A2 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_A3 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c218_B1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_A0 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c212_B1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_X (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c613_A0 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_A0 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_A3 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_B (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_c218_A2 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_c216_X (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_A0 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_A0 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_c221_X (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_A0 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_A2 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_c238_X (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone43_A (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout226_A (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_X (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_A1 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_A2 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_A0 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout225_A (.DIODE(net624));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_X (.DIODE(net624));
 sky130_fd_sc_hd__diode_2 ANTENNA_c765_A1 (.DIODE(net624));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A0 (.DIODE(net624));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_A2 (.DIODE(net624));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_X (.DIODE(net625));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge791_B1 (.DIODE(net625));
 sky130_fd_sc_hd__diode_2 ANTENNA_c769_A3 (.DIODE(net625));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_A0 (.DIODE(net625));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_A3 (.DIODE(net625));
 sky130_fd_sc_hd__diode_2 ANTENNA_c614_S0 (.DIODE(net625));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_C1 (.DIODE(net625));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_A (.DIODE(net625));
 sky130_fd_sc_hd__diode_2 ANTENNA_c265_A (.DIODE(net625));
 sky130_fd_sc_hd__diode_2 ANTENNA_c221_B1 (.DIODE(net625));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_X (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA_c747_A2 (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_S1 (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_B (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_A2 (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_A1 (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA_c434_C (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA_c402_C1 (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_A1 (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_A (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout223_A (.DIODE(net627));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout222_A (.DIODE(net627));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_X (.DIODE(net627));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_X (.DIODE(net628));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_A1 (.DIODE(net628));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_A0 (.DIODE(net628));
 sky130_fd_sc_hd__diode_2 ANTENNA_c410_A1 (.DIODE(net628));
 sky130_fd_sc_hd__diode_2 ANTENNA_c397_A (.DIODE(net628));
 sky130_fd_sc_hd__diode_2 ANTENNA_c241_C1 (.DIODE(net628));
 sky130_fd_sc_hd__diode_2 ANTENNA_c110_B (.DIODE(net628));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_X (.DIODE(net629));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_A3 (.DIODE(net629));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_A3 (.DIODE(net629));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_A0 (.DIODE(net629));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_A2 (.DIODE(net629));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_A3 (.DIODE(net629));
 sky130_fd_sc_hd__diode_2 ANTENNA_c614_S1 (.DIODE(net629));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_A0 (.DIODE(net629));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_S1 (.DIODE(net629));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_A (.DIODE(net629));
 sky130_fd_sc_hd__diode_2 ANTENNA_c111_B (.DIODE(net629));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_X (.DIODE(net630));
 sky130_fd_sc_hd__diode_2 ANTENNA_c180_A (.DIODE(net630));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_C (.DIODE(net630));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_A0 (.DIODE(net630));
 sky130_fd_sc_hd__diode_2 ANTENNA_c158_B (.DIODE(net630));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_B (.DIODE(net630));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_A1 (.DIODE(net630));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_X (.DIODE(net631));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_A1 (.DIODE(net631));
 sky130_fd_sc_hd__diode_2 ANTENNA_c411_A0 (.DIODE(net631));
 sky130_fd_sc_hd__diode_2 ANTENNA_c401_B (.DIODE(net631));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_A3 (.DIODE(net631));
 sky130_fd_sc_hd__diode_2 ANTENNA_c270_A (.DIODE(net631));
 sky130_fd_sc_hd__diode_2 ANTENNA_c129_A (.DIODE(net631));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_X (.DIODE(net632));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_A2 (.DIODE(net632));
 sky130_fd_sc_hd__diode_2 ANTENNA_c191_A0 (.DIODE(net632));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_C (.DIODE(net632));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_B (.DIODE(net632));
 sky130_fd_sc_hd__diode_2 ANTENNA_c130_A1 (.DIODE(net632));
 sky130_fd_sc_hd__diode_2 ANTENNA_c120_B1 (.DIODE(net632));
 sky130_fd_sc_hd__diode_2 ANTENNA_c102_A0 (.DIODE(net632));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone10_A3 (.DIODE(net633));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_X (.DIODE(net633));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_A2 (.DIODE(net633));
 sky130_fd_sc_hd__diode_2 ANTENNA_c158_A (.DIODE(net633));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_A3 (.DIODE(net633));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_B (.DIODE(net633));
 sky130_fd_sc_hd__diode_2 ANTENNA_c134_B (.DIODE(net633));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_A (.DIODE(net633));
 sky130_fd_sc_hd__diode_2 ANTENNA_c528_C (.DIODE(net634));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_X (.DIODE(net634));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge793_A1 (.DIODE(net634));
 sky130_fd_sc_hd__diode_2 ANTENNA_c533_S0 (.DIODE(net634));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_A2 (.DIODE(net634));
 sky130_fd_sc_hd__diode_2 ANTENNA_c274_B (.DIODE(net634));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_A (.DIODE(net634));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_A2 (.DIODE(net634));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_X (.DIODE(net635));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_A (.DIODE(net635));
 sky130_fd_sc_hd__diode_2 ANTENNA_c276_B (.DIODE(net635));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_A (.DIODE(net635));
 sky130_fd_sc_hd__diode_2 ANTENNA_c266_B (.DIODE(net635));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_A (.DIODE(net635));
 sky130_fd_sc_hd__diode_2 ANTENNA_c140_B (.DIODE(net635));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_X (.DIODE(net636));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_A (.DIODE(net636));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_B (.DIODE(net636));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_B (.DIODE(net636));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_A2 (.DIODE(net636));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_B (.DIODE(net636));
 sky130_fd_sc_hd__diode_2 ANTENNA_c117_C (.DIODE(net636));
 sky130_fd_sc_hd__diode_2 ANTENNA_c111_A (.DIODE(net636));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_X (.DIODE(net637));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_B (.DIODE(net637));
 sky130_fd_sc_hd__diode_2 ANTENNA_c531_B (.DIODE(net637));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_B (.DIODE(net637));
 sky130_fd_sc_hd__diode_2 ANTENNA_c408_B (.DIODE(net637));
 sky130_fd_sc_hd__diode_2 ANTENNA_c297_A0 (.DIODE(net637));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_C1 (.DIODE(net637));
 sky130_fd_sc_hd__diode_2 ANTENNA_c159_B1 (.DIODE(net637));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_A (.DIODE(net637));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_X (.DIODE(net638));
 sky130_fd_sc_hd__diode_2 ANTENNA_c369_D_N (.DIODE(net638));
 sky130_fd_sc_hd__diode_2 ANTENNA_c295_A (.DIODE(net638));
 sky130_fd_sc_hd__diode_2 ANTENNA_c260_S0 (.DIODE(net638));
 sky130_fd_sc_hd__diode_2 ANTENNA_c198_C (.DIODE(net638));
 sky130_fd_sc_hd__diode_2 ANTENNA_c122_A (.DIODE(net638));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_X (.DIODE(net639));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_A0 (.DIODE(net639));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_A3 (.DIODE(net639));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_A1 (.DIODE(net639));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_S1 (.DIODE(net639));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_A (.DIODE(net639));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_S1 (.DIODE(net639));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_X (.DIODE(net640));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_B1 (.DIODE(net640));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_B (.DIODE(net640));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_X (.DIODE(net641));
 sky130_fd_sc_hd__diode_2 ANTENNA_c759_A2 (.DIODE(net641));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_S0 (.DIODE(net641));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_A2 (.DIODE(net641));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_A (.DIODE(net641));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_C1 (.DIODE(net641));
 sky130_fd_sc_hd__diode_2 ANTENNA_c221_A1 (.DIODE(net641));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_B (.DIODE(net642));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_X (.DIODE(net642));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_A1 (.DIODE(net642));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_B1 (.DIODE(net642));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_A3 (.DIODE(net642));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_C (.DIODE(net642));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_B (.DIODE(net642));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_X (.DIODE(net643));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_A1 (.DIODE(net643));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_A1 (.DIODE(net643));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_B (.DIODE(net643));
 sky130_fd_sc_hd__diode_2 ANTENNA_c183_C (.DIODE(net643));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_A (.DIODE(net643));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_X (.DIODE(net644));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_A3 (.DIODE(net644));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_A1 (.DIODE(net644));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_D_N (.DIODE(net644));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_X (.DIODE(net645));
 sky130_fd_sc_hd__diode_2 ANTENNA_c760_A2 (.DIODE(net645));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_A3 (.DIODE(net645));
 sky130_fd_sc_hd__diode_2 ANTENNA_c610_A1 (.DIODE(net645));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_A1 (.DIODE(net645));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_C (.DIODE(net645));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_X (.DIODE(net646));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_B1 (.DIODE(net646));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_A (.DIODE(net646));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_B (.DIODE(net646));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_A (.DIODE(net646));
 sky130_fd_sc_hd__diode_2 ANTENNA_c136_B (.DIODE(net646));
 sky130_fd_sc_hd__diode_2 ANTENNA_c115_A (.DIODE(net646));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_X (.DIODE(net647));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_A1 (.DIODE(net647));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_A2 (.DIODE(net647));
 sky130_fd_sc_hd__diode_2 ANTENNA_c130_A2 (.DIODE(net647));
 sky130_fd_sc_hd__diode_2 ANTENNA_c113_A (.DIODE(net647));
 sky130_fd_sc_hd__diode_2 ANTENNA_c103_C_N (.DIODE(net647));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_X (.DIODE(net648));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_A1 (.DIODE(net648));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_A (.DIODE(net648));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_A0 (.DIODE(net648));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_S1 (.DIODE(net648));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_B (.DIODE(net648));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_X (.DIODE(net649));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_S0 (.DIODE(net649));
 sky130_fd_sc_hd__diode_2 ANTENNA_c496_A1 (.DIODE(net649));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_S1 (.DIODE(net649));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_B (.DIODE(net649));
 sky130_fd_sc_hd__diode_2 ANTENNA_c105_B (.DIODE(net649));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_B (.DIODE(net650));
 sky130_fd_sc_hd__diode_2 ANTENNA_input28_X (.DIODE(net650));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_A2 (.DIODE(net650));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_A0 (.DIODE(net650));
 sky130_fd_sc_hd__diode_2 ANTENNA_c587_S0 (.DIODE(net650));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_A1 (.DIODE(net650));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_S0 (.DIODE(net650));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_C1 (.DIODE(net650));
 sky130_fd_sc_hd__diode_2 ANTENNA_input29_X (.DIODE(net651));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_A0 (.DIODE(net651));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_A2 (.DIODE(net651));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_B (.DIODE(net651));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_D1 (.DIODE(net651));
 sky130_fd_sc_hd__diode_2 ANTENNA_c286_A (.DIODE(net651));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_S0 (.DIODE(net651));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_C_N (.DIODE(net651));
 sky130_fd_sc_hd__diode_2 ANTENNA_input31_X (.DIODE(net653));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_A1 (.DIODE(net653));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_A1 (.DIODE(net653));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_A3 (.DIODE(net653));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_S0 (.DIODE(net653));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_C (.DIODE(net653));
 sky130_fd_sc_hd__diode_2 ANTENNA_input32_X (.DIODE(net654));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_A (.DIODE(net654));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_C (.DIODE(net654));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_A (.DIODE(net654));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_A3 (.DIODE(net654));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_A2 (.DIODE(net654));
 sky130_fd_sc_hd__diode_2 ANTENNA_input33_X (.DIODE(net655));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_A0 (.DIODE(net655));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_D_N (.DIODE(net655));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_A (.DIODE(net655));
 sky130_fd_sc_hd__diode_2 ANTENNA_input34_X (.DIODE(net656));
 sky130_fd_sc_hd__diode_2 ANTENNA_c762_A1 (.DIODE(net656));
 sky130_fd_sc_hd__diode_2 ANTENNA_c745_A3 (.DIODE(net656));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_S1 (.DIODE(net656));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_C_N (.DIODE(net656));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_A2 (.DIODE(net656));
 sky130_fd_sc_hd__diode_2 ANTENNA_c428_A (.DIODE(net656));
 sky130_fd_sc_hd__diode_2 ANTENNA_c424_C_N (.DIODE(net656));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_A0 (.DIODE(net656));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_B (.DIODE(net657));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer109_A (.DIODE(net657));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer105_A (.DIODE(net657));
 sky130_fd_sc_hd__diode_2 ANTENNA_input35_X (.DIODE(net657));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_A3 (.DIODE(net657));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_SET_B (.DIODE(net657));
 sky130_fd_sc_hd__diode_2 ANTENNA_c267_A (.DIODE(net657));
 sky130_fd_sc_hd__diode_2 ANTENNA_input37_X (.DIODE(net659));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_A1 (.DIODE(net659));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_A (.DIODE(net659));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_A2 (.DIODE(net659));
 sky130_fd_sc_hd__diode_2 ANTENNA_input38_X (.DIODE(net660));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_B1 (.DIODE(net660));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_A3 (.DIODE(net660));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_RESET_B (.DIODE(net660));
 sky130_fd_sc_hd__diode_2 ANTENNA_c701_A1 (.DIODE(net660));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_D_N (.DIODE(net660));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_A1 (.DIODE(net660));
 sky130_fd_sc_hd__diode_2 ANTENNA_c565_S1 (.DIODE(net660));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_A (.DIODE(net660));
 sky130_fd_sc_hd__diode_2 ANTENNA_input39_X (.DIODE(net661));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_A (.DIODE(net661));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_B (.DIODE(net661));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_A2 (.DIODE(net661));
 sky130_fd_sc_hd__diode_2 ANTENNA_input40_X (.DIODE(net662));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_A1 (.DIODE(net662));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_S1 (.DIODE(net662));
 sky130_fd_sc_hd__diode_2 ANTENNA_c191_A3 (.DIODE(net662));
 sky130_fd_sc_hd__diode_2 ANTENNA_c104_B (.DIODE(net662));
 sky130_fd_sc_hd__diode_2 ANTENNA_input41_X (.DIODE(net663));
 sky130_fd_sc_hd__diode_2 ANTENNA_c127_A0 (.DIODE(net663));
 sky130_fd_sc_hd__diode_2 ANTENNA_c101_C (.DIODE(net663));
 sky130_fd_sc_hd__diode_2 ANTENNA_input42_X (.DIODE(net664));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_B (.DIODE(net664));
 sky130_fd_sc_hd__diode_2 ANTENNA_c259_S1 (.DIODE(net664));
 sky130_fd_sc_hd__diode_2 ANTENNA_c212_D1 (.DIODE(net664));
 sky130_fd_sc_hd__diode_2 ANTENNA_input45_X (.DIODE(net667));
 sky130_fd_sc_hd__diode_2 ANTENNA_c768_A2 (.DIODE(net667));
 sky130_fd_sc_hd__diode_2 ANTENNA_c757_A3 (.DIODE(net667));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A0 (.DIODE(net667));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_A2 (.DIODE(net667));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_S0 (.DIODE(net667));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_A3 (.DIODE(net667));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_D1 (.DIODE(net667));
 sky130_fd_sc_hd__diode_2 ANTENNA_c184_A3 (.DIODE(net667));
 sky130_fd_sc_hd__diode_2 ANTENNA_input46_X (.DIODE(net668));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A2 (.DIODE(net668));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_A0 (.DIODE(net668));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_A0 (.DIODE(net668));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_A2 (.DIODE(net668));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_A1 (.DIODE(net668));
 sky130_fd_sc_hd__diode_2 ANTENNA_c544_S1 (.DIODE(net668));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_A3 (.DIODE(net668));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_C_N (.DIODE(net668));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_B (.DIODE(net668));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_C_N (.DIODE(net668));
 sky130_fd_sc_hd__diode_2 ANTENNA_input47_X (.DIODE(net669));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_A1 (.DIODE(net669));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_A3 (.DIODE(net669));
 sky130_fd_sc_hd__diode_2 ANTENNA_c184_A0 (.DIODE(net669));
 sky130_fd_sc_hd__diode_2 ANTENNA_input48_X (.DIODE(net670));
 sky130_fd_sc_hd__diode_2 ANTENNA_c236_A0 (.DIODE(net670));
 sky130_fd_sc_hd__diode_2 ANTENNA_c206_C (.DIODE(net670));
 sky130_fd_sc_hd__diode_2 ANTENNA_c104_C (.DIODE(net670));
 sky130_fd_sc_hd__diode_2 ANTENNA_input49_X (.DIODE(net671));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_C1 (.DIODE(net671));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_A2 (.DIODE(net671));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_A0 (.DIODE(net671));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_C (.DIODE(net671));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_A2 (.DIODE(net671));
 sky130_fd_sc_hd__diode_2 ANTENNA_c180_B (.DIODE(net671));
 sky130_fd_sc_hd__diode_2 ANTENNA_input50_X (.DIODE(net672));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_A3 (.DIODE(net672));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_A0 (.DIODE(net672));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_B (.DIODE(net672));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_A3 (.DIODE(net672));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_B (.DIODE(net672));
 sky130_fd_sc_hd__diode_2 ANTENNA_c208_A2 (.DIODE(net672));
 sky130_fd_sc_hd__diode_2 ANTENNA_input51_X (.DIODE(net673));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_A2 (.DIODE(net673));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_C_N (.DIODE(net673));
 sky130_fd_sc_hd__diode_2 ANTENNA_c256_A2 (.DIODE(net673));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_A3 (.DIODE(net673));
 sky130_fd_sc_hd__diode_2 ANTENNA_c102_A1 (.DIODE(net673));
 sky130_fd_sc_hd__diode_2 ANTENNA_input52_X (.DIODE(net674));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_A0 (.DIODE(net674));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_A2 (.DIODE(net674));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_C1 (.DIODE(net674));
 sky130_fd_sc_hd__diode_2 ANTENNA_c190_C (.DIODE(net674));
 sky130_fd_sc_hd__diode_2 ANTENNA_input55_X (.DIODE(net677));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_A0 (.DIODE(net677));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_S0 (.DIODE(net677));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_A2 (.DIODE(net677));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_C1 (.DIODE(net677));
 sky130_fd_sc_hd__diode_2 ANTENNA_input56_X (.DIODE(net678));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_A0 (.DIODE(net678));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_A1 (.DIODE(net678));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_A1 (.DIODE(net678));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_A0 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_S1 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_A0 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_S1 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_A3 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_A (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_input57_X (.DIODE(net679));
 sky130_fd_sc_hd__diode_2 ANTENNA_c546_B (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c412_A1 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c344_B1 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_B1 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_input59_X (.DIODE(net681));
 sky130_fd_sc_hd__diode_2 ANTENNA_c765_A0 (.DIODE(net681));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A1 (.DIODE(net681));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_A3 (.DIODE(net681));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_S0 (.DIODE(net681));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_C1 (.DIODE(net681));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_S1 (.DIODE(net681));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_B (.DIODE(net681));
 sky130_fd_sc_hd__diode_2 ANTENNA_input61_X (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA_c767_A0 (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_A3 (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_A1 (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_A2 (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_A2 (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_B1 (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_C (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_S0 (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_B (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA_input63_X (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_A3 (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_A0 (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_A2 (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_A0 (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_C1 (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_A (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_C (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_B1 (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA_input65_X (.DIODE(net687));
 sky130_fd_sc_hd__diode_2 ANTENNA_c344_D1 (.DIODE(net687));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_A (.DIODE(net687));
 sky130_fd_sc_hd__diode_2 ANTENNA_input66_X (.DIODE(net688));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_A1 (.DIODE(net688));
 sky130_fd_sc_hd__diode_2 ANTENNA_input68_X (.DIODE(net690));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_A3 (.DIODE(net690));
 sky130_fd_sc_hd__diode_2 ANTENNA_c427_A (.DIODE(net690));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_A2 (.DIODE(net690));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_B (.DIODE(net690));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_S0 (.DIODE(net690));
 sky130_fd_sc_hd__diode_2 ANTENNA_c272_A (.DIODE(net690));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_D1 (.DIODE(net690));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_A2 (.DIODE(net690));
 sky130_fd_sc_hd__diode_2 ANTENNA_input69_X (.DIODE(net691));
 sky130_fd_sc_hd__diode_2 ANTENNA_c613_A3 (.DIODE(net691));
 sky130_fd_sc_hd__diode_2 ANTENNA_c482_A0 (.DIODE(net691));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_B (.DIODE(net691));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_B (.DIODE(net691));
 sky130_fd_sc_hd__diode_2 ANTENNA_c107_B1 (.DIODE(net691));
 sky130_fd_sc_hd__diode_2 ANTENNA_input70_X (.DIODE(net692));
 sky130_fd_sc_hd__diode_2 ANTENNA_c764_A0 (.DIODE(net692));
 sky130_fd_sc_hd__diode_2 ANTENNA_c743_A2 (.DIODE(net692));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_C1 (.DIODE(net692));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_A1 (.DIODE(net692));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_A1 (.DIODE(net692));
 sky130_fd_sc_hd__diode_2 ANTENNA_input74_X (.DIODE(net696));
 sky130_fd_sc_hd__diode_2 ANTENNA_c368_B (.DIODE(net696));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_A (.DIODE(net696));
 sky130_fd_sc_hd__diode_2 ANTENNA_c350_B1 (.DIODE(net696));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_C (.DIODE(net696));
 sky130_fd_sc_hd__diode_2 ANTENNA_input75_X (.DIODE(net697));
 sky130_fd_sc_hd__diode_2 ANTENNA_c370_A (.DIODE(net697));
 sky130_fd_sc_hd__diode_2 ANTENNA_c241_B1 (.DIODE(net697));
 sky130_fd_sc_hd__diode_2 ANTENNA_c221_A2 (.DIODE(net697));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_A2 (.DIODE(net697));
 sky130_fd_sc_hd__diode_2 ANTENNA_input76_X (.DIODE(net698));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge796_S1 (.DIODE(net698));
 sky130_fd_sc_hd__diode_2 ANTENNA_c767_A1 (.DIODE(net698));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_A2 (.DIODE(net698));
 sky130_fd_sc_hd__diode_2 ANTENNA_c228_B (.DIODE(net698));
 sky130_fd_sc_hd__diode_2 ANTENNA_c203_B (.DIODE(net698));
 sky130_fd_sc_hd__diode_2 ANTENNA_input77_X (.DIODE(net699));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_A2 (.DIODE(net699));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_A2 (.DIODE(net699));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_C_N (.DIODE(net699));
 sky130_fd_sc_hd__diode_2 ANTENNA_c236_A3 (.DIODE(net699));
 sky130_fd_sc_hd__diode_2 ANTENNA_c121_A1 (.DIODE(net699));
 sky130_fd_sc_hd__diode_2 ANTENNA_input78_X (.DIODE(net700));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_A0 (.DIODE(net700));
 sky130_fd_sc_hd__diode_2 ANTENNA_c102_A3 (.DIODE(net700));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout221_A (.DIODE(net701));
 sky130_fd_sc_hd__diode_2 ANTENNA_input79_X (.DIODE(net701));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_A1 (.DIODE(net701));
 sky130_fd_sc_hd__diode_2 ANTENNA_c746_A1 (.DIODE(net701));
 sky130_fd_sc_hd__diode_2 ANTENNA_input80_X (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA_c766_A0 (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_S0 (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_S0 (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_A2 (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_B (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA_c101_B (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA_input82_X (.DIODE(net704));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_C (.DIODE(net704));
 sky130_fd_sc_hd__diode_2 ANTENNA_c122_B (.DIODE(net704));
 sky130_fd_sc_hd__diode_2 ANTENNA_c121_S0 (.DIODE(net704));
 sky130_fd_sc_hd__diode_2 ANTENNA_c112_B (.DIODE(net704));
 sky130_fd_sc_hd__diode_2 ANTENNA_input83_X (.DIODE(net705));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_A0 (.DIODE(net705));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_A2 (.DIODE(net705));
 sky130_fd_sc_hd__diode_2 ANTENNA_input84_X (.DIODE(net706));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_D_N (.DIODE(net706));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_C1 (.DIODE(net706));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_A (.DIODE(net706));
 sky130_fd_sc_hd__diode_2 ANTENNA_c231_C (.DIODE(net706));
 sky130_fd_sc_hd__diode_2 ANTENNA_input85_X (.DIODE(net707));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_B1 (.DIODE(net707));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_A1 (.DIODE(net707));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_C1 (.DIODE(net707));
 sky130_fd_sc_hd__diode_2 ANTENNA_input86_X (.DIODE(net708));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge794_A3 (.DIODE(net708));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_S0 (.DIODE(net708));
 sky130_fd_sc_hd__diode_2 ANTENNA_c212_A2 (.DIODE(net708));
 sky130_fd_sc_hd__diode_2 ANTENNA_input87_X (.DIODE(net709));
 sky130_fd_sc_hd__diode_2 ANTENNA_c613_A1 (.DIODE(net709));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_A3 (.DIODE(net709));
 sky130_fd_sc_hd__diode_2 ANTENNA_c482_A3 (.DIODE(net709));
 sky130_fd_sc_hd__diode_2 ANTENNA_c262_A3 (.DIODE(net709));
 sky130_fd_sc_hd__diode_2 ANTENNA_c216_C1 (.DIODE(net709));
 sky130_fd_sc_hd__diode_2 ANTENNA_input88_X (.DIODE(net710));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_A (.DIODE(net710));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_A3 (.DIODE(net710));
 sky130_fd_sc_hd__diode_2 ANTENNA_c109_A3 (.DIODE(net710));
 sky130_fd_sc_hd__diode_2 ANTENNA_input89_X (.DIODE(net711));
 sky130_fd_sc_hd__diode_2 ANTENNA_c229_B (.DIODE(net711));
 sky130_fd_sc_hd__diode_2 ANTENNA_c109_S0 (.DIODE(net711));
 sky130_fd_sc_hd__diode_2 ANTENNA_c104_A (.DIODE(net711));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout3_A (.DIODE(net712));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone10_A2 (.DIODE(net712));
 sky130_fd_sc_hd__diode_2 ANTENNA_input90_X (.DIODE(net712));
 sky130_fd_sc_hd__diode_2 ANTENNA_input91_X (.DIODE(net713));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_A1 (.DIODE(net713));
 sky130_fd_sc_hd__diode_2 ANTENNA_c369_B (.DIODE(net713));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_S1 (.DIODE(net713));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_C1 (.DIODE(net713));
 sky130_fd_sc_hd__diode_2 ANTENNA_c236_A1 (.DIODE(net713));
 sky130_fd_sc_hd__diode_2 ANTENNA_c232_C1 (.DIODE(net713));
 sky130_fd_sc_hd__diode_2 ANTENNA_c105_A (.DIODE(net713));
 sky130_fd_sc_hd__diode_2 ANTENNA_input93_X (.DIODE(net715));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_A (.DIODE(net715));
 sky130_fd_sc_hd__diode_2 ANTENNA_c100_B (.DIODE(net715));
 sky130_fd_sc_hd__diode_2 ANTENNA_input95_X (.DIODE(net717));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_A1 (.DIODE(net717));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_A2 (.DIODE(net717));
 sky130_fd_sc_hd__diode_2 ANTENNA_c106_A (.DIODE(net717));
 sky130_fd_sc_hd__diode_2 ANTENNA_c100_C (.DIODE(net717));
 sky130_fd_sc_hd__diode_2 ANTENNA_input97_X (.DIODE(net719));
 sky130_fd_sc_hd__diode_2 ANTENNA_c114_A (.DIODE(net719));
 sky130_fd_sc_hd__diode_2 ANTENNA_c109_S1 (.DIODE(net719));
 sky130_fd_sc_hd__diode_2 ANTENNA_c105_C_N (.DIODE(net719));
 sky130_fd_sc_hd__diode_2 ANTENNA_input100_X (.DIODE(net722));
 sky130_fd_sc_hd__diode_2 ANTENNA_c761_A3 (.DIODE(net722));
 sky130_fd_sc_hd__diode_2 ANTENNA_c759_A0 (.DIODE(net722));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_S0 (.DIODE(net722));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_A3 (.DIODE(net722));
 sky130_fd_sc_hd__diode_2 ANTENNA_c221_D1 (.DIODE(net722));
 sky130_fd_sc_hd__diode_2 ANTENNA_c103_D_N (.DIODE(net722));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_C1 (.DIODE(net723));
 sky130_fd_sc_hd__diode_2 ANTENNA_output101_A (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_S0 (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_A3 (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_S0 (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_B1 (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_A2 (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c633_A2 (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c555_B (.DIODE(net723));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_X (.DIODE(net723));
 sky130_fd_sc_hd__diode_2 ANTENNA_output102_A (.DIODE(net724));
 sky130_fd_sc_hd__diode_2 ANTENNA_c761_S0 (.DIODE(net724));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_A3 (.DIODE(net724));
 sky130_fd_sc_hd__diode_2 ANTENNA_c686_B1 (.DIODE(net724));
 sky130_fd_sc_hd__diode_2 ANTENNA_c675_B (.DIODE(net724));
 sky130_fd_sc_hd__diode_2 ANTENNA_c674_X (.DIODE(net724));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout194_A (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA_output103_A (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA_c767_S0 (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_X (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA_output104_A (.DIODE(net726));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_C1 (.DIODE(net726));
 sky130_fd_sc_hd__diode_2 ANTENNA_c664_B (.DIODE(net726));
 sky130_fd_sc_hd__diode_2 ANTENNA_c615_A3 (.DIODE(net726));
 sky130_fd_sc_hd__diode_2 ANTENNA_c540_X (.DIODE(net726));
 sky130_fd_sc_hd__diode_2 ANTENNA_output109_A (.DIODE(net731));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_S1 (.DIODE(net731));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_A2 (.DIODE(net731));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_B (.DIODE(net731));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_B (.DIODE(net731));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_A3 (.DIODE(net731));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_B1 (.DIODE(net731));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_A (.DIODE(net731));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_X (.DIODE(net731));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout186_A (.DIODE(net733));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_S0 (.DIODE(net733));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_X (.DIODE(net733));
 sky130_fd_sc_hd__diode_2 ANTENNA_output112_A (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge868_Q_N (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA_c633_S0 (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_S0 (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_S0 (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_D1 (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_C1 (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_S1 (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout182_A (.DIODE(net735));
 sky130_fd_sc_hd__diode_2 ANTENNA_output113_A (.DIODE(net735));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_X (.DIODE(net735));
 sky130_fd_sc_hd__diode_2 ANTENNA_output115_A (.DIODE(net737));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_S0 (.DIODE(net737));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_A2 (.DIODE(net737));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_A2 (.DIODE(net737));
 sky130_fd_sc_hd__diode_2 ANTENNA_c446_X (.DIODE(net737));
 sky130_fd_sc_hd__diode_2 ANTENNA_output116_A (.DIODE(net738));
 sky130_fd_sc_hd__diode_2 ANTENNA_c765_A3 (.DIODE(net738));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A2 (.DIODE(net738));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_A3 (.DIODE(net738));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_A1 (.DIODE(net738));
 sky130_fd_sc_hd__diode_2 ANTENNA_c672_B (.DIODE(net738));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_B1 (.DIODE(net738));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_S0 (.DIODE(net738));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_X (.DIODE(net738));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone40_A (.DIODE(net740));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer21_A (.DIODE(net740));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout195_A (.DIODE(net740));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_X (.DIODE(net740));
 sky130_fd_sc_hd__diode_2 ANTENNA_output121_A (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge876_Q (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_S0 (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_S1 (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_S0 (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_S1 (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_S1 (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_C (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA_c577_C (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA_output122_A (.DIODE(net744));
 sky130_fd_sc_hd__diode_2 ANTENNA_c763_S1 (.DIODE(net744));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_S0 (.DIODE(net744));
 sky130_fd_sc_hd__diode_2 ANTENNA_c696_B (.DIODE(net744));
 sky130_fd_sc_hd__diode_2 ANTENNA_c678_SET_B (.DIODE(net744));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_A3 (.DIODE(net744));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_D1 (.DIODE(net744));
 sky130_fd_sc_hd__diode_2 ANTENNA_c279_D_N (.DIODE(net744));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_A3 (.DIODE(net744));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_A1 (.DIODE(net744));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_X (.DIODE(net744));
 sky130_fd_sc_hd__diode_2 ANTENNA_output124_A (.DIODE(net746));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_A2 (.DIODE(net746));
 sky130_fd_sc_hd__diode_2 ANTENNA_c496_A2 (.DIODE(net746));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_S1 (.DIODE(net746));
 sky130_fd_sc_hd__diode_2 ANTENNA_c257_A0 (.DIODE(net746));
 sky130_fd_sc_hd__diode_2 ANTENNA_c205_X (.DIODE(net746));
 sky130_fd_sc_hd__diode_2 ANTENNA_output125_A (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA_c571_S0 (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_A1 (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_SCD (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA_c566_X (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA_output127_A (.DIODE(net749));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_S0 (.DIODE(net749));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_B1 (.DIODE(net749));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_A3 (.DIODE(net749));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_A2 (.DIODE(net749));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_X (.DIODE(net749));
 sky130_fd_sc_hd__diode_2 ANTENNA_output128_A (.DIODE(net750));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_A3 (.DIODE(net750));
 sky130_fd_sc_hd__diode_2 ANTENNA_c369_X (.DIODE(net750));
 sky130_fd_sc_hd__diode_2 ANTENNA_output129_A (.DIODE(net751));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_A2 (.DIODE(net751));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_X (.DIODE(net751));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout217_A (.DIODE(net753));
 sky130_fd_sc_hd__diode_2 ANTENNA_output131_A (.DIODE(net753));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge867_Q (.DIODE(net753));
 sky130_fd_sc_hd__diode_2 ANTENNA_c757_S1 (.DIODE(net753));
 sky130_fd_sc_hd__diode_2 ANTENNA_output132_A (.DIODE(net754));
 sky130_fd_sc_hd__diode_2 ANTENNA_c502_A1 (.DIODE(net754));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_A3 (.DIODE(net754));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_A0 (.DIODE(net754));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_X (.DIODE(net754));
 sky130_fd_sc_hd__diode_2 ANTENNA_output133_A (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge790_S0 (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_A2 (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_A2 (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_X (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA_output135_A (.DIODE(net757));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge797_S0 (.DIODE(net757));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_S0 (.DIODE(net757));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_C1 (.DIODE(net757));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_A2 (.DIODE(net757));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_A3 (.DIODE(net757));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_C (.DIODE(net757));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_C (.DIODE(net757));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_X (.DIODE(net757));
 sky130_fd_sc_hd__diode_2 ANTENNA_output136_A (.DIODE(net758));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_A2 (.DIODE(net758));
 sky130_fd_sc_hd__diode_2 ANTENNA_c108_C1 (.DIODE(net758));
 sky130_fd_sc_hd__diode_2 ANTENNA_c105_X (.DIODE(net758));
 sky130_fd_sc_hd__diode_2 ANTENNA_output137_A (.DIODE(net759));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge873_Q (.DIODE(net759));
 sky130_fd_sc_hd__diode_2 ANTENNA_c764_S0 (.DIODE(net759));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_S1 (.DIODE(net759));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_S1 (.DIODE(net759));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_A3 (.DIODE(net759));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_S0 (.DIODE(net759));
 sky130_fd_sc_hd__diode_2 ANTENNA_c615_S0 (.DIODE(net759));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_S1 (.DIODE(net759));
 sky130_fd_sc_hd__diode_2 ANTENNA_output138_A (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_A2 (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA_c183_A (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_A3 (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_A (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_A0 (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_A2 (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_X (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA_c537_B (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_output139_A (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge794_A2 (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_S1 (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_B (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_C (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_A (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_X (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_output140_A (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_S0 (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_A1 (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_A2 (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_X (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout192_A (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_A3 (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_C (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_X (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA_output143_A (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_A2 (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_c230_X (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_c407_A (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer34_A (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_output145_A (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge795_S1 (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_c446_C (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_c402_X (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_output148_A (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_A2 (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_B1 (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_S1 (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_A1 (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_B (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_S1 (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_C1 (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_B1 (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_X (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer62_A (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_A (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c264_A (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_S1 (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_B1 (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_X (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_output151_A (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_A2 (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_X (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA_output152_A (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_c258_A2 (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_c220_C (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_c103_X (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_output155_A (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_S0 (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_c269_B (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_c220_B (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_C (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_A0 (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_A (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_c134_X (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_output158_A (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_A1 (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_C_N (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_B (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_B (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_X (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA_output160_A (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_B1 (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_A2 (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_A0 (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_c191_X (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer5_A (.DIODE(net783));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer4_A (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_output161_A (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c403_A (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c366_A2 (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c265_B (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_A1 (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c148_X (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_output165_A (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_B (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c220_X (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout213_A (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_output169_A (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_c262_S0 (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_c112_X (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_output174_A (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_A3 (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_A1 (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_B (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA_c180_X (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_D1 (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA_output175_A (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_B (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_A3 (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_A (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA_c159_X (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA_output176_A (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA_c120_D1 (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA_c118_X (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net799_A (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge881_GCLK (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_A2 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout182_X (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_A2 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_A3 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_A1 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_S1 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_S0 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_D1 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_C_N (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_B1 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_C (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout183_X (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_A2 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_A1 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_A1 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_A3 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_S1 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_S0 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_A2 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_S0 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_A2 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_A1 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout185_X (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_A0 (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_c695_B (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_c669_C1 (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_c662_D1 (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_S0 (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_c582_C_N (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_C (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_C1 (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_c560_C_N (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_S0 (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout186_X (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_A1 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_C_N (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c216_A2 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_output111_A (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_D1 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c256_A3 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c235_B1 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_A2 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c218_C1 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_A1 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout188_X (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_A3 (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_A3 (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge792_A2 (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_c238_B (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_c235_D1 (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_c212_C1 (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_C1 (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_c208_S0 (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_S1 (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_A2 (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout189_X (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_S0 (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_B (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_S1 (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_c230_B (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_c241_D1 (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_c237_C1 (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_c235_A1 (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_C1 (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_c232_D1 (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_c229_C (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout190_X (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_A2 (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_A3 (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_S0 (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_A2 (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout189_A (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_C1 (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout191_X (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_A3 (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_A2 (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_output110_A (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_A2 (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_A2 (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_A1 (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_A2 (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_B1 (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_C (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout192_X (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_c369_C_N (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_D1 (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_D1 (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_output141_A (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_B1 (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_C (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_S1 (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_C1 (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_B (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_C_N (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout193_X (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_S1 (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_A3 (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_S1 (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_c687_B1 (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_S0 (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_B (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_c544_A3 (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_B (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_c321_B1 (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_A1 (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout194_X (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_A3 (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_D1 (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c701_A2 (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_S0 (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_A3 (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_S0 (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_A2 (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c373_A2 (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_C1 (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_C_N (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout195_X (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_c665_C (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_c662_C1 (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_S0 (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_c402_A1 (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_A2 (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout196_X (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c757_A0 (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c720_A3 (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_C (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c273_B (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c566_S0 (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c554_C (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_A3 (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c277_A (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c276_A (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_B1 (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout197_X (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_D1 (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_S1 (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge790_S1 (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_S1 (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_S1 (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_C (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_D1 (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_D_N (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_C (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_B (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout198_X (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_output126_A (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_S1 (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_S0 (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_D1 (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_S1 (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_S1 (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout197_A (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout199_X (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_RESET_B (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_c671_B (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_c399_A (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_c428_B (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_c411_S0 (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_A3 (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_c297_S1 (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_c283_C (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_c272_C (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_c271_A (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_B1 (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout201_X (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_c560_D_N (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_c558_D_N (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_c537_D_N (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_C (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_C (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_C (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout200_A (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_c232_A2 (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout202_X (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_A3 (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_A3 (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_S0 (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_D_N (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout201_A (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout203_X (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_output108_A (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_A3 (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_A2 (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_A2 (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_c671_C (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_c660_C_N (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_S1 (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_S0 (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout202_A (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout206_X (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_B1 (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_C (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_S1 (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_D_N (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_S1 (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout204_A (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout205_A (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout207_X (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_D_N (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_S1 (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_D1 (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_S1 (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_C (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_C1 (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c232_B1 (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_C1 (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_D1 (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_S1 (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout208_X (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge793_S1 (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_SET_B (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA_c693_D_N (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA_c685_D_N (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_D_N (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_A2 (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout206_A (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout207_A (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_S0 (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_D1 (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone108_A (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c143_A (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout210_X (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_S1 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_S0 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_C1 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_C (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_C1 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout209_A (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout211_X (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_S1 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_D1 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_B1 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c539_A (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c410_S0 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_D1 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout210_A (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer98_A (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer97_A (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout212_X (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_C1 (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout211_A (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout213_X (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c127_S1 (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c123_B (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c119_C (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c114_B (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c113_B (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c129_B (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c125_B1 (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c124_C (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c121_A3 (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c118_C (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout214_X (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_S1 (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_D1 (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_S1 (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_S0 (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_S0 (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_S1 (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA_c263_S1 (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA_c261_S1 (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA_c234_A (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA_c222_A (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire215_X (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_output179_A (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_S0 (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_S1 (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_S0 (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout216_X (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_S1 (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_c764_A3 (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_S1 (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_D_N (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_S1 (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_D_N (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_D1 (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_D1 (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_S1 (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_D_N (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout217_X (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c691_S0 (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_S1 (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c742_A3 (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c562_D_N (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_S1 (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_D1 (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_S1 (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_A (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_A (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_C (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout218_X (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_c340_A (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_c239_A (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_D_N (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_c215_A (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_C1 (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_c371_D_N (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_c350_D1 (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_C_N (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_S1 (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_A (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout219_X (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_c759_S1 (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_S0 (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_S1 (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_S1 (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_S0 (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout218_A (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout220_X (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_A (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_c216_D1 (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_S1 (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_D1 (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_C (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_A (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_c263_S0 (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_c257_S1 (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_c261_S0 (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_c228_C (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_c143_C (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout221_X (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_A3 (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_A3 (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_S0 (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge793_S0 (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A2 (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_SCE (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c670_C (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_A3 (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c286_C (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout222_X (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_S0 (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_A3 (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_A2 (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_D_N (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_B1 (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_A (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c275_C (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_C (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_C (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c106_C (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout223_X (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_S0 (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_A3 (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A2 (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_S0 (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_c691_A2 (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout224_X (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_S0 (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_A3 (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_A3 (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_c587_S1 (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_A2 (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_B (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_A1 (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_B (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_S0 (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_C_N (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_c134_C (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout225_X (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_c720_S0 (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_S0 (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_c685_C_N (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_A2 (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_S0 (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_A2 (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_S0 (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_S0 (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_A2 (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout226_X (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_c532_B (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_c530_A (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_D_N (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_C (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_B (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_3__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_2__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_1__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_0__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_X (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge836_CLK (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge839_CLK (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge867_GATE_N (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge868_GATE_N (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge869_GATE (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge875_GATE (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge881_CLK (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge883_CLK (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_0__f_clk_X (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge858_CLK (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge862_CLK (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge866_CLK (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge873_GATE_N (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge878_CLK (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge879_CLK (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s885_CLK (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_1__f_clk_X (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_CLK_N (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c677_CLK_N (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c678_CLK (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_CLK_N (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_CLK_N (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge812_CLK (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge816_CLK (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge829_CLK_N (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge838_CLK (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge840_CLK (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge872_GATE_N (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge876_GATE (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s886_CLK (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_2__f_clk_X (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge865_CLK (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge870_GATE (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge871_GATE_N (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge877_GATE (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge880_CLK (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge882_CLK (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s884_CLK (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s887_CLK (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_3__f_clk_X (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_S1 (.DIODE(clknet_1_1__leaf_net615));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_S0 (.DIODE(clknet_1_1__leaf_net615));
 sky130_fd_sc_hd__diode_2 ANTENNA_c764_S1 (.DIODE(clknet_1_1__leaf_net615));
 sky130_fd_sc_hd__diode_2 ANTENNA_c769_S0 (.DIODE(clknet_1_1__leaf_net615));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net615_X (.DIODE(clknet_1_1__leaf_net615));
 sky130_fd_sc_hd__diode_2 ANTENNA_c240_C (.DIODE(clknet_1_0__leaf_net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c323_S1 (.DIODE(clknet_1_0__leaf_net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_D1 (.DIODE(clknet_1_0__leaf_net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_D_N (.DIODE(clknet_1_0__leaf_net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_C (.DIODE(clknet_1_0__leaf_net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_D_N (.DIODE(clknet_1_0__leaf_net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_S1 (.DIODE(clknet_1_0__leaf_net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_D1 (.DIODE(clknet_1_0__leaf_net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_D1 (.DIODE(clknet_1_0__leaf_net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_S1 (.DIODE(clknet_1_0__leaf_net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_S1 (.DIODE(clknet_1_0__leaf_net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net799_X (.DIODE(clknet_1_0__leaf_net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c236_S1 (.DIODE(clknet_1_1__leaf_net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c237_D1 (.DIODE(clknet_1_1__leaf_net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_S1 (.DIODE(clknet_1_1__leaf_net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c368_C (.DIODE(clknet_1_1__leaf_net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_S1 (.DIODE(clknet_1_1__leaf_net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c494_S1 (.DIODE(clknet_1_1__leaf_net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_S1 (.DIODE(clknet_1_1__leaf_net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_output177_A (.DIODE(clknet_1_1__leaf_net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net799_X (.DIODE(clknet_1_1__leaf_net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c610_S0 (.DIODE(clknet_1_0__leaf_net255));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_A2 (.DIODE(clknet_1_0__leaf_net255));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net255_X (.DIODE(clknet_1_0__leaf_net255));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_S0 (.DIODE(clknet_1_0__leaf_net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_A3 (.DIODE(clknet_1_0__leaf_net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_D1 (.DIODE(clknet_1_0__leaf_net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_B1 (.DIODE(clknet_1_0__leaf_net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_B1 (.DIODE(clknet_1_0__leaf_net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_D1 (.DIODE(clknet_1_0__leaf_net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge790_A1 (.DIODE(clknet_1_0__leaf_net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge797_A0 (.DIODE(clknet_1_0__leaf_net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net162_X (.DIODE(clknet_1_0__leaf_net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c611_S0 (.DIODE(clknet_1_1__leaf_net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_SCD (.DIODE(clknet_1_1__leaf_net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A3 (.DIODE(clknet_1_1__leaf_net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c743_A1 (.DIODE(clknet_1_1__leaf_net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c745_A0 (.DIODE(clknet_1_1__leaf_net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net162_X (.DIODE(clknet_1_1__leaf_net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer2_A (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c747_A0 (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_A3 (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_C1 (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer1_X (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_output149_A (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_D1 (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_S0 (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_B1 (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_A1 (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone10_X (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_D1 (.DIODE(net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer12_A (.DIODE(net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_A2 (.DIODE(net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer11_X (.DIODE(net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_output181_A (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_c259_A3 (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer13_X (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_output118_A (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer21_X (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_A2 (.DIODE(net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge795_A1 (.DIODE(net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer22_X (.DIODE(net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer32_A (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_c660_D_N (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer31_X (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_c662_A1 (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_c679_D1 (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer37_X (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_c724_B1 (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_A1 (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_S1 (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_A3 (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer39_A (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone40_X (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_C (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_C1 (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c110_A (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer42_A (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c262_S1 (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone43_X (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer45_A (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_output105_A (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_A2 (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer44_X (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_output130_A (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer56_X (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_A0 (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer59_A (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_A2 (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer58_X (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_c260_S1 (.DIODE(net910));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer62_X (.DIODE(net910));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_A2 (.DIODE(net916));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer68_X (.DIODE(net916));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_A3 (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_B1 (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer74_A (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer73_X (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_output106_A (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer75_A (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_S0 (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer74_X (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_A2 (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_A1 (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer78_X (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_A (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer106_A (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_A3 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer105_X (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_S1 (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_c148_D_N (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_C1 (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_c158_D_N (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone10_S1 (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone108_X (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout2_X (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone10_S0 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_C (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_D_N (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_S1 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c270_B (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c159_D1 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_D1 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_S0 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_S0 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_C (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout3_X (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c237_A1 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_A1 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c126_A (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c124_B (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c120_C1 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c108_D1 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_B (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_B (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_A2 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_A3 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(net553));
 sky130_fd_sc_hd__mux4_1 clone1 (.A0(net24),
    .A1(net20),
    .A2(net23),
    .A3(net760),
    .S0(net19),
    .S1(net831),
    .X(net963));
 sky130_fd_sc_hd__dlygate4sd3_1 rebuffer10 (.A(net29),
    .X(net964));
 sky130_fd_sc_hd__mux4_1 clone11 (.A0(net21),
    .A1(net28),
    .A2(net817),
    .A3(net744),
    .S0(net25),
    .S1(net969),
    .X(net965));
 sky130_fd_sc_hd__mux4_1 clone12 (.A0(net20),
    .A1(net27),
    .A2(net962),
    .A3(net633),
    .S0(net961),
    .S1(net831),
    .X(net966));
 sky130_fd_sc_hd__and3_1 clone13 (.A(net961),
    .B(net18),
    .C(net761),
    .X(net967));
 sky130_fd_sc_hd__and2_1 clone14 (.A(net17),
    .B(net635),
    .X(net968));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer38 (.A(net771),
    .X(net969));
 sky130_fd_sc_hd__clkbuf_1 clone39 (.A(net740),
    .X(net970));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer40 (.A(net825),
    .X(net971));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer43 (.A(net971),
    .X(net972));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer108 (.A(net972),
    .X(net973));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer110 (.A(net973),
    .X(net974));
 sky130_fd_sc_hd__or4bb_1 clone111 (.A(net18),
    .B(net24),
    .C_N(net19),
    .D_N(net956),
    .X(net975));
 sky130_fd_sc_hd__clkdlybuf4s50_1 rebuffer112 (.A(net142),
    .X(net976));
 sky130_fd_sc_hd__dlygate4sd3_1 rebuffer113 (.A(net976),
    .X(net977));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer114 (.A(net976),
    .X(net978));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer115 (.A(net976),
    .X(net979));
 sky130_fd_sc_hd__and2_1 clone116 (.A(net848),
    .B(net633),
    .X(net980));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer117 (.A(net723),
    .X(net981));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer118 (.A(net981),
    .X(net982));
 sky130_fd_sc_hd__clkbuf_1 rebuffer119 (.A(net982),
    .X(net983));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer120 (.A(net983),
    .X(net984));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer121 (.A(net225),
    .X(net985));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer122 (.A(net985),
    .X(net986));
 sky130_fd_sc_hd__and3_1 clone123 (.A(net988),
    .B(net131),
    .C(net642),
    .X(net987));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer124 (.A(net136),
    .X(net988));
 sky130_fd_sc_hd__clkbuf_1 clone125 (.A(in6),
    .X(net989));
 sky130_fd_sc_hd__clkbuf_1 clone126 (.A(net834),
    .X(net990));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_536 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_412 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_354 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_451 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_478 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_322 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_359 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_455 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_468 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_506 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_299 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_507 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_526 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_459 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_490 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_482 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_272 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_219 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_191 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_454 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_227 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_219 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_527 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_547 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_507 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_340 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_544 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_555 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_395 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_507 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_582 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_5 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_242 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_260 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_394 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_497 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_507 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_551 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_158 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_563 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_256 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_5 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_488 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_235 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_163 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_508 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_288 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_507 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_5 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_494 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_507 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_272 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_456 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_459 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_423 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_438 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_191 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_443 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_283 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_617 ();
endmodule
