module netlist_1 (clk,
    in0,
    in1,
    in10,
    in11,
    in12,
    in13,
    in14,
    in15,
    in16,
    in17,
    in18,
    in19,
    in2,
    in20,
    in21,
    in22,
    in23,
    in24,
    in25,
    in26,
    in27,
    in28,
    in29,
    in3,
    in30,
    in31,
    in32,
    in33,
    in34,
    in35,
    in36,
    in37,
    in38,
    in39,
    in4,
    in40,
    in41,
    in42,
    in43,
    in44,
    in45,
    in46,
    in47,
    in48,
    in49,
    in5,
    in50,
    in51,
    in52,
    in53,
    in54,
    in55,
    in56,
    in57,
    in58,
    in59,
    in6,
    in60,
    in61,
    in62,
    in63,
    in64,
    in65,
    in66,
    in67,
    in68,
    in69,
    in7,
    in70,
    in71,
    in72,
    in73,
    in74,
    in75,
    in76,
    in77,
    in78,
    in79,
    in8,
    in80,
    in81,
    in82,
    in83,
    in84,
    in85,
    in86,
    in87,
    in88,
    in89,
    in9,
    in90,
    in91,
    in92,
    in93,
    in94,
    in95,
    in96,
    in97,
    in98,
    in99,
    out0,
    out1,
    out10,
    out11,
    out12,
    out13,
    out14,
    out15,
    out16,
    out17,
    out18,
    out19,
    out2,
    out20,
    out21,
    out22,
    out23,
    out24,
    out25,
    out26,
    out27,
    out28,
    out29,
    out3,
    out30,
    out31,
    out32,
    out33,
    out34,
    out35,
    out36,
    out37,
    out38,
    out39,
    out4,
    out40,
    out41,
    out42,
    out43,
    out44,
    out45,
    out46,
    out47,
    out48,
    out49,
    out5,
    out50,
    out51,
    out52,
    out53,
    out54,
    out55,
    out56,
    out57,
    out58,
    out59,
    out6,
    out60,
    out61,
    out62,
    out63,
    out64,
    out65,
    out66,
    out67,
    out68,
    out69,
    out7,
    out70,
    out71,
    out72,
    out73,
    out74,
    out75,
    out76,
    out77,
    out78,
    out79,
    out8,
    out80,
    out81,
    out82,
    out83,
    out84,
    out85,
    out86,
    out87,
    out88,
    out89,
    out9,
    out90,
    out91,
    out92,
    out93,
    out94,
    out95,
    out96,
    out97,
    out98,
    out99,
    rst);
 input clk;
 input in0;
 input in1;
 input in10;
 input in11;
 input in12;
 input in13;
 input in14;
 input in15;
 input in16;
 input in17;
 input in18;
 input in19;
 input in2;
 input in20;
 input in21;
 input in22;
 input in23;
 input in24;
 input in25;
 input in26;
 input in27;
 input in28;
 input in29;
 input in3;
 input in30;
 input in31;
 input in32;
 input in33;
 input in34;
 input in35;
 input in36;
 input in37;
 input in38;
 input in39;
 input in4;
 input in40;
 input in41;
 input in42;
 input in43;
 input in44;
 input in45;
 input in46;
 input in47;
 input in48;
 input in49;
 input in5;
 input in50;
 input in51;
 input in52;
 input in53;
 input in54;
 input in55;
 input in56;
 input in57;
 input in58;
 input in59;
 input in6;
 input in60;
 input in61;
 input in62;
 input in63;
 input in64;
 input in65;
 input in66;
 input in67;
 input in68;
 input in69;
 input in7;
 input in70;
 input in71;
 input in72;
 input in73;
 input in74;
 input in75;
 input in76;
 input in77;
 input in78;
 input in79;
 input in8;
 input in80;
 input in81;
 input in82;
 input in83;
 input in84;
 input in85;
 input in86;
 input in87;
 input in88;
 input in89;
 input in9;
 input in90;
 input in91;
 input in92;
 input in93;
 input in94;
 input in95;
 input in96;
 input in97;
 input in98;
 input in99;
 output out0;
 output out1;
 output out10;
 output out11;
 output out12;
 output out13;
 output out14;
 output out15;
 output out16;
 output out17;
 output out18;
 output out19;
 output out2;
 output out20;
 output out21;
 output out22;
 output out23;
 output out24;
 output out25;
 output out26;
 output out27;
 output out28;
 output out29;
 output out3;
 output out30;
 output out31;
 output out32;
 output out33;
 output out34;
 output out35;
 output out36;
 output out37;
 output out38;
 output out39;
 output out4;
 output out40;
 output out41;
 output out42;
 output out43;
 output out44;
 output out45;
 output out46;
 output out47;
 output out48;
 output out49;
 output out5;
 output out50;
 output out51;
 output out52;
 output out53;
 output out54;
 output out55;
 output out56;
 output out57;
 output out58;
 output out59;
 output out6;
 output out60;
 output out61;
 output out62;
 output out63;
 output out64;
 output out65;
 output out66;
 output out67;
 output out68;
 output out69;
 output out7;
 output out70;
 output out71;
 output out72;
 output out73;
 output out74;
 output out75;
 output out76;
 output out77;
 output out78;
 output out79;
 output out8;
 output out80;
 output out81;
 output out82;
 output out83;
 output out84;
 output out85;
 output out86;
 output out87;
 output out88;
 output out89;
 output out9;
 output out90;
 output out91;
 output out92;
 output out93;
 output out94;
 output out95;
 output out96;
 output out97;
 output out98;
 output out99;
 input rst;

 wire net0;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net618;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net63;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net64;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net65;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net66;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net67;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net68;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net69;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net592;
 wire net604;
 wire net609;
 wire net617;
 wire net619;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire clknet_leaf_0_clk;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire clknet_0_net680;
 wire clknet_1_0__leaf_net680;
 wire clknet_1_1__leaf_net680;
 wire clknet_0_net679;
 wire clknet_1_0__leaf_net679;
 wire clknet_1_1__leaf_net679;
 wire clknet_0_net663;
 wire clknet_1_0__leaf_net663;
 wire clknet_1_1__leaf_net663;
 wire clknet_0_net327;
 wire clknet_1_0__leaf_net327;
 wire clknet_1_1__leaf_net327;
 wire clknet_0_net662;
 wire clknet_1_0__leaf_net662;
 wire clknet_1_1__leaf_net662;
 wire clknet_0_net419;
 wire clknet_1_0__leaf_net419;
 wire clknet_1_1__leaf_net419;
 wire clknet_0_net454;
 wire clknet_1_0__leaf_net454;
 wire clknet_1_1__leaf_net454;
 wire clknet_0_net455;
 wire clknet_1_0__leaf_net455;
 wire clknet_1_1__leaf_net455;
 wire clknet_0_net433;
 wire clknet_1_0__leaf_net433;
 wire clknet_1_1__leaf_net433;
 wire clknet_0_net421;
 wire clknet_1_0__leaf_net421;
 wire clknet_1_1__leaf_net421;
 wire clknet_0_net530;
 wire clknet_1_0__leaf_net530;
 wire clknet_1_1__leaf_net530;
 wire clknet_0_net423;
 wire clknet_1_0__leaf_net423;
 wire clknet_1_1__leaf_net423;
 wire clknet_0_net309;
 wire clknet_1_0__leaf_net309;
 wire clknet_1_1__leaf_net309;
 wire clknet_0_net288;
 wire clknet_1_0__leaf_net288;
 wire clknet_1_1__leaf_net288;
 wire clknet_0_net289;
 wire clknet_1_0__leaf_net289;
 wire clknet_1_1__leaf_net289;
 wire clknet_0_net643;
 wire clknet_1_0__leaf_net643;
 wire clknet_1_1__leaf_net643;
 wire clknet_0_net170;
 wire clknet_1_0__leaf_net170;
 wire clknet_1_1__leaf_net170;
 wire clknet_0_net184;
 wire clknet_1_0__leaf_net184;
 wire clknet_1_1__leaf_net184;
 wire clknet_0_net178;
 wire clknet_1_0__leaf_net178;
 wire clknet_1_1__leaf_net178;
 wire clknet_0_net175;
 wire clknet_1_0__leaf_net175;
 wire clknet_1_1__leaf_net175;
 wire clknet_0_net174;
 wire clknet_1_0__leaf_net174;
 wire clknet_1_1__leaf_net174;
 wire clknet_0_net173;
 wire clknet_1_0__leaf_net173;
 wire clknet_1_1__leaf_net173;
 wire clknet_0_net206;
 wire clknet_1_0__leaf_net206;
 wire clknet_1_1__leaf_net206;
 wire clknet_0_net185;
 wire clknet_1_0__leaf_net185;
 wire clknet_1_1__leaf_net185;
 wire clknet_0_net642;
 wire clknet_1_0__leaf_net642;
 wire clknet_1_1__leaf_net642;
 wire clknet_0_net602;
 wire clknet_1_0__leaf_net602;
 wire clknet_1_1__leaf_net602;
 wire clknet_0_net105;
 wire clknet_1_0__leaf_net105;
 wire clknet_1_1__leaf_net105;
 wire clknet_0_net806;
 wire clknet_1_0__leaf_net806;
 wire clknet_1_1__leaf_net806;
 wire clknet_0_net102;
 wire clknet_1_0__leaf_net102;
 wire clknet_1_1__leaf_net102;
 wire clknet_0_net106;
 wire clknet_1_0__leaf_net106;
 wire clknet_1_1__leaf_net106;
 wire clknet_0_net113;
 wire clknet_1_0__leaf_net113;
 wire clknet_1_1__leaf_net113;
 wire clknet_0_net111;
 wire clknet_1_0__leaf_net111;
 wire clknet_1_1__leaf_net111;
 wire clknet_0_net112;
 wire clknet_1_0__leaf_net112;
 wire clknet_1_1__leaf_net112;
 wire clknet_0_net108;
 wire clknet_1_0__leaf_net108;
 wire clknet_1_1__leaf_net108;
 wire clknet_0_net118;
 wire clknet_1_0__leaf_net118;
 wire clknet_1_1__leaf_net118;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;

 sky130_fd_sc_hd__mux4_1 c100 (.A0(net764),
    .A1(net778),
    .A2(net784),
    .A3(net773),
    .S0(net787),
    .S1(net780),
    .X(net0));
 sky130_fd_sc_hd__mux4_1 c101 (.A0(net788),
    .A1(net783),
    .A2(net780),
    .A3(net786),
    .S0(net759),
    .S1(net787),
    .X(net1));
 sky130_fd_sc_hd__mux4_1 c102 (.A0(net767),
    .A1(net777),
    .A2(net789),
    .A3(net776),
    .S0(net783),
    .S1(net780),
    .X(net2));
 sky130_fd_sc_hd__mux4_2 c103 (.A0(net785),
    .A1(net0),
    .A2(net787),
    .A3(net1),
    .S0(net2),
    .S1(net783),
    .X(net811));
 sky130_fd_sc_hd__mux4_1 c104 (.A0(net775),
    .A1(net774),
    .A2(net781),
    .A3(net782),
    .S0(net780),
    .S1(net787),
    .X(net3));
 sky130_fd_sc_hd__dlymetal6s2s_1 c121 (.A(net3),
    .X(net807));
 sky130_fd_sc_hd__clkbuf_1 c122 (.A(net807),
    .X(net817));
 sky130_fd_sc_hd__clkbuf_1 c123 (.X(net818));
 sky130_fd_sc_hd__clkbuf_1 c124 (.A(net591),
    .X(net814));
 sky130_fd_sc_hd__sdfrbp_1 c125 (.CLK(clknet_leaf_34_clk),
    .D(net818),
    .RESET_B(net807),
    .SCD(net817),
    .SCE(net814),
    .Q(net815),
    .Q_N(net816));
 sky130_fd_sc_hd__and2_1 c126 (.A(net747),
    .B(net699),
    .X(net4));
 sky130_fd_sc_hd__and2_1 c127 (.A(net4),
    .B(net696),
    .X(net5));
 sky130_fd_sc_hd__and3_1 c128 (.A(net5),
    .B(net619),
    .C(net700),
    .X(net6));
 sky130_fd_sc_hd__and3_1 c129 (.A(net4),
    .B(net609),
    .C(net5),
    .X(net7));
 sky130_fd_sc_hd__buf_1 c130 (.A(net611),
    .X(net8));
 sky130_fd_sc_hd__buf_1 c131 (.A(net611),
    .X(net9));
 sky130_fd_sc_hd__dfbbn_1 c132 (.CLK_N(clknet_leaf_9_clk),
    .D(net5),
    .RESET_B(net7),
    .SET_B(net9),
    .Q(net11),
    .Q_N(net10));
 sky130_fd_sc_hd__and3_1 c133 (.A(net714),
    .B(net4),
    .C(net736),
    .X(net12));
 sky130_fd_sc_hd__dfbbn_1 c134 (.CLK_N(clknet_leaf_9_clk),
    .D(net8),
    .RESET_B(net6),
    .SET_B(net869),
    .Q(net14),
    .Q_N(net13));
 sky130_fd_sc_hd__and3_1 c135 (.A(net11),
    .B(net14),
    .C(net4),
    .X(net15));
 sky130_fd_sc_hd__or4bb_1 c136 (.A(net12),
    .B(net15),
    .C_N(net4),
    .D_N(net758),
    .X(net16));
 sky130_fd_sc_hd__sdfbbn_1 c137 (.CLK_N(clknet_leaf_9_clk),
    .D(net16),
    .RESET_B(net604),
    .SCD(net911),
    .SCE(net779),
    .SET_B(net701),
    .Q(net18),
    .Q_N(net17));
 sky130_fd_sc_hd__a2111o_1 c138 (.A1(net9),
    .A2(net698),
    .B1(net17),
    .C1(net704),
    .D1(net8),
    .X(net19));
 sky130_fd_sc_hd__dfbbp_1 c139 (.CLK(clknet_leaf_9_clk),
    .D(net18),
    .RESET_B(net592),
    .SET_B(net16),
    .Q(net20));
 sky130_fd_sc_hd__sdfbbn_1 c140 (.CLK_N(clknet_leaf_8_clk),
    .D(net6),
    .RESET_B(net856),
    .SCD(net15),
    .SCE(net703),
    .SET_B(net8),
    .Q(net22),
    .Q_N(net21));
 sky130_fd_sc_hd__and3_1 c141 (.A(net14),
    .B(net20),
    .C(net22),
    .X(net23));
 sky130_fd_sc_hd__and3_1 c142 (.A(net725),
    .B(net15),
    .C(net21),
    .X(net24));
 sky130_fd_sc_hd__mux4_1 c143 (.A0(net19),
    .A1(net22),
    .A2(net24),
    .A3(net697),
    .S0(net5),
    .S1(net17),
    .X(net25));
 sky130_fd_sc_hd__sdfbbp_1 c144 (.CLK(clknet_leaf_8_clk),
    .D(net702),
    .RESET_B(net23),
    .SCD(net6),
    .SCE(net21),
    .SET_B(net845),
    .Q(net26));
 sky130_fd_sc_hd__sdfxbp_1 c145 (.CLK(clknet_leaf_8_clk),
    .D(net22),
    .SCD(net24),
    .SCE(net879),
    .Q(net27));
 sky130_fd_sc_hd__mux4_1 c146 (.A0(net26),
    .A1(net27),
    .A2(net15),
    .A3(net18),
    .S0(net19),
    .S1(net635),
    .X(net28));
 sky130_fd_sc_hd__and2_1 c147 (.A(net617),
    .B(net719),
    .X(net29));
 sky130_fd_sc_hd__and2_0 c148 (.A(net709),
    .B(net711),
    .X(net30));
 sky130_fd_sc_hd__and2_1 c149 (.A(net722),
    .B(net724),
    .X(net31));
 sky130_fd_sc_hd__and3_1 c150 (.A(net29),
    .B(net30),
    .C(net716),
    .X(net32));
 sky130_fd_sc_hd__and3_1 c151 (.A(net32),
    .B(net29),
    .C(net726),
    .X(net33));
 sky130_fd_sc_hd__and2_1 c152 (.A(net30),
    .B(net32),
    .X(net34));
 sky130_fd_sc_hd__sdfbbn_1 c153 (.CLK_N(clknet_leaf_0_clk),
    .D(net819),
    .RESET_B(net33),
    .SCD(net712),
    .SCE(net706),
    .SET_B(net32),
    .Q(net36),
    .Q_N(net35));
 sky130_fd_sc_hd__buf_1 c154 (.A(net598),
    .X(net37));
 sky130_fd_sc_hd__sdfxbp_1 c155 (.CLK(clknet_leaf_6_clk),
    .D(net31),
    .SCD(net37),
    .SCE(net819),
    .Q(net39),
    .Q_N(net38));
 sky130_fd_sc_hd__sdfxtp_1 c156 (.CLK(clknet_leaf_6_clk),
    .D(net723),
    .SCD(net862),
    .SCE(net819),
    .Q(net40));
 sky130_fd_sc_hd__buf_1 c157 (.A(net827),
    .X(net41));
 sky130_fd_sc_hd__sdfxtp_1 c158 (.CLK(clknet_leaf_6_clk),
    .D(net720),
    .SCD(net885),
    .SCE(net819),
    .Q(net42));
 sky130_fd_sc_hd__and3_1 c159 (.A(net40),
    .B(net42),
    .C(net31),
    .X(net43));
 sky130_fd_sc_hd__sdfbbn_1 c160 (.CLK_N(clknet_leaf_35_clk),
    .D(net30),
    .RESET_B(net40),
    .SCD(net41),
    .SCE(net819),
    .SET_B(net42),
    .Q(net45),
    .Q_N(net44));
 sky130_fd_sc_hd__sdfrbp_1 c161 (.CLK(clknet_leaf_6_clk),
    .D(net45),
    .RESET_B(net41),
    .SCD(net40),
    .SCE(net819),
    .Q(net47),
    .Q_N(net46));
 sky130_fd_sc_hd__mux4_1 c162 (.A0(net39),
    .A1(net33),
    .A2(net705),
    .A3(net47),
    .S0(net721),
    .S1(net819),
    .X(net48));
 sky130_fd_sc_hd__sdfbbp_1 c163 (.CLK(clknet_leaf_6_clk),
    .D(net859),
    .RESET_B(net885),
    .SCD(net43),
    .SCE(net34),
    .SET_B(net830),
    .Q(net50),
    .Q_N(net49));
 sky130_fd_sc_hd__mux4_1 c164 (.A0(net36),
    .A1(net37),
    .A2(net45),
    .A3(net713),
    .S0(net50),
    .S1(net819),
    .X(net51));
 sky130_fd_sc_hd__mux4_1 c165 (.A0(net43),
    .A1(net50),
    .A2(net42),
    .A3(net35),
    .S0(net637),
    .S1(net639),
    .X(net52));
 sky130_fd_sc_hd__mux4_1 c166 (.A0(net708),
    .A1(net44),
    .A2(net52),
    .A3(net819),
    .S0(net32),
    .S1(net830),
    .X(net53));
 sky130_fd_sc_hd__mux4_1 c167 (.A0(net52),
    .A1(net40),
    .A2(net46),
    .A3(net49),
    .S0(net639),
    .S1(net875),
    .X(net54));
 sky130_fd_sc_hd__and2_1 c168 (.A(net718),
    .B(net740),
    .X(net55));
 sky130_fd_sc_hd__and3_2 c169 (.A(net727),
    .B(net731),
    .C(net733),
    .X(net56));
 sky130_fd_sc_hd__and3_1 c170 (.A(net56),
    .B(net746),
    .C(net743),
    .X(net57));
 sky130_fd_sc_hd__and2_0 c171 (.A(net745),
    .B(net56),
    .X(net58));
 sky130_fd_sc_hd__and3_1 c172 (.A(net37),
    .B(net56),
    .C(net750),
    .X(net59));
 sky130_fd_sc_hd__a2111o_1 c173 (.A1(net55),
    .A2(net744),
    .B1(net56),
    .C1(net748),
    .D1(net729),
    .X(net60));
 sky130_fd_sc_hd__and3_1 c174 (.A(net59),
    .B(net56),
    .C(net741),
    .X(net61));
 sky130_fd_sc_hd__and3_1 c175 (.A(net58),
    .B(net56),
    .C(net60),
    .X(net62));
 sky130_fd_sc_hd__and3_1 c176 (.A(net32),
    .B(net56),
    .C(net57),
    .X(net63));
 sky130_fd_sc_hd__buf_1 c177 (.A(net695),
    .X(net64));
 sky130_fd_sc_hd__and3_1 c178 (.A(net29),
    .B(net57),
    .C(net64),
    .X(net65));
 sky130_fd_sc_hd__and2_0 c179 (.A(net60),
    .B(net64),
    .X(net66));
 sky130_fd_sc_hd__mux4_1 c180 (.A0(net64),
    .A1(net66),
    .A2(net63),
    .A3(net55),
    .S0(net61),
    .S1(net56),
    .X(net67));
 sky130_fd_sc_hd__buf_1 c181 (.A(net695),
    .X(net68));
 sky130_fd_sc_hd__and3_1 c182 (.A(net57),
    .B(net68),
    .C(clknet_1_1__leaf_net642),
    .X(net69));
 sky130_fd_sc_hd__and3_1 c183 (.A(net734),
    .B(net55),
    .C(net749),
    .X(net70));
 sky130_fd_sc_hd__sdfxtp_1 c184 (.CLK(clknet_leaf_35_clk),
    .D(net65),
    .SCD(net68),
    .SCE(net70),
    .Q(net71));
 sky130_fd_sc_hd__dfbbn_1 c185 (.CLK_N(clknet_leaf_35_clk),
    .D(net71),
    .RESET_B(net64),
    .SET_B(net63),
    .Q(net72));
 sky130_fd_sc_hd__mux4_1 c186 (.A0(net69),
    .A1(net70),
    .A2(net66),
    .A3(net728),
    .S0(net738),
    .S1(clknet_1_0__leaf_net642),
    .X(net73));
 sky130_fd_sc_hd__and3_1 c187 (.A(net68),
    .B(net72),
    .C(clknet_1_0__leaf_net643),
    .X(net74));
 sky130_fd_sc_hd__mux4_1 c188 (.A0(net74),
    .A1(net70),
    .A2(net64),
    .A3(net732),
    .S0(net735),
    .S1(clknet_1_0__leaf_net643),
    .X(net75));
 sky130_fd_sc_hd__and2_2 c189 (.A(net762),
    .B(net730),
    .X(net76));
 sky130_fd_sc_hd__and2_1 c190 (.A(net76),
    .B(net766),
    .X(net77));
 sky130_fd_sc_hd__and3_1 c191 (.A(net77),
    .B(net757),
    .C(net771),
    .X(net78));
 sky130_fd_sc_hd__and2_1 c192 (.A(net77),
    .B(net76),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_1 c193 (.A(net623),
    .X(net80));
 sky130_fd_sc_hd__clkbuf_1 c194 (.A(net622),
    .X(net81));
 sky130_fd_sc_hd__and3_1 c195 (.A(net76),
    .B(net81),
    .C(net769),
    .X(net82));
 sky130_fd_sc_hd__dfrbp_1 c196 (.CLK(clknet_leaf_33_clk),
    .D(net82),
    .RESET_B(net78),
    .Q(net84),
    .Q_N(net83));
 sky130_fd_sc_hd__and3_1 c197 (.A(net81),
    .B(net84),
    .C(net756),
    .X(net85));
 sky130_fd_sc_hd__buf_1 c198 (.A(net631),
    .X(net86));
 sky130_fd_sc_hd__sdfbbn_1 c199 (.CLK_N(clknet_leaf_33_clk),
    .D(net751),
    .RESET_B(net79),
    .SCD(net76),
    .SCE(net86),
    .SET_B(net78),
    .Q(net88),
    .Q_N(net87));
 sky130_fd_sc_hd__mux4_2 c200 (.A0(net88),
    .A1(net754),
    .A2(net86),
    .A3(net76),
    .S0(net84),
    .S1(net80),
    .X(net89));
 sky130_fd_sc_hd__and2_0 c201 (.A(net77),
    .B(net82),
    .X(net90));
 sky130_fd_sc_hd__sdfbbn_1 c202 (.CLK_N(clknet_leaf_33_clk),
    .D(net89),
    .RESET_B(net79),
    .SCD(net76),
    .SCE(net83),
    .SET_B(net761),
    .Q(net92),
    .Q_N(net91));
 sky130_fd_sc_hd__or4bb_4 c203 (.A(net84),
    .B(net89),
    .C_N(net86),
    .D_N(net772),
    .X(net93));
 sky130_fd_sc_hd__dfbbn_1 c204 (.CLK_N(clknet_leaf_32_clk),
    .D(net80),
    .RESET_B(net90),
    .SET_B(net83),
    .Q(net95),
    .Q_N(net94));
 sky130_fd_sc_hd__mux4_1 c205 (.A0(net95),
    .A1(net822),
    .A2(net77),
    .A3(net752),
    .S0(net85),
    .S1(net770),
    .X(net96));
 sky130_fd_sc_hd__and3_1 c206 (.A(net92),
    .B(net87),
    .C(net86),
    .X(net97));
 sky130_fd_sc_hd__mux4_1 c207 (.A0(net97),
    .A1(net94),
    .A2(net84),
    .A3(net76),
    .S0(net91),
    .S1(net763),
    .X(net98));
 sky130_fd_sc_hd__mux4_1 c208 (.A0(net93),
    .A1(net96),
    .A2(net97),
    .A3(net98),
    .S0(net78),
    .S1(net822),
    .X(net99));
 sky130_fd_sc_hd__dfbbp_1 c209 (.CLK(clknet_leaf_32_clk),
    .D(net98),
    .RESET_B(net93),
    .SET_B(net644),
    .Q(net100));
 sky130_fd_sc_hd__buf_1 c210 (.A(net811),
    .X(net101));
 sky130_fd_sc_hd__buf_1 c211 (.A(clknet_1_0__leaf_net602),
    .X(net102));
 sky130_fd_sc_hd__sdfxbp_1 c212 (.CLK(clknet_leaf_27_clk),
    .D(net86),
    .SCD(net101),
    .SCE(clknet_1_0__leaf_net102),
    .Q(net104),
    .Q_N(net103));
 sky130_fd_sc_hd__buf_1 c213 (.A(clknet_1_1__leaf_net602),
    .X(net105));
 sky130_fd_sc_hd__and2_0 c214 (.A(net760),
    .B(clknet_1_0__leaf_net102),
    .X(net106));
 sky130_fd_sc_hd__buf_1 c215 (.A(net632),
    .X(net107));
 sky130_fd_sc_hd__and2_0 c216 (.A(clknet_1_0__leaf_net106),
    .B(net107),
    .X(net108));
 sky130_fd_sc_hd__dfrbp_1 c217 (.CLK(clknet_leaf_28_clk),
    .D(clknet_1_0__leaf_net108),
    .RESET_B(net101),
    .Q(net110),
    .Q_N(net109));
 sky130_fd_sc_hd__and2_0 c218 (.A(clknet_1_1__leaf_net106),
    .B(net109),
    .X(net111));
 sky130_fd_sc_hd__and3_1 c219 (.A(net107),
    .B(clknet_1_1__leaf_net108),
    .C(clknet_1_0__leaf_net111),
    .X(net112));
 sky130_fd_sc_hd__and3_1 c220 (.A(clknet_1_0__leaf_net108),
    .B(clknet_1_0__leaf_net106),
    .C(clknet_1_0__leaf_net111),
    .X(net113));
 sky130_fd_sc_hd__dfrtn_1 c221 (.CLK_N(clknet_leaf_28_clk),
    .D(clknet_1_1__leaf_net113),
    .RESET_B(clknet_1_0__leaf_net112),
    .Q(net114));
 sky130_fd_sc_hd__sdfxbp_1 c222 (.CLK(clknet_leaf_26_clk),
    .D(clknet_1_1__leaf_net111),
    .SCD(clknet_1_1__leaf_net102),
    .SCE(clknet_1_0__leaf_net112),
    .Q(net808),
    .Q_N(net115));
 sky130_fd_sc_hd__mux4_1 c223 (.A0(net110),
    .A1(net114),
    .A2(clknet_1_0__leaf_net105),
    .A3(clknet_1_0__leaf_net112),
    .S0(clknet_1_0__leaf_net111),
    .S1(clknet_1_1__leaf_net108),
    .X(net116));
 sky130_fd_sc_hd__and2_1 c224 (.A(net114),
    .B(net808),
    .X(net117));
 sky130_fd_sc_hd__and3_1 c225 (.A(net104),
    .B(clknet_1_1__leaf_net108),
    .C(net114),
    .X(net118));
 sky130_fd_sc_hd__sdfxtp_1 c226 (.CLK(clknet_leaf_27_clk),
    .D(net903),
    .SCD(clknet_1_0__leaf_net118),
    .SCE(clknet_1_1__leaf_net102),
    .Q(net119));
 sky130_fd_sc_hd__sdfbbp_1 c227 (.CLK(clknet_leaf_27_clk),
    .D(clknet_1_0__leaf_net112),
    .RESET_B(net117),
    .SCD(clknet_1_0__leaf_net113),
    .SCE(clknet_1_0__leaf_net111),
    .SET_B(net831),
    .Q(net121),
    .Q_N(net120));
 sky130_fd_sc_hd__sdfrtn_1 c228 (.CLK_N(clknet_leaf_27_clk),
    .D(clknet_1_1__leaf_net118),
    .RESET_B(net825),
    .SCD(net119),
    .SCE(net120),
    .Q(net813));
 sky130_fd_sc_hd__a2111o_1 c229 (.A1(clknet_1_1__leaf_net105),
    .A2(net121),
    .B1(net117),
    .C1(net115),
    .D1(net813),
    .X(net806));
 sky130_fd_sc_hd__sdfrtp_1 c230 (.CLK(clknet_leaf_27_clk),
    .D(net831),
    .RESET_B(clknet_1_1__leaf_net112),
    .SCD(net121),
    .SCE(clknet_1_1__leaf_net806),
    .Q(net809));
 sky130_fd_sc_hd__buf_2 c252 (.X(net122));
 sky130_fd_sc_hd__clkbuf_1 c253 (.A(net820),
    .X(net123));
 sky130_fd_sc_hd__and2_1 c254 (.A(net123),
    .B(net820),
    .X(net124));
 sky130_fd_sc_hd__and2_0 c255 (.A(net820),
    .B(net124),
    .X(net125));
 sky130_fd_sc_hd__and2_1 c256 (.A(net123),
    .B(net820),
    .X(net126));
 sky130_fd_sc_hd__clkbuf_2 c257 (.A(net603),
    .X(net127));
 sky130_fd_sc_hd__and3_1 c258 (.A(net820),
    .B(net127),
    .C(net126),
    .X(net128));
 sky130_fd_sc_hd__and2_0 c259 (.A(net127),
    .B(net820),
    .X(net129));
 sky130_fd_sc_hd__sdfxtp_1 c260 (.CLK(clknet_leaf_6_clk),
    .D(net128),
    .SCD(net820),
    .SCE(net124),
    .Q(net130));
 sky130_fd_sc_hd__sdfxtp_1 c261 (.CLK(clknet_leaf_7_clk),
    .D(net909),
    .SCD(net128),
    .SCE(net127),
    .Q(net131));
 sky130_fd_sc_hd__sdfrtp_1 c262 (.CLK(clknet_leaf_8_clk),
    .D(net125),
    .RESET_B(net127),
    .SCD(net129),
    .SCE(net820),
    .Q(net132));
 sky130_fd_sc_hd__and3_1 c263 (.A(net131),
    .B(net132),
    .C(net130),
    .X(net133));
 sky130_fd_sc_hd__and3_1 c264 (.A(net133),
    .B(net131),
    .C(net820),
    .X(net134));
 sky130_fd_sc_hd__and3_1 c265 (.A(net134),
    .B(net133),
    .C(net130),
    .X(net135));
 sky130_fd_sc_hd__mux4_1 c266 (.A0(net132),
    .A1(net134),
    .A2(net130),
    .A3(net820),
    .S0(net127),
    .S1(net131),
    .X(net136));
 sky130_fd_sc_hd__dfbbn_1 c267 (.CLK_N(clknet_leaf_6_clk),
    .D(net124),
    .RESET_B(net135),
    .SET_B(net821),
    .Q(net138),
    .Q_N(net137));
 sky130_fd_sc_hd__mux4_1 c268 (.A0(net126),
    .A1(net136),
    .A2(net137),
    .A3(net135),
    .S0(net130),
    .S1(net134),
    .X(net139));
 sky130_fd_sc_hd__mux4_1 c269 (.A0(net129),
    .A1(net138),
    .A2(net821),
    .A3(net134),
    .S0(net130),
    .S1(net645),
    .X(net140));
 sky130_fd_sc_hd__sdfbbn_1 c270 (.CLK_N(clknet_leaf_7_clk),
    .D(net140),
    .RESET_B(net874),
    .SCD(net136),
    .SCE(net821),
    .SET_B(net841),
    .Q(net142),
    .Q_N(net141));
 sky130_fd_sc_hd__mux4_1 c271 (.A0(net138),
    .A1(net136),
    .A2(net133),
    .A3(net141),
    .S0(net126),
    .S1(net821),
    .X(net143));
 sky130_fd_sc_hd__a2111o_1 c272 (.A1(net142),
    .A2(net127),
    .B1(net821),
    .C1(net646),
    .D1(net647),
    .X(net144));
 sky130_fd_sc_hd__and2_2 c273 (.A(net715),
    .B(net641),
    .X(net145));
 sky130_fd_sc_hd__and2_2 c274 (.A(net31),
    .B(net145),
    .X(net146));
 sky130_fd_sc_hd__and2_1 c275 (.A(net717),
    .B(net146),
    .X(net147));
 sky130_fd_sc_hd__clkbuf_2 c276 (.X(net148));
 sky130_fd_sc_hd__and2_0 c277 (.A(net146),
    .B(net148),
    .X(net149));
 sky130_fd_sc_hd__dfbbn_1 c278 (.CLK_N(clknet_leaf_5_clk),
    .D(net149),
    .RESET_B(net146),
    .SET_B(net148),
    .Q(net151),
    .Q_N(net150));
 sky130_fd_sc_hd__and3_1 c279 (.A(net148),
    .B(net146),
    .C(net145),
    .X(net152));
 sky130_fd_sc_hd__and2_0 c280 (.A(net151),
    .B(net145),
    .X(net153));
 sky130_fd_sc_hd__and2_0 c281 (.A(net145),
    .B(net146),
    .X(net154));
 sky130_fd_sc_hd__sdfrtp_1 c282 (.CLK(clknet_leaf_5_clk),
    .D(net153),
    .RESET_B(net147),
    .SCD(net710),
    .SCE(net146),
    .Q(net155));
 sky130_fd_sc_hd__dfbbp_1 c283 (.CLK(clknet_leaf_5_clk),
    .D(net147),
    .RESET_B(net866),
    .SET_B(net832),
    .Q(net157),
    .Q_N(net156));
 sky130_fd_sc_hd__sdfbbn_1 c284 (.CLK_N(clknet_leaf_5_clk),
    .D(net146),
    .RESET_B(net145),
    .SCD(net148),
    .SCE(net150),
    .SET_B(net152),
    .Q(net159),
    .Q_N(net158));
 sky130_fd_sc_hd__and2_1 c285 (.A(net157),
    .B(net159),
    .X(net160));
 sky130_fd_sc_hd__mux4_1 c286 (.A0(net160),
    .A1(net158),
    .A2(net155),
    .A3(net147),
    .S0(net152),
    .S1(net145),
    .X(net161));
 sky130_fd_sc_hd__sdfxbp_1 c287 (.CLK(clknet_leaf_0_clk),
    .D(net154),
    .SCD(net152),
    .SCE(net160),
    .Q(net163),
    .Q_N(net162));
 sky130_fd_sc_hd__and3_1 c288 (.A(net155),
    .B(net160),
    .C(net148),
    .X(net164));
 sky130_fd_sc_hd__clkbuf_1 c289 (.A(net618),
    .X(net165));
 sky130_fd_sc_hd__mux4_1 c290 (.A0(net165),
    .A1(net155),
    .A2(net156),
    .A3(net148),
    .S0(net145),
    .S1(net649),
    .X(net166));
 sky130_fd_sc_hd__mux4_1 c291 (.A0(net163),
    .A1(net166),
    .A2(net160),
    .A3(net151),
    .S0(net145),
    .S1(net148),
    .X(net167));
 sky130_fd_sc_hd__sdfxbp_1 c292 (.CLK(clknet_leaf_1_clk),
    .D(net164),
    .SCD(net167),
    .SCE(net908),
    .Q(net168));
 sky130_fd_sc_hd__sdfxtp_1 c293 (.CLK(clknet_leaf_1_clk),
    .D(net152),
    .SCD(net847),
    .SCE(net160),
    .Q(net169));
 sky130_fd_sc_hd__and2_0 c294 (.A(net742),
    .B(clknet_1_1__leaf_net643),
    .X(net170));
 sky130_fd_sc_hd__clkbuf_1 c295 (.A(net601),
    .X(net171));
 sky130_fd_sc_hd__and2_2 c296 (.A(net171),
    .B(net739),
    .X(net172));
 sky130_fd_sc_hd__and2_0 c297 (.A(net172),
    .B(clknet_1_1__leaf_net170),
    .X(net173));
 sky130_fd_sc_hd__and2_0 c298 (.A(clknet_1_0__leaf_net170),
    .B(net172),
    .X(net174));
 sky130_fd_sc_hd__and2_0 c299 (.A(clknet_1_1__leaf_net170),
    .B(clknet_1_1__leaf_net173),
    .X(net175));
 sky130_fd_sc_hd__buf_1 c300 (.A(net601),
    .X(net176));
 sky130_fd_sc_hd__and2_0 c301 (.A(net176),
    .B(net172),
    .X(net177));
 sky130_fd_sc_hd__and3_1 c302 (.A(net171),
    .B(clknet_1_1__leaf_net170),
    .C(clknet_1_0__leaf_net173),
    .X(net178));
 sky130_fd_sc_hd__sdfxtp_1 c303 (.CLK(clknet_leaf_31_clk),
    .D(clknet_1_0__leaf_net175),
    .SCD(net172),
    .SCE(clknet_1_1__leaf_net178),
    .Q(net179));
 sky130_fd_sc_hd__sdfxtp_1 c304 (.CLK(clknet_leaf_31_clk),
    .D(clknet_1_1__leaf_net178),
    .SCD(net176),
    .SCE(net899),
    .Q(net180));
 sky130_fd_sc_hd__mux4_1 c305 (.A0(net63),
    .A1(net177),
    .A2(net180),
    .A3(net176),
    .S0(clknet_1_0__leaf_net174),
    .S1(clknet_1_0__leaf_net170),
    .X(net181));
 sky130_fd_sc_hd__sdfsbp_1 c306 (.CLK(clknet_leaf_31_clk),
    .D(net177),
    .SCD(clknet_1_0__leaf_net178),
    .SCE(clknet_1_0__leaf_net173),
    .SET_B(clknet_1_1__leaf_net170),
    .Q(net183),
    .Q_N(net182));
 sky130_fd_sc_hd__mux4_1 c307 (.A0(net180),
    .A1(clknet_1_0__leaf_net170),
    .A2(net182),
    .A3(clknet_1_0__leaf_net173),
    .S0(net179),
    .S1(net650),
    .X(net184));
 sky130_fd_sc_hd__or4bb_1 c308 (.A(net179),
    .B(net180),
    .C_N(clknet_1_0__leaf_net173),
    .D_N(net172),
    .X(net185));
 sky130_fd_sc_hd__dfbbn_1 c309 (.CLK_N(clknet_leaf_31_clk),
    .D(clknet_1_0__leaf_net174),
    .RESET_B(clknet_1_0__leaf_net185),
    .SET_B(net176),
    .Q(net187),
    .Q_N(net186));
 sky130_fd_sc_hd__sdfsbp_1 c310 (.CLK(clknet_leaf_31_clk),
    .D(clknet_1_1__leaf_net185),
    .SCD(net187),
    .SCE(net899),
    .SET_B(clknet_1_0__leaf_net178),
    .Q(net189),
    .Q_N(net188));
 sky130_fd_sc_hd__and2_0 c311 (.A(net187),
    .B(net189),
    .X(net190));
 sky130_fd_sc_hd__or4bb_1 c312 (.A(net186),
    .B(net916),
    .C_N(net172),
    .D_N(net650),
    .X(net191));
 sky130_fd_sc_hd__mux4_1 c313 (.A0(net189),
    .A1(clknet_1_0__leaf_net184),
    .A2(net190),
    .A3(net191),
    .S0(clknet_1_0__leaf_net173),
    .S1(net172),
    .X(net192));
 sky130_fd_sc_hd__mux4_1 c314 (.A0(net190),
    .A1(net188),
    .A2(net191),
    .A3(clknet_1_1__leaf_net170),
    .S0(clknet_1_1__leaf_net184),
    .S1(net651),
    .X(net193));
 sky130_fd_sc_hd__dlymetal6s2s_1 c315 (.A(net652),
    .X(net194));
 sky130_fd_sc_hd__and2_1 c316 (.A(net100),
    .B(net194),
    .X(net195));
 sky130_fd_sc_hd__and3_1 c317 (.A(net85),
    .B(net195),
    .C(net194),
    .X(net196));
 sky130_fd_sc_hd__and2_1 c318 (.A(net195),
    .B(net755),
    .X(net197));
 sky130_fd_sc_hd__buf_1 c319 (.A(net615),
    .X(net198));
 sky130_fd_sc_hd__dfbbn_1 c320 (.CLK_N(clknet_leaf_32_clk),
    .D(net197),
    .RESET_B(net198),
    .SET_B(net194),
    .Q(net200),
    .Q_N(net199));
 sky130_fd_sc_hd__and2_0 c321 (.A(net194),
    .B(net198),
    .X(net201));
 sky130_fd_sc_hd__and2_1 c322 (.A(net194),
    .B(net201),
    .X(net202));
 sky130_fd_sc_hd__buf_1 c323 (.A(net614),
    .X(net203));
 sky130_fd_sc_hd__and2_1 c324 (.A(net183),
    .B(net198),
    .X(net204));
 sky130_fd_sc_hd__and2_1 c325 (.A(net198),
    .B(net204),
    .X(net205));
 sky130_fd_sc_hd__and3_1 c326 (.A(clknet_1_1__leaf_net173),
    .B(net195),
    .C(net204),
    .X(net206));
 sky130_fd_sc_hd__clkbuf_1 c327 (.A(net629),
    .X(net207));
 sky130_fd_sc_hd__and2_1 c328 (.A(net205),
    .B(net207),
    .X(net208));
 sky130_fd_sc_hd__dfbbp_1 c329 (.CLK(clknet_leaf_32_clk),
    .D(net207),
    .RESET_B(net196),
    .SET_B(net202),
    .Q(net210),
    .Q_N(net209));
 sky130_fd_sc_hd__sdfxbp_1 c330 (.CLK(clknet_leaf_28_clk),
    .D(net204),
    .SCD(clknet_1_0__leaf_net206),
    .SCE(net203),
    .Q(net212),
    .Q_N(net211));
 sky130_fd_sc_hd__sdfxbp_1 c331 (.CLK(clknet_leaf_31_clk),
    .D(net191),
    .SCD(net195),
    .SCE(net208),
    .Q(net214),
    .Q_N(net213));
 sky130_fd_sc_hd__sdfbbp_1 c332 (.CLK(clknet_leaf_31_clk),
    .D(net200),
    .RESET_B(net210),
    .SCD(net208),
    .SCE(net886),
    .SET_B(net887),
    .Q(net216),
    .Q_N(net215));
 sky130_fd_sc_hd__mux4_1 c333 (.A0(net208),
    .A1(net214),
    .A2(net210),
    .A3(net215),
    .S0(net195),
    .S1(net194),
    .X(net217));
 sky130_fd_sc_hd__mux4_1 c334 (.A0(net216),
    .A1(net211),
    .A2(net209),
    .A3(net204),
    .S0(net199),
    .S1(net653),
    .X(net218));
 sky130_fd_sc_hd__mux4_1 c335 (.A0(net201),
    .A1(net212),
    .A2(net218),
    .A3(net209),
    .S0(net205),
    .S1(net653),
    .X(net801));
 sky130_fd_sc_hd__and2_2 c336 (.A(net808),
    .B(net765),
    .X(net219));
 sky130_fd_sc_hd__buf_1 c337 (.A(net219),
    .X(net220));
 sky130_fd_sc_hd__and2_2 c338 (.A(net203),
    .B(net220),
    .X(net221));
 sky130_fd_sc_hd__clkbuf_1 c339 (.X(net613));
 sky130_fd_sc_hd__buf_1 c340 (.A(net834),
    .X(net223));
 sky130_fd_sc_hd__and2_1 c341 (.A(net223),
    .B(net222),
    .X(net224));
 sky130_fd_sc_hd__sdfbbn_1 c342 (.CLK_N(clknet_leaf_25_clk),
    .D(net219),
    .RESET_B(net224),
    .SCD(net220),
    .SCE(net222),
    .SET_B(net221),
    .Q(net226),
    .Q_N(net225));
 sky130_fd_sc_hd__sdfxtp_1 c343 (.CLK(clknet_leaf_27_clk),
    .D(net813),
    .SCD(net219),
    .SCE(net221),
    .Q(net803));
 sky130_fd_sc_hd__a2111o_1 c344 (.A1(net222),
    .A2(net220),
    .B1(net223),
    .C1(net224),
    .D1(net803),
    .X(net227));
 sky130_fd_sc_hd__sdfxtp_1 c345 (.CLK(clknet_leaf_26_clk),
    .D(net224),
    .SCD(net227),
    .SCE(net920),
    .Q(net228));
 sky130_fd_sc_hd__and3_1 c346 (.A(net228),
    .B(net220),
    .C(net224),
    .X(net229));
 sky130_fd_sc_hd__sdfbbn_1 c347 (.CLK_N(clknet_leaf_26_clk),
    .D(net229),
    .RESET_B(net227),
    .SCD(net803),
    .SCE(net220),
    .SET_B(net219),
    .Q(net231),
    .Q_N(net230));
 sky130_fd_sc_hd__and3_2 c348 (.A(net220),
    .B(net231),
    .C(net224),
    .X(net805));
 sky130_fd_sc_hd__sdfstp_1 c349 (.CLK(clknet_leaf_26_clk),
    .D(net221),
    .SCD(net803),
    .SCE(net227),
    .SET_B(net223),
    .Q(net232));
 sky130_fd_sc_hd__mux4_1 c350 (.A0(net232),
    .A1(net229),
    .A2(net223),
    .A3(net222),
    .S0(net805),
    .S1(net219),
    .X(net233));
 sky130_fd_sc_hd__and3_1 c351 (.A(net232),
    .B(net225),
    .C(net810),
    .X(net802));
 sky130_fd_sc_hd__mux4_1 c352 (.A0(net227),
    .A1(net221),
    .A2(net232),
    .A3(net230),
    .S0(net222),
    .S1(net905),
    .X(net234));
 sky130_fd_sc_hd__sdfxtp_1 c353 (.CLK(clknet_leaf_25_clk),
    .D(net224),
    .SCD(net805),
    .SCE(net858),
    .Q(net235));
 sky130_fd_sc_hd__mux4_1 c354 (.A0(net231),
    .A1(net228),
    .A2(net906),
    .A3(net219),
    .S0(net221),
    .S1(net858),
    .X(net236));
 sky130_fd_sc_hd__or4bb_1 c355 (.A(net232),
    .B(net803),
    .C_N(net655),
    .D_N(net658),
    .X(net237));
 sky130_fd_sc_hd__mux4_1 c356 (.A0(net235),
    .A1(net226),
    .A2(net237),
    .A3(net654),
    .S0(net656),
    .S1(net658),
    .X(net804));
 sky130_fd_sc_hd__buf_1 c378 (.A(net144),
    .X(net238));
 sky130_fd_sc_hd__buf_2 c379 (.A(net238),
    .X(net239));
 sky130_fd_sc_hd__clkbuf_1 c380 (.X(net240));
 sky130_fd_sc_hd__clkbuf_1 c381 (.A(net616),
    .X(net241));
 sky130_fd_sc_hd__dfrtp_1 c382 (.CLK(clknet_leaf_10_clk),
    .D(net240),
    .RESET_B(net239),
    .Q(net242));
 sky130_fd_sc_hd__dfrtp_1 c383 (.CLK(clknet_leaf_10_clk),
    .D(net833),
    .RESET_B(net239),
    .Q(net243));
 sky130_fd_sc_hd__and3_1 c384 (.A(net243),
    .B(net242),
    .C(net241),
    .X(net244));
 sky130_fd_sc_hd__dfrtp_1 c385 (.CLK(clknet_leaf_5_clk),
    .D(net239),
    .RESET_B(net238),
    .Q(net245));
 sky130_fd_sc_hd__sdfbbp_1 c386 (.CLK(clknet_leaf_7_clk),
    .D(net238),
    .RESET_B(net863),
    .SCD(net241),
    .SCE(net244),
    .SET_B(net239),
    .Q(net247),
    .Q_N(net246));
 sky130_fd_sc_hd__sdfstp_1 c387 (.CLK(clknet_leaf_10_clk),
    .D(net140),
    .SCD(net889),
    .SCE(net244),
    .SET_B(net239),
    .Q(net248));
 sky130_fd_sc_hd__and3_1 c388 (.A(net241),
    .B(net240),
    .C(net246),
    .X(net249));
 sky130_fd_sc_hd__and2_1 c389 (.A(net248),
    .B(net247),
    .X(net250));
 sky130_fd_sc_hd__and2_0 c390 (.A(net250),
    .B(net245),
    .X(net251));
 sky130_fd_sc_hd__sdfstp_1 c391 (.CLK(clknet_leaf_4_clk),
    .D(net244),
    .SCD(net251),
    .SCE(net250),
    .SET_B(net239),
    .Q(net252));
 sky130_fd_sc_hd__mux4_1 c392 (.A0(net251),
    .A1(net250),
    .A2(net239),
    .A3(net249),
    .S0(net252),
    .S1(net863),
    .X(net253));
 sky130_fd_sc_hd__or4bb_1 c393 (.A(net889),
    .B(net249),
    .C_N(net238),
    .D_N(net917),
    .X(net254));
 sky130_fd_sc_hd__and2_0 c394 (.A(net245),
    .B(net249),
    .X(net255));
 sky130_fd_sc_hd__sedfxbp_1 c395 (.CLK(clknet_leaf_12_clk),
    .D(net255),
    .DE(net250),
    .SCD(net254),
    .SCE(net912),
    .Q(net257),
    .Q_N(net256));
 sky130_fd_sc_hd__or4bb_1 c396 (.A(net255),
    .B(net251),
    .C_N(net244),
    .D_N(net648),
    .X(net258));
 sky130_fd_sc_hd__sedfxbp_1 c397 (.CLK(clknet_leaf_12_clk),
    .D(net247),
    .DE(net258),
    .SCD(net250),
    .SCE(net256),
    .Q(net259));
 sky130_fd_sc_hd__sedfxtp_1 c398 (.CLK(clknet_leaf_12_clk),
    .D(net249),
    .DE(net257),
    .SCD(net857),
    .SCE(net258),
    .Q(net260));
 sky130_fd_sc_hd__buf_1 c399 (.A(net921),
    .X(net261));
 sky130_fd_sc_hd__clkbuf_2 c400 (.A(net261),
    .X(net262));
 sky130_fd_sc_hd__and2_1 c401 (.A(net261),
    .B(net262),
    .X(net263));
 sky130_fd_sc_hd__clkbuf_1 c402 (.X(net264));
 sky130_fd_sc_hd__and2_1 c403 (.A(net895),
    .B(net262),
    .X(net265));
 sky130_fd_sc_hd__buf_1 c404 (.A(net612),
    .X(net266));
 sky130_fd_sc_hd__dfbbn_1 c405 (.CLK_N(clknet_leaf_2_clk),
    .D(net252),
    .RESET_B(net265),
    .SET_B(net266),
    .Q(net268),
    .Q_N(net267));
 sky130_fd_sc_hd__dfbbn_1 c406 (.CLK_N(clknet_leaf_2_clk),
    .D(net263),
    .RESET_B(net266),
    .SET_B(net842),
    .Q(net270),
    .Q_N(net269));
 sky130_fd_sc_hd__and3_1 c407 (.A(net261),
    .B(net267),
    .C(net262),
    .X(net271));
 sky130_fd_sc_hd__dfsbp_1 c408 (.CLK(clknet_leaf_2_clk),
    .D(net265),
    .SET_B(net269),
    .Q(net273),
    .Q_N(net272));
 sky130_fd_sc_hd__dfbbp_1 c409 (.CLK(clknet_leaf_2_clk),
    .D(net907),
    .RESET_B(net270),
    .SET_B(net271),
    .Q(net275),
    .Q_N(net274));
 sky130_fd_sc_hd__or4bb_1 c410 (.A(net270),
    .B(net268),
    .C_N(net272),
    .D_N(net262),
    .X(net276));
 sky130_fd_sc_hd__and3_1 c411 (.A(net262),
    .B(net275),
    .C(net272),
    .X(net277));
 sky130_fd_sc_hd__sdfxbp_1 c412 (.CLK(clknet_leaf_2_clk),
    .D(net266),
    .SCD(net276),
    .SCE(net274),
    .Q(net279),
    .Q_N(net278));
 sky130_fd_sc_hd__sdfxbp_1 c413 (.CLK(clknet_leaf_3_clk),
    .D(net846),
    .SCD(net277),
    .SCE(net276),
    .Q(net281),
    .Q_N(net280));
 sky130_fd_sc_hd__and3_1 c414 (.A(net275),
    .B(net273),
    .C(net280),
    .X(net282));
 sky130_fd_sc_hd__sdfxtp_1 c415 (.CLK(clknet_leaf_30_clk),
    .D(net839),
    .SCD(net282),
    .SCE(net263),
    .Q(net283));
 sky130_fd_sc_hd__mux4_1 c416 (.A0(net265),
    .A1(net283),
    .A2(net262),
    .A3(net272),
    .S0(net895),
    .S1(net263),
    .X(net284));
 sky130_fd_sc_hd__and3_1 c417 (.A(net268),
    .B(net278),
    .C(net660),
    .X(net285));
 sky130_fd_sc_hd__mux4_1 c418 (.A0(net263),
    .A1(net282),
    .A2(net285),
    .A3(net283),
    .S0(net262),
    .S1(net261),
    .X(net286));
 sky130_fd_sc_hd__and3_1 c419 (.A(net282),
    .B(net660),
    .C(net661),
    .X(net287));
 sky130_fd_sc_hd__buf_1 c420 (.A(net287),
    .X(net288));
 sky130_fd_sc_hd__buf_1 c421 (.X(net289));
 sky130_fd_sc_hd__buf_1 c422 (.A(net610),
    .X(net290));
 sky130_fd_sc_hd__dfsbp_1 c423 (.CLK(clknet_leaf_30_clk),
    .D(clknet_1_0__leaf_net289),
    .SET_B(clknet_1_0__leaf_net288),
    .Q(net292),
    .Q_N(net291));
 sky130_fd_sc_hd__and2_1 c424 (.A(net292),
    .B(net290),
    .X(net293));
 sky130_fd_sc_hd__buf_1 c425 (.A(net633),
    .X(net294));
 sky130_fd_sc_hd__and2_1 c426 (.A(net293),
    .B(net290),
    .X(net295));
 sky130_fd_sc_hd__and3_1 c427 (.A(net293),
    .B(net292),
    .C(net295),
    .X(net296));
 sky130_fd_sc_hd__dfstp_1 c428 (.CLK(clknet_leaf_30_clk),
    .D(net296),
    .SET_B(net295),
    .Q(net297));
 sky130_fd_sc_hd__sdfxtp_1 c429 (.CLK(clknet_leaf_30_clk),
    .D(net907),
    .SCD(net865),
    .SCE(clknet_1_0__leaf_net288),
    .Q(net298));
 sky130_fd_sc_hd__sdfxtp_1 c430 (.CLK(clknet_leaf_30_clk),
    .D(net296),
    .SCD(net293),
    .SCE(net892),
    .Q(net299));
 sky130_fd_sc_hd__and2_1 c431 (.A(net295),
    .B(net290),
    .X(net300));
 sky130_fd_sc_hd__dfstp_1 c432 (.CLK(clknet_leaf_30_clk),
    .D(net838),
    .SET_B(net300),
    .Q(net301));
 sky130_fd_sc_hd__sedfxtp_1 c433 (.CLK(clknet_leaf_30_clk),
    .D(net271),
    .DE(net298),
    .SCD(net300),
    .SCE(net297),
    .Q(net302));
 sky130_fd_sc_hd__mux4_1 c434 (.A0(net300),
    .A1(net299),
    .A2(net298),
    .A3(net297),
    .S0(clknet_1_1__leaf_net288),
    .S1(net293),
    .X(net303));
 sky130_fd_sc_hd__dfbbn_1 c435 (.CLK_N(clknet_leaf_30_clk),
    .D(net290),
    .RESET_B(net300),
    .SET_B(net868),
    .Q(net305),
    .Q_N(net304));
 sky130_fd_sc_hd__and3_1 c436 (.A(net892),
    .B(net302),
    .C(net294),
    .X(net306));
 sky130_fd_sc_hd__and3_1 c437 (.A(net301),
    .B(net306),
    .C(net304),
    .X(net307));
 sky130_fd_sc_hd__and2_0 c438 (.A(clknet_1_0__leaf_net289),
    .B(net297),
    .X(net308));
 sky130_fd_sc_hd__or4bb_1 c439 (.A(net305),
    .B(net307),
    .C_N(net308),
    .D_N(clknet_1_0__leaf_net662),
    .X(net309));
 sky130_fd_sc_hd__dfbbn_1 c440 (.CLK_N(clknet_leaf_29_clk),
    .D(net302),
    .RESET_B(net306),
    .SET_B(clknet_1_0__leaf_net309),
    .Q(net310));
 sky130_fd_sc_hd__buf_1 c441 (.A(net600),
    .X(net311));
 sky130_fd_sc_hd__and2_1 c442 (.A(net310),
    .B(net311),
    .X(net312));
 sky130_fd_sc_hd__and2_2 c443 (.A(net294),
    .B(net312),
    .X(net313));
 sky130_fd_sc_hd__and2_1 c444 (.A(net311),
    .B(net313),
    .X(net314));
 sky130_fd_sc_hd__and2_0 c445 (.A(net311),
    .B(net313),
    .X(net315));
 sky130_fd_sc_hd__buf_1 c446 (.A(net891),
    .X(net316));
 sky130_fd_sc_hd__and3_2 c447 (.A(net313),
    .B(net316),
    .C(net312),
    .X(net317));
 sky130_fd_sc_hd__dfbbp_1 c448 (.CLK(clknet_leaf_26_clk),
    .D(clknet_1_1__leaf_net206),
    .RESET_B(net317),
    .SET_B(net313),
    .Q(net319),
    .Q_N(net318));
 sky130_fd_sc_hd__buf_1 c449 (.A(net630),
    .X(net320));
 sky130_fd_sc_hd__sdfbbn_1 c450 (.CLK_N(clknet_leaf_29_clk),
    .D(net314),
    .RESET_B(net316),
    .SCD(net312),
    .SCE(net313),
    .SET_B(net317),
    .Q(net322),
    .Q_N(net321));
 sky130_fd_sc_hd__and2_1 c451 (.A(net297),
    .B(net320),
    .X(net323));
 sky130_fd_sc_hd__clkbuf_1 c452 (.A(net633),
    .X(net324));
 sky130_fd_sc_hd__mux4_1 c453 (.A0(net316),
    .A1(net317),
    .A2(net324),
    .A3(net323),
    .S0(net321),
    .S1(net313),
    .X(net325));
 sky130_fd_sc_hd__sedfxtp_1 c454 (.CLK(clknet_leaf_29_clk),
    .D(net323),
    .DE(net317),
    .SCD(net313),
    .SCE(clknet_1_0__leaf_net663),
    .Q(net326));
 sky130_fd_sc_hd__mux4_1 c455 (.A0(net210),
    .A1(net326),
    .A2(net320),
    .A3(net323),
    .S0(net313),
    .S1(clknet_1_0__leaf_net663),
    .X(net327));
 sky130_fd_sc_hd__mux4_1 c456 (.A0(net324),
    .A1(clknet_1_0__leaf_net327),
    .A2(net322),
    .A3(net318),
    .S0(net313),
    .S1(net317),
    .X(net328));
 sky130_fd_sc_hd__mux4_1 c457 (.A0(net326),
    .A1(net314),
    .A2(net315),
    .A3(net317),
    .S0(clknet_1_0__leaf_net327),
    .S1(clknet_1_1__leaf_net663),
    .X(net329));
 sky130_fd_sc_hd__mux4_1 c458 (.A0(net319),
    .A1(net316),
    .A2(clknet_1_1__leaf_net327),
    .A3(clknet_1_1__leaf_net663),
    .S0(net664),
    .S1(net667),
    .X(net330));
 sky130_fd_sc_hd__mux4_1 c459 (.A0(net214),
    .A1(net322),
    .A2(net323),
    .A3(net317),
    .S0(net666),
    .S1(net668),
    .X(net331));
 sky130_fd_sc_hd__mux4_1 c460 (.A0(net317),
    .A1(net311),
    .A2(net665),
    .A3(net666),
    .S0(net799),
    .S1(net792),
    .X(net332));
 sky130_fd_sc_hd__mux4_1 c461 (.A0(net320),
    .A1(net321),
    .A2(net667),
    .A3(net799),
    .S0(net792),
    .S1(net669),
    .X(net797));
 sky130_fd_sc_hd__buf_1 c462 (.A(net668),
    .X(net333));
 sky130_fd_sc_hd__clkbuf_1 c463 (.A(net333),
    .X(net334));
 sky130_fd_sc_hd__and2_1 c464 (.A(net334),
    .B(net333),
    .X(net335));
 sky130_fd_sc_hd__buf_1 c465 (.X(net800));
 sky130_fd_sc_hd__clkbuf_1 c466 (.A(net608),
    .X(net336));
 sky130_fd_sc_hd__and2_0 c467 (.A(net334),
    .B(net336),
    .X(net337));
 sky130_fd_sc_hd__clkbuf_1 c468 (.A(net853),
    .X(net338));
 sky130_fd_sc_hd__and2_1 c469 (.A(net336),
    .B(net338),
    .X(net339));
 sky130_fd_sc_hd__and2_1 c470 (.A(net338),
    .B(net339),
    .X(net340));
 sky130_fd_sc_hd__dfstp_1 c471 (.CLK(clknet_leaf_23_clk),
    .D(net337),
    .SET_B(net340),
    .Q(net794));
 sky130_fd_sc_hd__sdfxbp_1 c472 (.CLK(clknet_leaf_23_clk),
    .D(net339),
    .SCD(net335),
    .SCE(net794),
    .Q(net342),
    .Q_N(net341));
 sky130_fd_sc_hd__sdfxbp_1 c473 (.CLK(clknet_leaf_23_clk),
    .D(net335),
    .SCD(net883),
    .SCE(net339),
    .Q(net344),
    .Q_N(net343));
 sky130_fd_sc_hd__and3_1 c474 (.A(net344),
    .B(net340),
    .C(net339),
    .X(net345));
 sky130_fd_sc_hd__sdfxtp_1 c475 (.CLK(clknet_leaf_22_clk),
    .D(net844),
    .SCD(net345),
    .SCE(net794),
    .Q(net346));
 sky130_fd_sc_hd__sdfxtp_1 c476 (.CLK(clknet_leaf_23_clk),
    .D(net333),
    .SCD(net881),
    .SCE(net345),
    .Q(net347));
 sky130_fd_sc_hd__and3_1 c477 (.A(net347),
    .B(net339),
    .C(net346),
    .X(net348));
 sky130_fd_sc_hd__and3_1 c478 (.A(net348),
    .B(net346),
    .C(net340),
    .X(net798));
 sky130_fd_sc_hd__sdfxtp_1 c479 (.CLK(clknet_leaf_22_clk),
    .D(net798),
    .SCD(net345),
    .SCE(net852),
    .Q(net349));
 sky130_fd_sc_hd__dfbbn_1 c480 (.CLK_N(clknet_leaf_22_clk),
    .D(net346),
    .RESET_B(net348),
    .SET_B(net345),
    .Q(net351),
    .Q_N(net350));
 sky130_fd_sc_hd__dfbbn_1 c481 (.CLK_N(clknet_leaf_22_clk),
    .D(clknet_1_1__leaf_net309),
    .RESET_B(net349),
    .SET_B(net871),
    .Q(net791),
    .Q_N(net795));
 sky130_fd_sc_hd__or4bb_1 c482 (.A(net349),
    .B(net351),
    .C_N(net348),
    .D_N(net795),
    .X(net793));
 sky130_fd_sc_hd__buf_1 c504 (.A(net260),
    .X(net352));
 sky130_fd_sc_hd__clkbuf_2 c505 (.A(net352),
    .X(net353));
 sky130_fd_sc_hd__and2_2 c506 (.A(net353),
    .B(net352),
    .X(net354));
 sky130_fd_sc_hd__buf_1 c507 (.A(net621),
    .X(net355));
 sky130_fd_sc_hd__dlymetal6s2s_1 c508 (.A(net620),
    .X(net356));
 sky130_fd_sc_hd__dfbbp_1 c509 (.CLK(clknet_leaf_10_clk),
    .D(net353),
    .RESET_B(net356),
    .SET_B(net354),
    .Q(net358),
    .Q_N(net357));
 sky130_fd_sc_hd__and3_1 c510 (.A(net355),
    .B(net356),
    .C(net353),
    .X(net359));
 sky130_fd_sc_hd__and3_1 c511 (.A(net355),
    .B(net357),
    .C(net356),
    .X(net360));
 sky130_fd_sc_hd__sdfxbp_1 c512 (.CLK(clknet_leaf_11_clk),
    .D(net254),
    .SCD(net359),
    .SCE(net356),
    .Q(net362),
    .Q_N(net361));
 sky130_fd_sc_hd__sdfxbp_1 c513 (.CLK(clknet_leaf_10_clk),
    .D(net884),
    .SCD(net356),
    .SCE(net354),
    .Q(net364),
    .Q_N(net363));
 sky130_fd_sc_hd__and3_1 c514 (.A(net358),
    .B(net364),
    .C(net353),
    .X(net365));
 sky130_fd_sc_hd__sdfxtp_1 c515 (.CLK(clknet_leaf_11_clk),
    .D(net354),
    .SCD(net884),
    .SCE(net365),
    .Q(net366));
 sky130_fd_sc_hd__sdfxtp_1 c516 (.CLK(clknet_leaf_11_clk),
    .D(net365),
    .SCD(net870),
    .SCE(net913),
    .Q(net367));
 sky130_fd_sc_hd__and3_1 c517 (.A(net360),
    .B(net367),
    .C(net362),
    .X(net368));
 sky130_fd_sc_hd__sdfbbn_1 c518 (.CLK_N(clknet_leaf_10_clk),
    .D(net368),
    .RESET_B(net363),
    .SCD(net356),
    .SCE(net354),
    .SET_B(net353),
    .Q(net370),
    .Q_N(net369));
 sky130_fd_sc_hd__mux4_1 c519 (.A0(net356),
    .A1(net366),
    .A2(net368),
    .A3(net361),
    .S0(net355),
    .S1(net353),
    .X(net371));
 sky130_fd_sc_hd__and3_1 c520 (.A(net370),
    .B(net352),
    .C(net360),
    .X(net372));
 sky130_fd_sc_hd__sdfxtp_1 c521 (.CLK(clknet_leaf_11_clk),
    .D(net359),
    .SCD(net368),
    .SCE(net371),
    .Q(net373));
 sky130_fd_sc_hd__a2111o_1 c522 (.A1(net373),
    .A2(net364),
    .B1(net353),
    .C1(net372),
    .D1(net362),
    .X(net374));
 sky130_fd_sc_hd__mux4_1 c523 (.A0(net372),
    .A1(net374),
    .A2(net371),
    .A3(net373),
    .S0(net354),
    .S1(net353),
    .X(net375));
 sky130_fd_sc_hd__mux4_1 c524 (.A0(net366),
    .A1(net371),
    .A2(net374),
    .A3(net372),
    .S0(net369),
    .S1(net361),
    .X(net376));
 sky130_fd_sc_hd__dlymetal6s2s_1 c525 (.A(net670),
    .X(net377));
 sky130_fd_sc_hd__buf_1 c526 (.A(net377),
    .X(net378));
 sky130_fd_sc_hd__and2_1 c527 (.A(net377),
    .B(net378),
    .X(net379));
 sky130_fd_sc_hd__and2_2 c528 (.A(net378),
    .B(net377),
    .X(net380));
 sky130_fd_sc_hd__clkbuf_1 c529 (.A(net596),
    .X(net381));
 sky130_fd_sc_hd__clkbuf_1 c530 (.A(net595),
    .X(net382));
 sky130_fd_sc_hd__dfbbn_1 c531 (.CLK_N(clknet_leaf_4_clk),
    .D(net382),
    .RESET_B(net377),
    .SET_B(net379),
    .Q(net384),
    .Q_N(net383));
 sky130_fd_sc_hd__dlrbn_1 c532 (.D(net377),
    .GATE_N(clknet_leaf_12_clk),
    .RESET_B(net380),
    .Q(net386),
    .Q_N(net385));
 sky130_fd_sc_hd__dfbbn_1 c533 (.CLK_N(clknet_leaf_4_clk),
    .D(net877),
    .RESET_B(net382),
    .SET_B(net380),
    .Q(net388),
    .Q_N(net387));
 sky130_fd_sc_hd__dlrbn_1 c534 (.D(net388),
    .GATE_N(clknet_leaf_4_clk),
    .RESET_B(net379),
    .Q(net390),
    .Q_N(net389));
 sky130_fd_sc_hd__and3_1 c535 (.A(net390),
    .B(net386),
    .C(net377),
    .X(net391));
 sky130_fd_sc_hd__dlrbp_1 c536 (.D(net386),
    .GATE(clknet_leaf_12_clk),
    .RESET_B(net380),
    .Q(net393),
    .Q_N(net392));
 sky130_fd_sc_hd__and3_1 c537 (.A(net854),
    .B(net391),
    .C(net385),
    .X(net394));
 sky130_fd_sc_hd__dlrbp_1 c538 (.D(net394),
    .GATE(clknet_leaf_13_clk),
    .RESET_B(net877),
    .Q(net396),
    .Q_N(net395));
 sky130_fd_sc_hd__and3_1 c539 (.A(net381),
    .B(net392),
    .C(net395),
    .X(net397));
 sky130_fd_sc_hd__and3_1 c540 (.A(net397),
    .B(net384),
    .C(net389),
    .X(net398));
 sky130_fd_sc_hd__sdfbbp_1 c541 (.CLK(clknet_leaf_4_clk),
    .D(net854),
    .RESET_B(net398),
    .SCD(net890),
    .SCE(net380),
    .SET_B(net383),
    .Q(net400),
    .Q_N(net399));
 sky130_fd_sc_hd__dfbbp_1 c542 (.CLK(clknet_leaf_3_clk),
    .D(net391),
    .RESET_B(net394),
    .SET_B(net837),
    .Q(net402),
    .Q_N(net401));
 sky130_fd_sc_hd__and3_1 c543 (.A(net400),
    .B(net387),
    .C(net381),
    .X(net403));
 sky130_fd_sc_hd__mux4_1 c544 (.A0(net277),
    .A1(net402),
    .A2(net397),
    .A3(net403),
    .S0(net398),
    .S1(net379),
    .X(net404));
 sky130_fd_sc_hd__sdfbbn_1 c545 (.CLK_N(clknet_leaf_3_clk),
    .D(net403),
    .RESET_B(net401),
    .SCD(net380),
    .SCE(net383),
    .SET_B(net672),
    .Q(net406),
    .Q_N(net405));
 sky130_fd_sc_hd__clkbuf_2 c546 (.A(net405),
    .X(net407));
 sky130_fd_sc_hd__clkbuf_2 c547 (.A(net628),
    .X(net408));
 sky130_fd_sc_hd__and2_1 c548 (.A(net408),
    .B(net407),
    .X(net409));
 sky130_fd_sc_hd__and2_0 c549 (.A(net408),
    .B(net407),
    .X(net410));
 sky130_fd_sc_hd__and2_2 c550 (.A(net409),
    .B(net407),
    .X(net411));
 sky130_fd_sc_hd__and2_1 c551 (.A(net408),
    .B(net409),
    .X(net412));
 sky130_fd_sc_hd__sdfxbp_1 c552 (.CLK(clknet_leaf_13_clk),
    .D(net412),
    .SCD(net410),
    .SCE(net411),
    .Q(net414),
    .Q_N(net413));
 sky130_fd_sc_hd__sdfxbp_1 c553 (.CLK(clknet_leaf_3_clk),
    .D(net407),
    .SCD(net408),
    .SCE(net411),
    .Q(net416),
    .Q_N(net415));
 sky130_fd_sc_hd__clkbuf_1 c554 (.A(net628),
    .X(net417));
 sky130_fd_sc_hd__sdfxtp_1 c555 (.CLK(clknet_leaf_30_clk),
    .D(net409),
    .SCD(net411),
    .SCE(net412),
    .Q(net418));
 sky130_fd_sc_hd__and2_0 c556 (.A(net418),
    .B(clknet_1_1__leaf_net662),
    .X(net419));
 sky130_fd_sc_hd__dlrtn_1 c557 (.D(net411),
    .GATE_N(clknet_leaf_3_clk),
    .RESET_B(net829),
    .Q(net420));
 sky130_fd_sc_hd__and3_1 c558 (.A(net418),
    .B(clknet_1_0__leaf_net419),
    .C(net417),
    .X(net421));
 sky130_fd_sc_hd__and3_1 c559 (.A(net420),
    .B(net407),
    .C(net850),
    .X(net422));
 sky130_fd_sc_hd__and3_1 c560 (.A(net407),
    .B(clknet_1_0__leaf_net421),
    .C(net420),
    .X(net423));
 sky130_fd_sc_hd__sdfbbn_1 c561 (.CLK_N(clknet_leaf_18_clk),
    .D(clknet_1_0__leaf_net423),
    .RESET_B(net411),
    .SCD(clknet_1_0__leaf_net419),
    .SCE(clknet_1_0__leaf_net421),
    .SET_B(net407),
    .Q(net425),
    .Q_N(net424));
 sky130_fd_sc_hd__and3_1 c562 (.A(net410),
    .B(net422),
    .C(net409),
    .X(net426));
 sky130_fd_sc_hd__mux4_1 c563 (.A0(net425),
    .A1(net420),
    .A2(clknet_1_1__leaf_net421),
    .A3(net426),
    .S0(clknet_1_1__leaf_net423),
    .S1(net408),
    .X(net427));
 sky130_fd_sc_hd__mux4_1 c564 (.A0(net285),
    .A1(net417),
    .A2(clknet_1_0__leaf_net421),
    .A3(net424),
    .S0(net408),
    .S1(net420),
    .X(net428));
 sky130_fd_sc_hd__mux4_1 c565 (.A0(net426),
    .A1(net428),
    .A2(net424),
    .A3(net411),
    .S0(clknet_1_1__leaf_net421),
    .S1(net673),
    .X(net429));
 sky130_fd_sc_hd__sdfrbp_1 c566 (.CLK(clknet_leaf_19_clk),
    .D(net425),
    .RESET_B(net426),
    .SCD(net888),
    .SCE(net896),
    .Q(net430));
 sky130_fd_sc_hd__buf_1 c567 (.A(net430),
    .X(net431));
 sky130_fd_sc_hd__buf_1 c568 (.A(net431),
    .X(net432));
 sky130_fd_sc_hd__and2_0 c569 (.A(clknet_1_1__leaf_net419),
    .B(net432),
    .X(net433));
 sky130_fd_sc_hd__and2_1 c570 (.A(net432),
    .B(net431),
    .X(net434));
 sky130_fd_sc_hd__buf_1 c571 (.A(net626),
    .X(net435));
 sky130_fd_sc_hd__buf_1 c572 (.A(net625),
    .X(net436));
 sky130_fd_sc_hd__dlrtn_1 c573 (.D(net436),
    .GATE_N(clknet_leaf_19_clk),
    .RESET_B(clknet_1_0__leaf_net433),
    .Q(net437));
 sky130_fd_sc_hd__sdfxtp_1 c574 (.CLK(clknet_leaf_19_clk),
    .D(net437),
    .SCD(net434),
    .SCE(net435),
    .Q(net438));
 sky130_fd_sc_hd__and3_1 c575 (.A(net438),
    .B(net437),
    .C(net436),
    .X(net439));
 sky130_fd_sc_hd__and2_0 c576 (.A(net438),
    .B(net439),
    .X(net440));
 sky130_fd_sc_hd__sdfxtp_1 c577 (.CLK(clknet_leaf_19_clk),
    .D(net434),
    .SCD(net440),
    .SCE(net436),
    .Q(net441));
 sky130_fd_sc_hd__dfbbn_1 c578 (.CLK_N(clknet_leaf_29_clk),
    .D(net314),
    .RESET_B(net441),
    .SET_B(net867),
    .Q(net442));
 sky130_fd_sc_hd__and3_1 c579 (.A(net432),
    .B(net435),
    .C(net431),
    .X(net443));
 sky130_fd_sc_hd__and2_0 c580 (.A(net435),
    .B(net437),
    .X(net444));
 sky130_fd_sc_hd__and2_1 c581 (.A(net431),
    .B(net439),
    .X(net445));
 sky130_fd_sc_hd__and3_1 c582 (.A(net444),
    .B(net445),
    .C(net439),
    .X(net446));
 sky130_fd_sc_hd__a2111o_1 c583 (.A1(net441),
    .A2(net898),
    .B1(net435),
    .C1(net445),
    .D1(net436),
    .X(net447));
 sky130_fd_sc_hd__dfbbn_1 c584 (.CLK_N(clknet_leaf_19_clk),
    .D(net439),
    .RESET_B(net447),
    .SET_B(net445),
    .Q(net449),
    .Q_N(net448));
 sky130_fd_sc_hd__sdfbbp_1 c585 (.CLK(clknet_leaf_19_clk),
    .D(net440),
    .RESET_B(net446),
    .SCD(net449),
    .SCE(net445),
    .SET_B(net437),
    .Q(net451),
    .Q_N(net450));
 sky130_fd_sc_hd__mux4_1 c586 (.A0(net449),
    .A1(net451),
    .A2(net444),
    .A3(net432),
    .S0(net443),
    .S1(clknet_1_1__leaf_net433),
    .X(net452));
 sky130_fd_sc_hd__mux4_1 c587 (.A0(net450),
    .A1(net448),
    .A2(net446),
    .A3(net441),
    .S0(net668),
    .S1(net878),
    .X(net453));
 sky130_fd_sc_hd__buf_1 c588 (.A(clknet_1_1__leaf_net419),
    .X(net454));
 sky130_fd_sc_hd__buf_1 c589 (.A(clknet_1_1__leaf_net454),
    .X(net455));
 sky130_fd_sc_hd__clkbuf_1 c590 (.A(net901),
    .X(net456));
 sky130_fd_sc_hd__dfbbp_1 c591 (.CLK(clknet_leaf_21_clk),
    .D(net456),
    .RESET_B(clknet_1_1__leaf_net455),
    .SET_B(clknet_1_1__leaf_net454),
    .Q(net458),
    .Q_N(net457));
 sky130_fd_sc_hd__buf_1 c592 (.A(net605),
    .X(net459));
 sky130_fd_sc_hd__and2_2 c593 (.A(net459),
    .B(net458),
    .X(net460));
 sky130_fd_sc_hd__sdfxbp_1 c594 (.CLK(clknet_leaf_23_clk),
    .D(clknet_1_0__leaf_net455),
    .SCD(clknet_1_0__leaf_net454),
    .SCE(net459),
    .Q(net462),
    .Q_N(net461));
 sky130_fd_sc_hd__and3_1 c595 (.A(net460),
    .B(net459),
    .C(net835),
    .X(net463));
 sky130_fd_sc_hd__clkbuf_1 c596 (.A(net634),
    .X(net464));
 sky130_fd_sc_hd__sdfxbp_1 c597 (.CLK(clknet_leaf_20_clk),
    .D(net460),
    .SCD(clknet_1_1__leaf_net455),
    .SCE(net872),
    .Q(net466),
    .Q_N(net465));
 sky130_fd_sc_hd__and2_2 c598 (.A(net466),
    .B(net460),
    .X(net790));
 sky130_fd_sc_hd__mux4_1 c599 (.A0(net464),
    .A1(net465),
    .A2(net459),
    .A3(net460),
    .S0(net458),
    .S1(net790),
    .X(net467));
 sky130_fd_sc_hd__or4bb_1 c600 (.A(net823),
    .B(net463),
    .C_N(net459),
    .D_N(net790),
    .X(net468));
 sky130_fd_sc_hd__sdfxtp_1 c601 (.CLK(clknet_leaf_21_clk),
    .D(net468),
    .SCD(net460),
    .SCE(net790),
    .Q(net469));
 sky130_fd_sc_hd__sdfrbp_1 c602 (.CLK(clknet_leaf_21_clk),
    .D(net848),
    .RESET_B(net836),
    .SCD(net460),
    .SCE(net790),
    .Q(net471),
    .Q_N(net470));
 sky130_fd_sc_hd__sdfxtp_1 c603 (.CLK(clknet_leaf_22_clk),
    .D(net840),
    .SCD(net790),
    .SCE(net467),
    .Q(net472));
 sky130_fd_sc_hd__mux4_1 c604 (.A0(net462),
    .A1(net463),
    .A2(net472),
    .A3(clknet_1_0__leaf_net454),
    .S0(clknet_1_0__leaf_net455),
    .S1(net460),
    .X(net473));
 sky130_fd_sc_hd__mux4_1 c605 (.A0(net472),
    .A1(net467),
    .A2(net459),
    .A3(clknet_1_0__leaf_net455),
    .S0(clknet_1_0__leaf_net454),
    .S1(net464),
    .X(net474));
 sky130_fd_sc_hd__sdfbbn_1 c606 (.CLK_N(clknet_leaf_21_clk),
    .D(clknet_1_1__leaf_net454),
    .RESET_B(net468),
    .SCD(net790),
    .SCE(net460),
    .SET_B(net678),
    .Q(net476),
    .Q_N(net475));
 sky130_fd_sc_hd__mux4_1 c607 (.A0(net476),
    .A1(net472),
    .A2(net469),
    .A3(net790),
    .S0(net678),
    .S1(clknet_1_0__leaf_net679),
    .X(net477));
 sky130_fd_sc_hd__mux4_1 c608 (.A0(net477),
    .A1(net475),
    .A2(net456),
    .A3(net470),
    .S0(net678),
    .S1(clknet_1_1__leaf_net679),
    .X(net478));
 sky130_fd_sc_hd__clkbuf_2 c630 (.A(net670),
    .X(net479));
 sky130_fd_sc_hd__buf_1 c631 (.A(net479),
    .X(net480));
 sky130_fd_sc_hd__and2_0 c632 (.A(net367),
    .B(net479),
    .X(net481));
 sky130_fd_sc_hd__and2_1 c633 (.A(net480),
    .B(net479),
    .X(net482));
 sky130_fd_sc_hd__and2_0 c634 (.A(net480),
    .B(net479),
    .X(net483));
 sky130_fd_sc_hd__buf_1 c635 (.X(net484));
 sky130_fd_sc_hd__and2_0 c636 (.A(net484),
    .B(net671),
    .X(net485));
 sky130_fd_sc_hd__clkbuf_1 c637 (.A(net607),
    .X(net486));
 sky130_fd_sc_hd__dlrtn_1 c638 (.D(net485),
    .GATE_N(clknet_leaf_11_clk),
    .RESET_B(net482),
    .Q(net487));
 sky130_fd_sc_hd__and2_0 c639 (.A(net487),
    .B(net486),
    .X(net488));
 sky130_fd_sc_hd__sdfxtp_1 c640 (.CLK(clknet_leaf_14_clk),
    .D(net479),
    .SCD(net482),
    .SCE(net483),
    .Q(net489));
 sky130_fd_sc_hd__and2_1 c641 (.A(net489),
    .B(net487),
    .X(net490));
 sky130_fd_sc_hd__or4bb_1 c642 (.A(net488),
    .B(net490),
    .C_N(net489),
    .D_N(net481),
    .X(net491));
 sky130_fd_sc_hd__and3_1 c643 (.A(net486),
    .B(net490),
    .C(net484),
    .X(net492));
 sky130_fd_sc_hd__a2111o_1 c644 (.A1(net484),
    .A2(net492),
    .B1(net487),
    .C1(net490),
    .D1(net479),
    .X(net493));
 sky130_fd_sc_hd__sdfrtn_1 c645 (.CLK_N(clknet_leaf_11_clk),
    .D(net493),
    .RESET_B(net828),
    .SCD(net490),
    .SCE(net489),
    .Q(net494));
 sky130_fd_sc_hd__mux4_1 c646 (.A0(net491),
    .A1(net487),
    .A2(net493),
    .A3(net479),
    .S0(net494),
    .S1(net480),
    .X(net495));
 sky130_fd_sc_hd__dfbbn_1 c647 (.CLK_N(clknet_leaf_15_clk),
    .D(net491),
    .RESET_B(net489),
    .SET_B(clknet_1_0__leaf_net680),
    .Q(net497),
    .Q_N(net496));
 sky130_fd_sc_hd__mux4_1 c648 (.A0(net485),
    .A1(net494),
    .A2(net489),
    .A3(net482),
    .S0(net496),
    .S1(net479),
    .X(net498));
 sky130_fd_sc_hd__mux4_1 c649 (.A0(net481),
    .A1(net494),
    .A2(net484),
    .A3(net479),
    .S0(clknet_1_1__leaf_net680),
    .S1(net682),
    .X(net499));
 sky130_fd_sc_hd__sdfrtp_1 c650 (.CLK(clknet_leaf_15_clk),
    .D(net497),
    .RESET_B(net499),
    .SCD(net494),
    .SCE(net681),
    .Q(net500));
 sky130_fd_sc_hd__buf_1 c651 (.A(net500),
    .X(net501));
 sky130_fd_sc_hd__buf_1 c652 (.A(net501),
    .X(net502));
 sky130_fd_sc_hd__and2_0 c653 (.A(net501),
    .B(net502),
    .X(net503));
 sky130_fd_sc_hd__dlymetal6s2s_1 c654 (.A(net624),
    .X(net504));
 sky130_fd_sc_hd__and2_1 c655 (.A(net406),
    .B(net502),
    .X(net505));
 sky130_fd_sc_hd__clkbuf_2 c656 (.A(net624),
    .X(net506));
 sky130_fd_sc_hd__and2_0 c657 (.A(net502),
    .B(net506),
    .X(net507));
 sky130_fd_sc_hd__dlrtp_1 c658 (.D(net507),
    .GATE(clknet_leaf_12_clk),
    .RESET_B(net506),
    .Q(net508));
 sky130_fd_sc_hd__dfbbn_1 c659 (.CLK_N(clknet_leaf_12_clk),
    .D(net490),
    .RESET_B(net507),
    .SET_B(net506),
    .Q(net509));
 sky130_fd_sc_hd__and3_1 c660 (.A(net506),
    .B(net501),
    .C(net504),
    .X(net510));
 sky130_fd_sc_hd__dfbbp_1 c661 (.CLK(clknet_leaf_12_clk),
    .D(net509),
    .RESET_B(net505),
    .SET_B(net849),
    .Q(net512),
    .Q_N(net511));
 sky130_fd_sc_hd__and3_1 c662 (.A(net508),
    .B(net506),
    .C(net504),
    .X(net513));
 sky130_fd_sc_hd__and3_1 c663 (.A(net510),
    .B(net512),
    .C(net513),
    .X(net514));
 sky130_fd_sc_hd__and3_1 c664 (.A(net512),
    .B(net513),
    .C(net508),
    .X(net515));
 sky130_fd_sc_hd__sdfxbp_1 c665 (.CLK(clknet_leaf_13_clk),
    .D(net380),
    .SCD(net904),
    .SCE(net504),
    .Q(net517),
    .Q_N(net516));
 sky130_fd_sc_hd__mux4_1 c666 (.A0(net492),
    .A1(net514),
    .A2(net511),
    .A3(net516),
    .S0(net513),
    .S1(net504),
    .X(net518));
 sky130_fd_sc_hd__sdfxbp_1 c667 (.CLK(clknet_leaf_13_clk),
    .D(net843),
    .SCD(net505),
    .SCE(net513),
    .Q(net519));
 sky130_fd_sc_hd__and3_1 c668 (.A(net513),
    .B(net919),
    .C(net506),
    .X(net520));
 sky130_fd_sc_hd__sdfxtp_1 c669 (.CLK(clknet_leaf_14_clk),
    .D(net501),
    .SCD(net520),
    .SCE(net505),
    .Q(net521));
 sky130_fd_sc_hd__and3_1 c670 (.A(net515),
    .B(net915),
    .C(net502),
    .X(net522));
 sky130_fd_sc_hd__sdfxtp_1 c671 (.CLK(clknet_leaf_13_clk),
    .D(net504),
    .SCD(net522),
    .SCE(net683),
    .Q(net523));
 sky130_fd_sc_hd__and2_1 c672 (.A(net422),
    .B(net523),
    .X(net524));
 sky130_fd_sc_hd__clkbuf_1 c673 (.X(net590));
 sky130_fd_sc_hd__buf_1 c674 (.A(net590),
    .X(net526));
 sky130_fd_sc_hd__dlrtp_1 c675 (.D(net482),
    .GATE(clknet_leaf_14_clk),
    .RESET_B(net525),
    .Q(net527));
 sky130_fd_sc_hd__and3_1 c676 (.A(net396),
    .B(net527),
    .C(net525),
    .X(net528));
 sky130_fd_sc_hd__and3_1 c677 (.A(net526),
    .B(net528),
    .C(net525),
    .X(net529));
 sky130_fd_sc_hd__and3_1 c678 (.A(clknet_1_1__leaf_net421),
    .B(net526),
    .C(net525),
    .X(net530));
 sky130_fd_sc_hd__and2_1 c679 (.A(net529),
    .B(net525),
    .X(net531));
 sky130_fd_sc_hd__dlrtp_1 c680 (.D(net531),
    .GATE(clknet_leaf_14_clk),
    .RESET_B(net525),
    .Q(net532));
 sky130_fd_sc_hd__sdfxtp_1 c681 (.CLK(clknet_leaf_13_clk),
    .D(net528),
    .SCD(net531),
    .SCE(net900),
    .Q(net533));
 sky130_fd_sc_hd__or4bb_2 c682 (.A(net532),
    .B(net528),
    .C_N(net533),
    .D_N(net525),
    .X(net534));
 sky130_fd_sc_hd__and3_1 c683 (.A(net529),
    .B(net534),
    .C(net527),
    .X(net535));
 sky130_fd_sc_hd__mux4_1 c684 (.A0(net527),
    .A1(net534),
    .A2(net533),
    .A3(net535),
    .S0(net525),
    .S1(net531),
    .X(net536));
 sky130_fd_sc_hd__mux4_1 c685 (.A0(clknet_1_0__leaf_net530),
    .A1(net532),
    .A2(net531),
    .A3(net527),
    .S0(net533),
    .S1(net525),
    .X(net537));
 sky130_fd_sc_hd__mux4_1 c686 (.A0(net534),
    .A1(net527),
    .A2(net533),
    .A3(net531),
    .S0(net524),
    .S1(net685),
    .X(net538));
 sky130_fd_sc_hd__mux4_1 c687 (.A0(net535),
    .A1(net527),
    .A2(net524),
    .A3(net525),
    .S0(net686),
    .S1(net687),
    .X(net539));
 sky130_fd_sc_hd__mux4_1 c688 (.A0(net534),
    .A1(net524),
    .A2(net525),
    .A3(net685),
    .S0(net687),
    .S1(net688),
    .X(net540));
 sky130_fd_sc_hd__mux4_1 c689 (.A0(net533),
    .A1(net531),
    .A2(net534),
    .A3(net686),
    .S0(net687),
    .S1(net689),
    .X(net541));
 sky130_fd_sc_hd__sdfbbn_1 c690 (.CLK_N(clknet_leaf_17_clk),
    .D(net524),
    .RESET_B(clknet_1_1__leaf_net530),
    .SCD(net525),
    .SCE(net687),
    .SET_B(net689),
    .Q(net543),
    .Q_N(net542));
 sky130_fd_sc_hd__mux4_1 c691 (.A0(net525),
    .A1(net535),
    .A2(net542),
    .A3(clknet_1_1__leaf_net530),
    .S0(net686),
    .S1(net687),
    .X(net544));
 sky130_fd_sc_hd__mux4_1 c692 (.A0(net543),
    .A1(clknet_1_0__leaf_net530),
    .A2(net525),
    .A3(net684),
    .S0(net687),
    .S1(net691),
    .X(net545));
 sky130_fd_sc_hd__clkbuf_2 c693 (.A(net627),
    .X(net546));
 sky130_fd_sc_hd__buf_1 c694 (.A(net546),
    .X(net547));
 sky130_fd_sc_hd__and2_0 c695 (.A(net546),
    .B(net547),
    .X(net548));
 sky130_fd_sc_hd__and2_0 c696 (.A(net546),
    .B(net692),
    .X(net549));
 sky130_fd_sc_hd__and2_1 c697 (.A(net414),
    .B(net547),
    .X(net550));
 sky130_fd_sc_hd__and2_1 c698 (.A(net546),
    .B(net550),
    .X(net551));
 sky130_fd_sc_hd__and2_1 c699 (.A(net549),
    .B(net546),
    .X(net552));
 sky130_fd_sc_hd__and2_1 c700 (.A(net547),
    .B(net548),
    .X(net553));
 sky130_fd_sc_hd__buf_1 c701 (.A(net918),
    .X(net554));
 sky130_fd_sc_hd__dfbbn_1 c702 (.CLK_N(clknet_leaf_17_clk),
    .D(net553),
    .RESET_B(net552),
    .SET_B(net554),
    .Q(net556),
    .Q_N(net555));
 sky130_fd_sc_hd__sdfrtp_1 c703 (.CLK(clknet_leaf_19_clk),
    .D(net547),
    .RESET_B(net553),
    .SCD(net548),
    .SCE(net546),
    .Q(net557));
 sky130_fd_sc_hd__and2_1 c704 (.A(net548),
    .B(net552),
    .X(net558));
 sky130_fd_sc_hd__dfbbn_1 c705 (.CLK_N(clknet_leaf_17_clk),
    .D(net552),
    .RESET_B(net558),
    .SET_B(net873),
    .Q(net560),
    .Q_N(net559));
 sky130_fd_sc_hd__sdfrtp_1 c706 (.CLK(clknet_leaf_17_clk),
    .D(net378),
    .RESET_B(net560),
    .SCD(net553),
    .SCE(net555),
    .Q(net561));
 sky130_fd_sc_hd__and2_0 c707 (.A(net556),
    .B(net690),
    .X(net562));
 sky130_fd_sc_hd__or4bb_1 c708 (.A(net562),
    .B(net560),
    .C_N(net555),
    .D_N(net557),
    .X(net563));
 sky130_fd_sc_hd__or4bb_1 c709 (.A(net914),
    .B(net555),
    .C_N(net563),
    .D_N(net688),
    .X(net564));
 sky130_fd_sc_hd__mux4_1 c710 (.A0(net922),
    .A1(net554),
    .A2(net556),
    .A3(net564),
    .S0(net547),
    .S1(net551),
    .X(net565));
 sky130_fd_sc_hd__sdfsbp_1 c711 (.CLK(clknet_leaf_16_clk),
    .D(net563),
    .SCD(net547),
    .SCE(net553),
    .SET_B(net824),
    .Q(net567),
    .Q_N(net566));
 sky130_fd_sc_hd__mux4_1 c712 (.A0(net564),
    .A1(net567),
    .A2(net559),
    .A3(net563),
    .S0(net558),
    .S1(net824),
    .X(net568));
 sky130_fd_sc_hd__sdfbbp_1 c713 (.CLK(clknet_leaf_16_clk),
    .D(net558),
    .RESET_B(net554),
    .SCD(net860),
    .SCE(net564),
    .SET_B(net826),
    .Q(net569));
 sky130_fd_sc_hd__clkbuf_1 c714 (.A(net550),
    .X(net570));
 sky130_fd_sc_hd__buf_1 c715 (.X(net594));
 sky130_fd_sc_hd__buf_1 c716 (.A(net593),
    .X(net572));
 sky130_fd_sc_hd__and2_1 c717 (.A(net572),
    .B(net571),
    .X(net573));
 sky130_fd_sc_hd__and2_2 c718 (.A(net571),
    .B(net573),
    .X(net574));
 sky130_fd_sc_hd__edfxbp_1 c719 (.CLK(clknet_leaf_16_clk),
    .D(net570),
    .DE(net573),
    .Q(net576),
    .Q_N(net575));
 sky130_fd_sc_hd__and3_1 c720 (.A(net576),
    .B(net571),
    .C(net574),
    .X(net577));
 sky130_fd_sc_hd__and2_1 c721 (.A(net573),
    .B(net575),
    .X(net578));
 sky130_fd_sc_hd__dfbbp_1 c722 (.CLK(clknet_leaf_16_clk),
    .D(net578),
    .RESET_B(net577),
    .SET_B(net572),
    .Q(net580),
    .Q_N(net579));
 sky130_fd_sc_hd__and3_1 c723 (.A(net574),
    .B(net579),
    .C(net571),
    .X(net581));
 sky130_fd_sc_hd__sdfxbp_1 c724 (.CLK(clknet_leaf_16_clk),
    .D(net851),
    .SCD(net581),
    .SCE(net578),
    .Q(net583),
    .Q_N(net582));
 sky130_fd_sc_hd__sdfxbp_1 c725 (.CLK(clknet_leaf_16_clk),
    .D(net794),
    .SCD(net580),
    .SCE(net577),
    .Q(net584));
 sky130_fd_sc_hd__and3_1 c726 (.A(net910),
    .B(net583),
    .C(net574),
    .X(net585));
 sky130_fd_sc_hd__sdfsbp_1 c727 (.CLK(clknet_leaf_16_clk),
    .D(net577),
    .SCD(net581),
    .SCE(net897),
    .SET_B(net574),
    .Q(net586));
 sky130_fd_sc_hd__sdfxtp_1 c728 (.CLK(clknet_leaf_16_clk),
    .D(net882),
    .SCD(net585),
    .SCE(net574),
    .Q(net587));
 sky130_fd_sc_hd__sdfxtp_1 c729 (.CLK(clknet_leaf_16_clk),
    .D(net585),
    .SCD(net855),
    .SCE(net572),
    .Q(net588));
 sky130_fd_sc_hd__and3_1 c730 (.A(net583),
    .B(net893),
    .C(net855),
    .X(net589));
 sky130_fd_sc_hd__sdfxtp_4 c731 (.CLK(clknet_leaf_16_clk),
    .D(net894),
    .SCD(net581),
    .SCE(net574));
 sky130_fd_sc_hd__edfxtp_1 merge732 (.CLK(clknet_leaf_18_clk),
    .D(net524),
    .Q(net590));
 sky130_fd_sc_hd__dfbbn_1 merge733 (.CLK_N(clknet_leaf_34_clk),
    .D(net817),
    .RESET_B(net807),
    .Q(net818),
    .Q_N(net591));
 sky130_fd_sc_hd__dfbbn_1 merge734 (.CLK_N(clknet_leaf_16_clk),
    .D(net569),
    .RESET_B(net570),
    .Q(net594),
    .Q_N(net593));
 sky130_fd_sc_hd__dfbbp_1 merge735 (.CLK(clknet_leaf_4_clk),
    .D(net380),
    .RESET_B(net377),
    .SET_B(net379),
    .Q(net596),
    .Q_N(net595));
 sky130_fd_sc_hd__mux4_1 merge736 (.A0(net61),
    .A1(net55),
    .A2(net56),
    .A3(net62),
    .S0(net737),
    .S1(clknet_1_0__leaf_net642),
    .X(net597));
 sky130_fd_sc_hd__sdfstp_1 merge737 (.CLK(clknet_leaf_6_clk),
    .D(net819),
    .SCD(net902),
    .SCE(net33),
    .SET_B(net707),
    .Q(net598));
 sky130_fd_sc_hd__sdfxbp_1 merge738 (.CLK(clknet_leaf_29_clk),
    .D(net801),
    .SCD(net312),
    .SCE(net314),
    .Q(net600),
    .Q_N(net599));
 sky130_fd_sc_hd__sdfstp_1 merge739 (.CLK(clknet_leaf_2_clk),
    .D(net75),
    .SCD(clknet_1_0__leaf_net170),
    .SCE(clknet_1_1__leaf_net174),
    .SET_B(clknet_1_0__leaf_net175),
    .Q(net601));
 sky130_fd_sc_hd__sdlclkp_1 merge740 (.CLK(clknet_leaf_27_clk),
    .GATE(net101),
    .SCE(net864),
    .GCLK(net602));
 sky130_fd_sc_hd__sdfbbn_2 merge741 (.CLK_N(clknet_leaf_8_clk),
    .D(net28),
    .RESET_B(net768),
    .SCD(net125),
    .SCE(net126),
    .Q(net122),
    .Q_N(net603));
 sky130_fd_sc_hd__sdfxbp_1 merge742 (.CLK(clknet_leaf_20_clk),
    .D(net443),
    .SCD(clknet_1_1__leaf_net455),
    .SCE(net457),
    .Q(net606),
    .Q_N(net605));
 sky130_fd_sc_hd__sdfstp_1 merge743 (.CLK(clknet_leaf_14_clk),
    .D(net483),
    .SCD(net480),
    .SCE(net482),
    .Q(net484));
 sky130_fd_sc_hd__sedfxbp_1 merge744 (.CLK(clknet_leaf_23_clk),
    .D(net335),
    .DE(net805),
    .SCE(net792),
    .Q(net800),
    .Q_N(net608));
 sky130_fd_sc_hd__sdlclkp_2 merge745 (.CLK(clknet_leaf_30_clk),
    .GATE(clknet_1_0__leaf_net288),
    .GCLK(net289));
 sky130_fd_sc_hd__sdfxtp_1 merge746 (.CLK(clknet_leaf_9_clk),
    .D(net4),
    .SCD(net6),
    .SCE(net7),
    .Q(net611));
 sky130_fd_sc_hd__sdfxtp_1 merge747 (.CLK(clknet_leaf_2_clk),
    .D(net262),
    .SCD(net263),
    .Q(net264));
 sky130_fd_sc_hd__sdfxtp_1 merge748 (.CLK(clknet_leaf_26_clk),
    .D(net880),
    .SCD(net221),
    .Q(net613));
 sky130_fd_sc_hd__dfbbn_1 merge749 (.CLK_N(clknet_leaf_28_clk),
    .D(net196),
    .RESET_B(net195),
    .SET_B(net202),
    .Q(net615),
    .Q_N(net614));
 sky130_fd_sc_hd__dfbbn_1 merge750 (.CLK_N(clknet_leaf_7_clk),
    .D(net239),
    .RESET_B(net238),
    .Q(net240),
    .Q_N(net616));
 sky130_fd_sc_hd__sedfxbp_2 merge751 (.CLK(clknet_leaf_5_clk),
    .D(net147),
    .DE(net146),
    .SCD(net149),
    .Q(net148),
    .Q_N(net618));
 sky130_fd_sc_hd__dfbbp_1 merge752 (.CLK(clknet_leaf_10_clk),
    .D(net354),
    .RESET_B(net353),
    .SET_B(net833),
    .Q(net621),
    .Q_N(net620));
 sky130_fd_sc_hd__sdfxbp_1 merge753 (.CLK(clknet_leaf_33_clk),
    .D(net78),
    .SCD(net753),
    .SCE(net79),
    .Q(net623),
    .Q_N(net622));
 sky130_fd_sc_hd__sedfxtp_1 merge754 (.CLK(clknet_leaf_14_clk),
    .D(net503),
    .DE(net502),
    .SCD(net505),
    .SCE(net501),
    .Q(net624));
 sky130_fd_sc_hd__sdfxbp_1 merge755 (.CLK(clknet_leaf_19_clk),
    .D(net434),
    .SCD(net432),
    .SCE(clknet_1_0__leaf_net433),
    .Q(net626),
    .Q_N(net625));
 sky130_fd_sc_hd__sedfxtp_1 merge756 (.CLK(clknet_leaf_21_clk),
    .D(clknet_1_1__leaf_net433),
    .DE(net551),
    .SCD(net553),
    .SCE(net550),
    .Q(net627));
 sky130_fd_sc_hd__sedfxtp_1 merge757 (.CLK(clknet_leaf_30_clk),
    .D(clknet_1_1__leaf_net175),
    .DE(net407),
    .SCD(net861),
    .SCE(net412),
    .Q(net628));
 sky130_fd_sc_hd__sdfrbp_1 merge758 (.CLK(clknet_leaf_29_clk),
    .D(net313),
    .RESET_B(net317),
    .SCD(net198),
    .SCE(net197),
    .Q(net630),
    .Q_N(net629));
 sky130_fd_sc_hd__sdfrbp_1 merge759 (.CLK(clknet_leaf_28_clk),
    .D(clknet_1_0__leaf_net102),
    .RESET_B(net101),
    .SCD(net79),
    .SCE(net83),
    .Q(net632),
    .Q_N(net631));
 sky130_fd_sc_hd__sdfrtn_1 merge760 (.CLK_N(clknet_leaf_29_clk),
    .D(clknet_1_1__leaf_net288),
    .RESET_B(clknet_1_1__leaf_net289),
    .SCD(net315),
    .SCE(net320),
    .Q(net633));
 sky130_fd_sc_hd__sdfrtp_1 merge761 (.CLK(clknet_leaf_23_clk),
    .D(net337),
    .RESET_B(net823),
    .SCD(net463),
    .SCE(clknet_1_0__leaf_net455),
    .Q(net634));
 sky130_fd_sc_hd__dfxbp_1 s762 (.CLK(clknet_leaf_8_clk),
    .D(net25),
    .Q(net636),
    .Q_N(net635));
 sky130_fd_sc_hd__dfxbp_1 s763 (.CLK(clknet_leaf_5_clk),
    .D(net48),
    .Q(net638),
    .Q_N(net637));
 sky130_fd_sc_hd__dfxtp_1 s764 (.CLK(clknet_leaf_0_clk),
    .D(net51),
    .Q(net639));
 sky130_fd_sc_hd__dfxtp_1 s765 (.CLK(clknet_leaf_0_clk),
    .D(net53),
    .Q(net640));
 sky130_fd_sc_hd__dfxtp_1 s766 (.CLK(clknet_leaf_0_clk),
    .D(net876),
    .Q(net641));
 sky130_fd_sc_hd__dlclkp_1 s767 (.CLK(clknet_leaf_35_clk),
    .GATE(net67),
    .GCLK(net642));
 sky130_fd_sc_hd__dlclkp_2 s768 (.CLK(clknet_leaf_35_clk),
    .GATE(net73),
    .GCLK(net643));
 sky130_fd_sc_hd__dlclkp_4 s769 (.CLK(clknet_leaf_32_clk),
    .GATE(net99),
    .GCLK(net644));
 sky130_fd_sc_hd__dlxbn_1 s770 (.D(net116),
    .GATE_N(clknet_leaf_24_clk),
    .Q(net810),
    .Q_N(net812));
 sky130_fd_sc_hd__dlxbn_1 s771 (.D(net139),
    .GATE_N(clknet_leaf_7_clk),
    .Q(net646),
    .Q_N(net645));
 sky130_fd_sc_hd__dlxbp_1 s772 (.D(net143),
    .GATE(clknet_leaf_7_clk),
    .Q(net648),
    .Q_N(net647));
 sky130_fd_sc_hd__dlxtn_1 s773 (.D(net161),
    .GATE_N(clknet_leaf_4_clk),
    .Q(net649));
 sky130_fd_sc_hd__dlxtn_1 s774 (.D(net181),
    .GATE_N(clknet_leaf_31_clk),
    .Q(net650));
 sky130_fd_sc_hd__dlxtn_1 s775 (.D(net192),
    .GATE_N(clknet_leaf_31_clk),
    .Q(net651));
 sky130_fd_sc_hd__dlxtp_1 s776 (.D(net193),
    .GATE(clknet_leaf_32_clk),
    .Q(net652));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s777 (.D(net217),
    .SLEEP_B(clknet_leaf_29_clk),
    .Q(net653));
 sky130_fd_sc_hd__dfxbp_1 s778 (.CLK(clknet_leaf_25_clk),
    .D(net233),
    .Q(net655),
    .Q_N(net654));
 sky130_fd_sc_hd__dfxbp_1 s779 (.CLK(clknet_leaf_24_clk),
    .D(net234),
    .Q(net657),
    .Q_N(net656));
 sky130_fd_sc_hd__dfxtp_1 s780 (.CLK(clknet_leaf_25_clk),
    .D(net236),
    .Q(net658));
 sky130_fd_sc_hd__dfxtp_1 s781 (.CLK(clknet_leaf_4_clk),
    .D(net253),
    .Q(net659));
 sky130_fd_sc_hd__dfxtp_1 s782 (.CLK(clknet_leaf_2_clk),
    .D(net284),
    .Q(net660));
 sky130_fd_sc_hd__dlclkp_1 s783 (.CLK(clknet_leaf_30_clk),
    .GATE(net286),
    .GCLK(net661));
 sky130_fd_sc_hd__dlclkp_2 s784 (.CLK(clknet_leaf_18_clk),
    .GATE(net303),
    .GCLK(net662));
 sky130_fd_sc_hd__dlclkp_4 s785 (.CLK(clknet_leaf_20_clk),
    .GATE(net325),
    .GCLK(net663));
 sky130_fd_sc_hd__dlxbn_1 s786 (.D(net328),
    .GATE_N(clknet_leaf_26_clk),
    .Q(net665),
    .Q_N(net664));
 sky130_fd_sc_hd__dlxbn_1 s787 (.D(net329),
    .GATE_N(clknet_leaf_20_clk),
    .Q(net667),
    .Q_N(net666));
 sky130_fd_sc_hd__dlxbp_1 s788 (.D(net330),
    .GATE(clknet_leaf_23_clk),
    .Q(net668),
    .Q_N(net799));
 sky130_fd_sc_hd__dlxtn_1 s789 (.D(net331),
    .GATE_N(clknet_leaf_23_clk),
    .Q(net792));
 sky130_fd_sc_hd__dlxtn_1 s790 (.D(net332),
    .GATE_N(clknet_leaf_23_clk),
    .Q(net669));
 sky130_fd_sc_hd__dlxtn_1 s791 (.D(net375),
    .GATE_N(clknet_leaf_11_clk),
    .Q(net670));
 sky130_fd_sc_hd__dlxtp_1 s792 (.D(net376),
    .GATE(clknet_leaf_11_clk),
    .Q(net671));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s793 (.D(net404),
    .SLEEP_B(clknet_leaf_3_clk),
    .Q(net672));
 sky130_fd_sc_hd__dfxbp_1 s794 (.CLK(clknet_leaf_18_clk),
    .D(net427),
    .Q(net674),
    .Q_N(net673));
 sky130_fd_sc_hd__dfxbp_1 s795 (.CLK(clknet_leaf_19_clk),
    .D(net429),
    .Q(net675));
 sky130_fd_sc_hd__dfxtp_1 s796 (.CLK(clknet_leaf_20_clk),
    .D(net452),
    .Q(net676));
 sky130_fd_sc_hd__dfxtp_1 s797 (.CLK(clknet_leaf_20_clk),
    .D(net453),
    .Q(net677));
 sky130_fd_sc_hd__dfxtp_1 s798 (.CLK(clknet_leaf_22_clk),
    .D(net473),
    .Q(net678));
 sky130_fd_sc_hd__dlclkp_1 s799 (.CLK(clknet_leaf_22_clk),
    .GATE(net474),
    .GCLK(net679));
 sky130_fd_sc_hd__dlclkp_2 s800 (.CLK(clknet_leaf_22_clk),
    .GATE(net478),
    .GCLK(net796));
 sky130_fd_sc_hd__dlclkp_4 s801 (.CLK(clknet_leaf_15_clk),
    .GATE(net495),
    .GCLK(net680));
 sky130_fd_sc_hd__dlxbn_1 s802 (.D(net498),
    .GATE_N(clknet_leaf_15_clk),
    .Q(net682),
    .Q_N(net681));
 sky130_fd_sc_hd__dlxbn_1 s803 (.D(net518),
    .GATE_N(clknet_leaf_13_clk),
    .Q(net683));
 sky130_fd_sc_hd__dlxbp_1 s804 (.D(net536),
    .GATE(clknet_leaf_14_clk),
    .Q(net685),
    .Q_N(net684));
 sky130_fd_sc_hd__dlxtn_1 s805 (.D(net537),
    .GATE_N(clknet_leaf_14_clk),
    .Q(net686));
 sky130_fd_sc_hd__dlxtn_2 s806 (.D(net538),
    .GATE_N(clknet_leaf_14_clk),
    .Q(net687));
 sky130_fd_sc_hd__dlxtn_1 s807 (.D(net539),
    .GATE_N(clknet_leaf_18_clk),
    .Q(net688));
 sky130_fd_sc_hd__dlxtp_1 s808 (.D(net540),
    .GATE(clknet_leaf_17_clk),
    .Q(net689));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s809 (.D(net541),
    .SLEEP_B(clknet_leaf_17_clk),
    .Q(net690));
 sky130_fd_sc_hd__dfxbp_1 s810 (.CLK(clknet_leaf_17_clk),
    .D(net544),
    .Q(net691));
 sky130_fd_sc_hd__dfxbp_1 s811 (.CLK(clknet_leaf_17_clk),
    .D(net545),
    .Q(net692));
 sky130_fd_sc_hd__dfxtp_1 s812 (.CLK(clknet_leaf_21_clk),
    .D(net565),
    .Q(net693));
 sky130_fd_sc_hd__dfxtp_1 s813 (.CLK(clknet_leaf_16_clk),
    .D(net568),
    .Q(net694));
 sky130_fd_sc_hd__dfxtp_1 s814 (.CLK(clknet_leaf_35_clk),
    .D(net597),
    .Q(net695));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Right_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Right_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Right_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Right_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Right_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Right_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Right_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Right_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Right_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Right_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Right_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Right_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Right_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Right_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Right_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Right_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Right_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Right_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Right_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Right_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Right_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_161 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_162 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_163 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_164 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_165 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_166 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_167 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_168 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_169 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_170 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_171 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_172 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_173 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_174 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_175 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_176 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_177 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_178 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_179 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_180 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_181 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_182 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Left_183 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Left_184 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Left_185 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Left_186 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Left_187 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Left_188 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Left_189 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Left_190 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Left_191 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Left_192 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Left_193 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Left_194 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Left_195 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Left_196 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Left_197 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Left_198 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Left_199 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Left_200 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Left_201 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Left_202 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Left_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1347 ();
 sky130_fd_sc_hd__buf_1 input1 (.A(in0),
    .X(net592));
 sky130_fd_sc_hd__buf_1 input2 (.A(in1),
    .X(net604));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(in10),
    .X(net609));
 sky130_fd_sc_hd__buf_1 input4 (.A(in11),
    .X(net617));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(in12),
    .X(net619));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(in13),
    .X(net696));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(in14),
    .X(net697));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(in15),
    .X(net698));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(in16),
    .X(net699));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(in17),
    .X(net700));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(in18),
    .X(net701));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(in19),
    .X(net702));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(in2),
    .X(net703));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(in20),
    .X(net704));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(in21),
    .X(net705));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(in22),
    .X(net706));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(in23),
    .X(net707));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(in24),
    .X(net708));
 sky130_fd_sc_hd__clkbuf_1 input19 (.A(in25),
    .X(net709));
 sky130_fd_sc_hd__buf_1 input20 (.A(in26),
    .X(net710));
 sky130_fd_sc_hd__clkbuf_1 input21 (.A(in27),
    .X(net711));
 sky130_fd_sc_hd__clkbuf_1 input22 (.A(in28),
    .X(net712));
 sky130_fd_sc_hd__clkbuf_1 input23 (.A(in29),
    .X(net713));
 sky130_fd_sc_hd__clkbuf_1 input24 (.A(in3),
    .X(net714));
 sky130_fd_sc_hd__clkbuf_1 input25 (.A(in30),
    .X(net715));
 sky130_fd_sc_hd__clkbuf_1 input26 (.A(in31),
    .X(net716));
 sky130_fd_sc_hd__clkbuf_1 input27 (.A(in32),
    .X(net717));
 sky130_fd_sc_hd__clkbuf_1 input28 (.A(in33),
    .X(net718));
 sky130_fd_sc_hd__clkbuf_1 input29 (.A(in34),
    .X(net719));
 sky130_fd_sc_hd__clkbuf_1 input30 (.A(in35),
    .X(net720));
 sky130_fd_sc_hd__clkbuf_1 input31 (.A(in36),
    .X(net721));
 sky130_fd_sc_hd__clkbuf_1 input32 (.A(in37),
    .X(net722));
 sky130_fd_sc_hd__clkbuf_1 input33 (.A(in38),
    .X(net723));
 sky130_fd_sc_hd__clkbuf_1 input34 (.A(in39),
    .X(net724));
 sky130_fd_sc_hd__clkbuf_1 input35 (.A(in4),
    .X(net725));
 sky130_fd_sc_hd__clkbuf_1 input36 (.A(in40),
    .X(net726));
 sky130_fd_sc_hd__clkbuf_1 input37 (.A(in41),
    .X(net727));
 sky130_fd_sc_hd__clkbuf_1 input38 (.A(in42),
    .X(net728));
 sky130_fd_sc_hd__clkbuf_1 input39 (.A(in43),
    .X(net729));
 sky130_fd_sc_hd__clkbuf_1 input40 (.A(in44),
    .X(net730));
 sky130_fd_sc_hd__buf_1 input41 (.A(in45),
    .X(net731));
 sky130_fd_sc_hd__clkbuf_1 input42 (.A(in46),
    .X(net732));
 sky130_fd_sc_hd__clkbuf_1 input43 (.A(in47),
    .X(net733));
 sky130_fd_sc_hd__clkbuf_1 input44 (.A(in48),
    .X(net734));
 sky130_fd_sc_hd__buf_1 input45 (.A(in49),
    .X(net735));
 sky130_fd_sc_hd__clkbuf_1 input46 (.A(in5),
    .X(net736));
 sky130_fd_sc_hd__clkbuf_1 input47 (.A(in50),
    .X(net737));
 sky130_fd_sc_hd__clkbuf_1 input48 (.A(in51),
    .X(net738));
 sky130_fd_sc_hd__buf_1 input49 (.A(in52),
    .X(net739));
 sky130_fd_sc_hd__clkbuf_1 input50 (.A(in53),
    .X(net740));
 sky130_fd_sc_hd__clkbuf_1 input51 (.A(in54),
    .X(net741));
 sky130_fd_sc_hd__clkbuf_1 input52 (.A(in55),
    .X(net742));
 sky130_fd_sc_hd__clkbuf_1 input53 (.A(in56),
    .X(net743));
 sky130_fd_sc_hd__clkbuf_1 input54 (.A(in57),
    .X(net744));
 sky130_fd_sc_hd__clkbuf_1 input55 (.A(in58),
    .X(net745));
 sky130_fd_sc_hd__buf_1 input56 (.A(in59),
    .X(net746));
 sky130_fd_sc_hd__clkbuf_1 input57 (.A(in6),
    .X(net747));
 sky130_fd_sc_hd__clkbuf_1 input58 (.A(in60),
    .X(net748));
 sky130_fd_sc_hd__clkbuf_1 input59 (.A(in61),
    .X(net749));
 sky130_fd_sc_hd__clkbuf_1 input60 (.A(in62),
    .X(net750));
 sky130_fd_sc_hd__clkbuf_1 input61 (.A(in63),
    .X(net751));
 sky130_fd_sc_hd__clkbuf_1 input62 (.A(in64),
    .X(net752));
 sky130_fd_sc_hd__buf_1 input63 (.A(in65),
    .X(net753));
 sky130_fd_sc_hd__buf_1 input64 (.A(in66),
    .X(net754));
 sky130_fd_sc_hd__clkbuf_1 input65 (.A(in67),
    .X(net755));
 sky130_fd_sc_hd__clkbuf_1 input66 (.A(in68),
    .X(net756));
 sky130_fd_sc_hd__clkbuf_1 input67 (.A(in69),
    .X(net757));
 sky130_fd_sc_hd__clkbuf_1 input68 (.A(in7),
    .X(net758));
 sky130_fd_sc_hd__buf_1 input69 (.A(in70),
    .X(net759));
 sky130_fd_sc_hd__clkbuf_1 input70 (.A(in71),
    .X(net760));
 sky130_fd_sc_hd__clkbuf_1 input71 (.A(in72),
    .X(net761));
 sky130_fd_sc_hd__clkbuf_1 input72 (.A(in74),
    .X(net762));
 sky130_fd_sc_hd__clkbuf_1 input73 (.A(in75),
    .X(net763));
 sky130_fd_sc_hd__clkbuf_1 input74 (.A(in76),
    .X(net764));
 sky130_fd_sc_hd__clkbuf_1 input75 (.A(in77),
    .X(net765));
 sky130_fd_sc_hd__clkbuf_1 input76 (.A(in78),
    .X(net766));
 sky130_fd_sc_hd__clkbuf_1 input77 (.A(in79),
    .X(net767));
 sky130_fd_sc_hd__clkbuf_1 input78 (.A(in8),
    .X(net768));
 sky130_fd_sc_hd__clkbuf_1 input79 (.A(in80),
    .X(net769));
 sky130_fd_sc_hd__clkbuf_1 input80 (.A(in81),
    .X(net770));
 sky130_fd_sc_hd__clkbuf_1 input81 (.A(in82),
    .X(net771));
 sky130_fd_sc_hd__clkbuf_1 input82 (.A(in83),
    .X(net772));
 sky130_fd_sc_hd__clkbuf_1 input83 (.A(in84),
    .X(net773));
 sky130_fd_sc_hd__clkbuf_1 input84 (.A(in85),
    .X(net774));
 sky130_fd_sc_hd__clkbuf_1 input85 (.A(in86),
    .X(net775));
 sky130_fd_sc_hd__clkbuf_1 input86 (.A(in87),
    .X(net776));
 sky130_fd_sc_hd__clkbuf_1 input87 (.A(in88),
    .X(net777));
 sky130_fd_sc_hd__clkbuf_1 input88 (.A(in89),
    .X(net778));
 sky130_fd_sc_hd__clkbuf_1 input89 (.A(in9),
    .X(net779));
 sky130_fd_sc_hd__buf_1 input90 (.A(in90),
    .X(net780));
 sky130_fd_sc_hd__clkbuf_1 input91 (.A(in91),
    .X(net781));
 sky130_fd_sc_hd__clkbuf_1 input92 (.A(in92),
    .X(net782));
 sky130_fd_sc_hd__buf_1 input93 (.A(in93),
    .X(net783));
 sky130_fd_sc_hd__clkbuf_1 input94 (.A(in94),
    .X(net784));
 sky130_fd_sc_hd__clkbuf_1 input95 (.A(in95),
    .X(net785));
 sky130_fd_sc_hd__clkbuf_1 input96 (.A(in96),
    .X(net786));
 sky130_fd_sc_hd__dlymetal6s2s_1 input97 (.A(in97),
    .X(net787));
 sky130_fd_sc_hd__clkbuf_1 input98 (.A(in98),
    .X(net788));
 sky130_fd_sc_hd__clkbuf_1 input99 (.A(in99),
    .X(net789));
 sky130_fd_sc_hd__buf_2 output100 (.A(net790),
    .X(out10));
 sky130_fd_sc_hd__buf_2 output101 (.A(net791),
    .X(out19));
 sky130_fd_sc_hd__buf_2 output102 (.A(net792),
    .X(out21));
 sky130_fd_sc_hd__buf_2 output103 (.A(net793),
    .X(out23));
 sky130_fd_sc_hd__buf_2 output104 (.A(net794),
    .X(out25));
 sky130_fd_sc_hd__buf_2 output105 (.A(net795),
    .X(out26));
 sky130_fd_sc_hd__clkbuf_1 output106 (.A(net796),
    .X(out3));
 sky130_fd_sc_hd__buf_2 output107 (.A(net797),
    .X(out32));
 sky130_fd_sc_hd__buf_2 output108 (.A(net798),
    .X(out33));
 sky130_fd_sc_hd__buf_2 output109 (.A(net799),
    .X(out35));
 sky130_fd_sc_hd__buf_2 output110 (.A(net800),
    .X(out36));
 sky130_fd_sc_hd__buf_2 output111 (.A(net801),
    .X(out44));
 sky130_fd_sc_hd__buf_2 output112 (.A(net802),
    .X(out47));
 sky130_fd_sc_hd__buf_2 output113 (.A(net803),
    .X(out49));
 sky130_fd_sc_hd__buf_2 output114 (.A(net804),
    .X(out50));
 sky130_fd_sc_hd__buf_2 output115 (.A(net805),
    .X(out54));
 sky130_fd_sc_hd__clkbuf_1 output116 (.A(clknet_1_0__leaf_net806),
    .X(out65));
 sky130_fd_sc_hd__buf_2 output117 (.A(net807),
    .X(out66));
 sky130_fd_sc_hd__buf_2 output118 (.A(net808),
    .X(out70));
 sky130_fd_sc_hd__buf_2 output119 (.A(net809),
    .X(out71));
 sky130_fd_sc_hd__buf_2 output120 (.A(net810),
    .X(out73));
 sky130_fd_sc_hd__buf_2 output121 (.A(net811),
    .X(out79));
 sky130_fd_sc_hd__buf_2 output122 (.A(net812),
    .X(out80));
 sky130_fd_sc_hd__buf_2 output123 (.A(net813),
    .X(out83));
 sky130_fd_sc_hd__buf_2 output124 (.A(net814),
    .X(out84));
 sky130_fd_sc_hd__buf_2 output125 (.A(net815),
    .X(out92));
 sky130_fd_sc_hd__buf_2 output126 (.A(net816),
    .X(out93));
 sky130_fd_sc_hd__buf_2 output127 (.A(net817),
    .X(out94));
 sky130_fd_sc_hd__buf_2 output128 (.A(net818),
    .X(out98));
 sky130_fd_sc_hd__clkbuf_4 fanout129 (.A(net34),
    .X(net819));
 sky130_fd_sc_hd__clkbuf_2 fanout130 (.A(net821),
    .X(net820));
 sky130_fd_sc_hd__clkbuf_2 fanout131 (.A(net122),
    .X(net821));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_0_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_1_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_2_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_3_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_4_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_5_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_6_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_7_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_8_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_9_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_9_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_10_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_11_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_12_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_13_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_14_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_15_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_16_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_17_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_18_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_19_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_20_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_21_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_22_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_22_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_23_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_24_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_24_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_25_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_25_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_26_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_26_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_27_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_27_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_28_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_28_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_29_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_29_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_30_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_30_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_31_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_31_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_32_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_32_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_33_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_33_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_34_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_34_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_35_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_35_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net680 (.A(net680),
    .X(clknet_0_net680));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net680 (.A(clknet_0_net680),
    .X(clknet_1_0__leaf_net680));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net680 (.A(clknet_0_net680),
    .X(clknet_1_1__leaf_net680));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net679 (.A(net679),
    .X(clknet_0_net679));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net679 (.A(clknet_0_net679),
    .X(clknet_1_0__leaf_net679));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net679 (.A(clknet_0_net679),
    .X(clknet_1_1__leaf_net679));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net663 (.A(net663),
    .X(clknet_0_net663));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net663 (.A(clknet_0_net663),
    .X(clknet_1_0__leaf_net663));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net663 (.A(clknet_0_net663),
    .X(clknet_1_1__leaf_net663));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net327 (.A(net327),
    .X(clknet_0_net327));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net327 (.A(clknet_0_net327),
    .X(clknet_1_0__leaf_net327));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net327 (.A(clknet_0_net327),
    .X(clknet_1_1__leaf_net327));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net662 (.A(net662),
    .X(clknet_0_net662));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net662 (.A(clknet_0_net662),
    .X(clknet_1_0__leaf_net662));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net662 (.A(clknet_0_net662),
    .X(clknet_1_1__leaf_net662));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net419 (.A(net419),
    .X(clknet_0_net419));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net419 (.A(clknet_0_net419),
    .X(clknet_1_0__leaf_net419));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net419 (.A(clknet_0_net419),
    .X(clknet_1_1__leaf_net419));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net454 (.A(net454),
    .X(clknet_0_net454));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net454 (.A(clknet_0_net454),
    .X(clknet_1_0__leaf_net454));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net454 (.A(clknet_0_net454),
    .X(clknet_1_1__leaf_net454));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net455 (.A(net455),
    .X(clknet_0_net455));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net455 (.A(clknet_0_net455),
    .X(clknet_1_0__leaf_net455));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net455 (.A(clknet_0_net455),
    .X(clknet_1_1__leaf_net455));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net433 (.A(net433),
    .X(clknet_0_net433));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net433 (.A(clknet_0_net433),
    .X(clknet_1_0__leaf_net433));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net433 (.A(clknet_0_net433),
    .X(clknet_1_1__leaf_net433));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net421 (.A(net421),
    .X(clknet_0_net421));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net421 (.A(clknet_0_net421),
    .X(clknet_1_0__leaf_net421));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net421 (.A(clknet_0_net421),
    .X(clknet_1_1__leaf_net421));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net530 (.A(net530),
    .X(clknet_0_net530));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net530 (.A(clknet_0_net530),
    .X(clknet_1_0__leaf_net530));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net530 (.A(clknet_0_net530),
    .X(clknet_1_1__leaf_net530));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net423 (.A(net423),
    .X(clknet_0_net423));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net423 (.A(clknet_0_net423),
    .X(clknet_1_0__leaf_net423));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net423 (.A(clknet_0_net423),
    .X(clknet_1_1__leaf_net423));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net309 (.A(net309),
    .X(clknet_0_net309));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net309 (.A(clknet_0_net309),
    .X(clknet_1_0__leaf_net309));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net309 (.A(clknet_0_net309),
    .X(clknet_1_1__leaf_net309));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net288 (.A(net288),
    .X(clknet_0_net288));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net288 (.A(clknet_0_net288),
    .X(clknet_1_0__leaf_net288));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net288 (.A(clknet_0_net288),
    .X(clknet_1_1__leaf_net288));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net289 (.A(net289),
    .X(clknet_0_net289));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net289 (.A(clknet_0_net289),
    .X(clknet_1_0__leaf_net289));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net289 (.A(clknet_0_net289),
    .X(clknet_1_1__leaf_net289));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net643 (.A(net643),
    .X(clknet_0_net643));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net643 (.A(clknet_0_net643),
    .X(clknet_1_0__leaf_net643));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net643 (.A(clknet_0_net643),
    .X(clknet_1_1__leaf_net643));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net170 (.A(net170),
    .X(clknet_0_net170));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net170 (.A(clknet_0_net170),
    .X(clknet_1_0__leaf_net170));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net170 (.A(clknet_0_net170),
    .X(clknet_1_1__leaf_net170));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net184 (.A(net184),
    .X(clknet_0_net184));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net184 (.A(clknet_0_net184),
    .X(clknet_1_0__leaf_net184));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net184 (.A(clknet_0_net184),
    .X(clknet_1_1__leaf_net184));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net178 (.A(net178),
    .X(clknet_0_net178));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net178 (.A(clknet_0_net178),
    .X(clknet_1_0__leaf_net178));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net178 (.A(clknet_0_net178),
    .X(clknet_1_1__leaf_net178));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net175 (.A(net175),
    .X(clknet_0_net175));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net175 (.A(clknet_0_net175),
    .X(clknet_1_0__leaf_net175));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net175 (.A(clknet_0_net175),
    .X(clknet_1_1__leaf_net175));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net174 (.A(net174),
    .X(clknet_0_net174));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net174 (.A(clknet_0_net174),
    .X(clknet_1_0__leaf_net174));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net174 (.A(clknet_0_net174),
    .X(clknet_1_1__leaf_net174));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net173 (.A(net173),
    .X(clknet_0_net173));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net173 (.A(clknet_0_net173),
    .X(clknet_1_0__leaf_net173));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net173 (.A(clknet_0_net173),
    .X(clknet_1_1__leaf_net173));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net206 (.A(net206),
    .X(clknet_0_net206));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net206 (.A(clknet_0_net206),
    .X(clknet_1_0__leaf_net206));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net206 (.A(clknet_0_net206),
    .X(clknet_1_1__leaf_net206));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net185 (.A(net185),
    .X(clknet_0_net185));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net185 (.A(clknet_0_net185),
    .X(clknet_1_0__leaf_net185));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net185 (.A(clknet_0_net185),
    .X(clknet_1_1__leaf_net185));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net642 (.A(net642),
    .X(clknet_0_net642));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net642 (.A(clknet_0_net642),
    .X(clknet_1_0__leaf_net642));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net642 (.A(clknet_0_net642),
    .X(clknet_1_1__leaf_net642));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net602 (.A(net602),
    .X(clknet_0_net602));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net602 (.A(clknet_0_net602),
    .X(clknet_1_0__leaf_net602));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net602 (.A(clknet_0_net602),
    .X(clknet_1_1__leaf_net602));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net105 (.A(net105),
    .X(clknet_0_net105));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net105 (.A(clknet_0_net105),
    .X(clknet_1_0__leaf_net105));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net105 (.A(clknet_0_net105),
    .X(clknet_1_1__leaf_net105));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net806 (.A(net806),
    .X(clknet_0_net806));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net806 (.A(clknet_0_net806),
    .X(clknet_1_0__leaf_net806));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net806 (.A(clknet_0_net806),
    .X(clknet_1_1__leaf_net806));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net102 (.A(net102),
    .X(clknet_0_net102));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net102 (.A(clknet_0_net102),
    .X(clknet_1_0__leaf_net102));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net102 (.A(clknet_0_net102),
    .X(clknet_1_1__leaf_net102));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net106 (.A(net106),
    .X(clknet_0_net106));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net106 (.A(clknet_0_net106),
    .X(clknet_1_0__leaf_net106));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net106 (.A(clknet_0_net106),
    .X(clknet_1_1__leaf_net106));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net113 (.A(net113),
    .X(clknet_0_net113));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net113 (.A(clknet_0_net113),
    .X(clknet_1_0__leaf_net113));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net113 (.A(clknet_0_net113),
    .X(clknet_1_1__leaf_net113));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net111 (.A(net111),
    .X(clknet_0_net111));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net111 (.A(clknet_0_net111),
    .X(clknet_1_0__leaf_net111));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net111 (.A(clknet_0_net111),
    .X(clknet_1_1__leaf_net111));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net112 (.A(net112),
    .X(clknet_0_net112));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net112 (.A(clknet_0_net112),
    .X(clknet_1_0__leaf_net112));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net112 (.A(clknet_0_net112),
    .X(clknet_1_1__leaf_net112));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net108 (.A(net108),
    .X(clknet_0_net108));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net108 (.A(clknet_0_net108),
    .X(clknet_1_0__leaf_net108));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net108 (.A(clknet_0_net108),
    .X(clknet_1_1__leaf_net108));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net118 (.A(net118),
    .X(clknet_0_net118));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net118 (.A(clknet_0_net118),
    .X(clknet_1_0__leaf_net118));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net118 (.A(clknet_0_net118),
    .X(clknet_1_1__leaf_net118));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer1 (.A(net89),
    .X(net822));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(net800),
    .X(net823));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(net693),
    .X(net824));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(net117),
    .X(net825));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(net694),
    .X(net826));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(net598),
    .X(net827));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(net488),
    .X(net828));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(net416),
    .X(net829));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(net638),
    .X(net830));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(net119),
    .X(net831));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(net155),
    .X(net832));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(net242),
    .X(net833));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(net613),
    .X(net834));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(net461),
    .X(net835));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(net468),
    .X(net836));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(net399),
    .X(net837));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(net299),
    .X(net838));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(net281),
    .X(net839));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(net471),
    .X(net840));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(net646),
    .X(net841));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(net649),
    .X(net842));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(net517),
    .X(net843));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(net342),
    .X(net844));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(net9),
    .X(net845));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(net279),
    .X(net846));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(net168),
    .X(net847));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(net469),
    .X(net848));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(net506),
    .X(net849));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(net413),
    .X(net850));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(net576),
    .X(net851));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(net347),
    .X(net852));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(net634),
    .X(net853));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(net393),
    .X(net854));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(net587),
    .X(net855));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(net18),
    .X(net856));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(net259),
    .X(net857));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(net657),
    .X(net858));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(net47),
    .X(net859));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(net566),
    .X(net860));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(net415),
    .X(net861));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(net39),
    .X(net862));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(net245),
    .X(net863));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(net103),
    .X(net864));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(net291),
    .X(net865));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(net148),
    .X(net866));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(net437),
    .X(net867));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(net294),
    .X(net868));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(net10),
    .X(net869));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(net366),
    .X(net870));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(net350),
    .X(net871));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(net677),
    .X(net872));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(net556),
    .X(net873));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(net137),
    .X(net874));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(net640),
    .X(net875));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(net54),
    .X(net876));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(net384),
    .X(net877));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(net676),
    .X(net878));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(net636),
    .X(net879));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(net115),
    .X(net880));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(net343),
    .X(net881));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(net586),
    .X(net882));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(net341),
    .X(net883));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(net362),
    .X(net884));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(net40),
    .X(net885));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(net213),
    .X(net886));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(net204),
    .X(net887));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(net674),
    .X(net888));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(net243),
    .X(net889));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(net396),
    .X(net890));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(net599),
    .X(net891));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(net298),
    .X(net892));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(net588),
    .X(net893));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(net589),
    .X(net894));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(net264),
    .X(net895));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(net675),
    .X(net896));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(net582),
    .X(net897));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(net442),
    .X(net898));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(net179),
    .X(net899));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(net526),
    .X(net900));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(net606),
    .X(net901));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(net38),
    .X(net902));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(net107),
    .X(net903));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(net511),
    .X(net904));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(net655),
    .X(net905));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(net235),
    .X(net906));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(net273),
    .X(net907));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(net162),
    .X(net908));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(net130),
    .X(net909));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(net584),
    .X(net910));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(net13),
    .X(net911));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(net248),
    .X(net912));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(net361),
    .X(net913));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(net561),
    .X(net914));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(net521),
    .X(net915));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(net188),
    .X(net916));
 sky130_fd_sc_hd__dlygate4sd3_1 hold96 (.A(net659),
    .X(net917));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(net627),
    .X(net918));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(net519),
    .X(net919));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(net803),
    .X(net920));
 sky130_fd_sc_hd__dlygate4sd3_1 hold100 (.A(net169),
    .X(net921));
 sky130_fd_sc_hd__dlygate4sd3_1 hold101 (.A(net557),
    .X(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_A (.DIODE(clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(in0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(in1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(in10));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(in11));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(in12));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(in13));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(in14));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(in15));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(in16));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(in17));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(in18));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(in19));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(in2));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(in20));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(in21));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(in22));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(in23));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(in24));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(in25));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(in26));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(in27));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_A (.DIODE(in28));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_A (.DIODE(in29));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_A (.DIODE(in3));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_A (.DIODE(in30));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_A (.DIODE(in31));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_A (.DIODE(in32));
 sky130_fd_sc_hd__diode_2 ANTENNA_input28_A (.DIODE(in33));
 sky130_fd_sc_hd__diode_2 ANTENNA_input29_A (.DIODE(in34));
 sky130_fd_sc_hd__diode_2 ANTENNA_input30_A (.DIODE(in35));
 sky130_fd_sc_hd__diode_2 ANTENNA_input31_A (.DIODE(in36));
 sky130_fd_sc_hd__diode_2 ANTENNA_input32_A (.DIODE(in37));
 sky130_fd_sc_hd__diode_2 ANTENNA_input33_A (.DIODE(in38));
 sky130_fd_sc_hd__diode_2 ANTENNA_input34_A (.DIODE(in39));
 sky130_fd_sc_hd__diode_2 ANTENNA_input35_A (.DIODE(in4));
 sky130_fd_sc_hd__diode_2 ANTENNA_input36_A (.DIODE(in40));
 sky130_fd_sc_hd__diode_2 ANTENNA_input37_A (.DIODE(in41));
 sky130_fd_sc_hd__diode_2 ANTENNA_input38_A (.DIODE(in42));
 sky130_fd_sc_hd__diode_2 ANTENNA_input39_A (.DIODE(in43));
 sky130_fd_sc_hd__diode_2 ANTENNA_input40_A (.DIODE(in44));
 sky130_fd_sc_hd__diode_2 ANTENNA_input41_A (.DIODE(in45));
 sky130_fd_sc_hd__diode_2 ANTENNA_input42_A (.DIODE(in46));
 sky130_fd_sc_hd__diode_2 ANTENNA_input43_A (.DIODE(in47));
 sky130_fd_sc_hd__diode_2 ANTENNA_input44_A (.DIODE(in48));
 sky130_fd_sc_hd__diode_2 ANTENNA_input45_A (.DIODE(in49));
 sky130_fd_sc_hd__diode_2 ANTENNA_input46_A (.DIODE(in5));
 sky130_fd_sc_hd__diode_2 ANTENNA_input47_A (.DIODE(in50));
 sky130_fd_sc_hd__diode_2 ANTENNA_input48_A (.DIODE(in51));
 sky130_fd_sc_hd__diode_2 ANTENNA_input49_A (.DIODE(in52));
 sky130_fd_sc_hd__diode_2 ANTENNA_input50_A (.DIODE(in53));
 sky130_fd_sc_hd__diode_2 ANTENNA_input51_A (.DIODE(in54));
 sky130_fd_sc_hd__diode_2 ANTENNA_input52_A (.DIODE(in55));
 sky130_fd_sc_hd__diode_2 ANTENNA_input53_A (.DIODE(in56));
 sky130_fd_sc_hd__diode_2 ANTENNA_input54_A (.DIODE(in57));
 sky130_fd_sc_hd__diode_2 ANTENNA_input55_A (.DIODE(in58));
 sky130_fd_sc_hd__diode_2 ANTENNA_input56_A (.DIODE(in59));
 sky130_fd_sc_hd__diode_2 ANTENNA_input57_A (.DIODE(in6));
 sky130_fd_sc_hd__diode_2 ANTENNA_input58_A (.DIODE(in60));
 sky130_fd_sc_hd__diode_2 ANTENNA_input59_A (.DIODE(in61));
 sky130_fd_sc_hd__diode_2 ANTENNA_input60_A (.DIODE(in62));
 sky130_fd_sc_hd__diode_2 ANTENNA_input61_A (.DIODE(in63));
 sky130_fd_sc_hd__diode_2 ANTENNA_input62_A (.DIODE(in64));
 sky130_fd_sc_hd__diode_2 ANTENNA_input63_A (.DIODE(in65));
 sky130_fd_sc_hd__diode_2 ANTENNA_input64_A (.DIODE(in66));
 sky130_fd_sc_hd__diode_2 ANTENNA_input65_A (.DIODE(in67));
 sky130_fd_sc_hd__diode_2 ANTENNA_input66_A (.DIODE(in68));
 sky130_fd_sc_hd__diode_2 ANTENNA_input67_A (.DIODE(in69));
 sky130_fd_sc_hd__diode_2 ANTENNA_input68_A (.DIODE(in7));
 sky130_fd_sc_hd__diode_2 ANTENNA_input69_A (.DIODE(in70));
 sky130_fd_sc_hd__diode_2 ANTENNA_input70_A (.DIODE(in71));
 sky130_fd_sc_hd__diode_2 ANTENNA_input71_A (.DIODE(in72));
 sky130_fd_sc_hd__diode_2 ANTENNA_input72_A (.DIODE(in74));
 sky130_fd_sc_hd__diode_2 ANTENNA_input73_A (.DIODE(in75));
 sky130_fd_sc_hd__diode_2 ANTENNA_input74_A (.DIODE(in76));
 sky130_fd_sc_hd__diode_2 ANTENNA_input75_A (.DIODE(in77));
 sky130_fd_sc_hd__diode_2 ANTENNA_input76_A (.DIODE(in78));
 sky130_fd_sc_hd__diode_2 ANTENNA_input77_A (.DIODE(in79));
 sky130_fd_sc_hd__diode_2 ANTENNA_input78_A (.DIODE(in8));
 sky130_fd_sc_hd__diode_2 ANTENNA_input79_A (.DIODE(in80));
 sky130_fd_sc_hd__diode_2 ANTENNA_input80_A (.DIODE(in81));
 sky130_fd_sc_hd__diode_2 ANTENNA_input81_A (.DIODE(in82));
 sky130_fd_sc_hd__diode_2 ANTENNA_input82_A (.DIODE(in83));
 sky130_fd_sc_hd__diode_2 ANTENNA_input83_A (.DIODE(in84));
 sky130_fd_sc_hd__diode_2 ANTENNA_input84_A (.DIODE(in85));
 sky130_fd_sc_hd__diode_2 ANTENNA_input85_A (.DIODE(in86));
 sky130_fd_sc_hd__diode_2 ANTENNA_input86_A (.DIODE(in87));
 sky130_fd_sc_hd__diode_2 ANTENNA_input87_A (.DIODE(in88));
 sky130_fd_sc_hd__diode_2 ANTENNA_input88_A (.DIODE(in89));
 sky130_fd_sc_hd__diode_2 ANTENNA_input89_A (.DIODE(in9));
 sky130_fd_sc_hd__diode_2 ANTENNA_input90_A (.DIODE(in90));
 sky130_fd_sc_hd__diode_2 ANTENNA_input91_A (.DIODE(in91));
 sky130_fd_sc_hd__diode_2 ANTENNA_input92_A (.DIODE(in92));
 sky130_fd_sc_hd__diode_2 ANTENNA_input93_A (.DIODE(in93));
 sky130_fd_sc_hd__diode_2 ANTENNA_input94_A (.DIODE(in94));
 sky130_fd_sc_hd__diode_2 ANTENNA_input95_A (.DIODE(in95));
 sky130_fd_sc_hd__diode_2 ANTENNA_input96_A (.DIODE(in96));
 sky130_fd_sc_hd__diode_2 ANTENNA_input97_A (.DIODE(in97));
 sky130_fd_sc_hd__diode_2 ANTENNA_input98_A (.DIODE(in98));
 sky130_fd_sc_hd__diode_2 ANTENNA_input99_A (.DIODE(in99));
 sky130_fd_sc_hd__diode_2 ANTENNA_s770_D (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_X (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_A0 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_SET_B (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_c180_A2 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_X (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_X (.DIODE(net592));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_RESET_B (.DIODE(net592));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_X (.DIODE(net604));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_RESET_B (.DIODE(net604));
 sky130_fd_sc_hd__diode_2 ANTENNA_input45_X (.DIODE(net735));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_S0 (.DIODE(net735));
 sky130_fd_sc_hd__diode_2 ANTENNA_input49_X (.DIODE(net739));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_B (.DIODE(net739));
 sky130_fd_sc_hd__diode_2 ANTENNA_input63_X (.DIODE(net753));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge753_SCD (.DIODE(net753));
 sky130_fd_sc_hd__diode_2 ANTENNA_output102_A (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_s789_Q (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge744_SCE (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_S0 (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_S1 (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_output104_A (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_D (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_SCE (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_SCE (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_Q (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_output109_A (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_s788_Q_N (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_A3 (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_S0 (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold99_A (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA_output113_A (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_B (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_SCD (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_SCD (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA_c344_D1 (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_Q (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA_output117_A (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge733_RESET_B (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_c125_RESET_B (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_c122_A (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_c121_X (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_output118_A (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_A (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_B (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c222_Q (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_output121_A (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_A (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_c103_X (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_output123_A (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_D (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c229_D1 (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c228_Q (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_3__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_2__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_1__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_0__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_X (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_35_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_34_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_33_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_31_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_3_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_2_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_1_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_0_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_0__f_clk_X (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_13_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_12_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_11_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_10_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_9_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_8_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_7_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_6_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_5_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_4_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_1__f_clk_X (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_32_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_29_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_28_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_27_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_26_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_25_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_24_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_23_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_22_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_20_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_2__f_clk_X (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_30_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_21_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_19_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_18_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_17_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_16_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_15_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_14_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_3__f_clk_X (.DIODE(clknet_2_3__leaf_clk));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_396 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_506 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_357 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_270 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_303 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_476 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_488 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_607 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_8 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_594 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_606 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_624 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_8 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_368 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_20 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_539 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_560 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_619 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_359 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_20 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_584 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_623 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_8 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_553 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_247 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_14 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_480 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_618 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_16 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_8 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_527 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_476 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_510 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_506 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_609 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_581 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_228 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_553 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_367 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_312 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_310 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_60 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_62 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_172 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_115 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_86 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_282 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_8 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_8 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_8 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_617 ();
endmodule
