module netlist_1 (clk,
    in0,
    in1,
    in10,
    in11,
    in12,
    in13,
    in14,
    in15,
    in16,
    in17,
    in18,
    in19,
    in2,
    in20,
    in21,
    in22,
    in23,
    in24,
    in25,
    in26,
    in27,
    in28,
    in29,
    in3,
    in30,
    in31,
    in32,
    in33,
    in34,
    in35,
    in36,
    in37,
    in38,
    in39,
    in4,
    in40,
    in41,
    in42,
    in43,
    in44,
    in45,
    in46,
    in47,
    in48,
    in49,
    in5,
    in50,
    in51,
    in52,
    in53,
    in54,
    in55,
    in56,
    in57,
    in58,
    in59,
    in6,
    in60,
    in61,
    in7,
    in8,
    in9,
    out0,
    out1,
    out10,
    out11,
    out12,
    out13,
    out14,
    out15,
    out16,
    out17,
    out18,
    out19,
    out2,
    out20,
    out21,
    out22,
    out23,
    out24,
    out25,
    out26,
    out27,
    out28,
    out29,
    out3,
    out30,
    out31,
    out32,
    out33,
    out34,
    out35,
    out36,
    out37,
    out38,
    out39,
    out4,
    out40,
    out41,
    out42,
    out43,
    out44,
    out45,
    out46,
    out47,
    out48,
    out49,
    out5,
    out50,
    out51,
    out52,
    out53,
    out54,
    out55,
    out56,
    out57,
    out58,
    out59,
    out6,
    out60,
    out61,
    out7,
    out8,
    out9,
    rst);
 input clk;
 input in0;
 input in1;
 input in10;
 input in11;
 input in12;
 input in13;
 input in14;
 input in15;
 input in16;
 input in17;
 input in18;
 input in19;
 input in2;
 input in20;
 input in21;
 input in22;
 input in23;
 input in24;
 input in25;
 input in26;
 input in27;
 input in28;
 input in29;
 input in3;
 input in30;
 input in31;
 input in32;
 input in33;
 input in34;
 input in35;
 input in36;
 input in37;
 input in38;
 input in39;
 input in4;
 input in40;
 input in41;
 input in42;
 input in43;
 input in44;
 input in45;
 input in46;
 input in47;
 input in48;
 input in49;
 input in5;
 input in50;
 input in51;
 input in52;
 input in53;
 input in54;
 input in55;
 input in56;
 input in57;
 input in58;
 input in59;
 input in6;
 input in60;
 input in61;
 input in7;
 input in8;
 input in9;
 output out0;
 output out1;
 output out10;
 output out11;
 output out12;
 output out13;
 output out14;
 output out15;
 output out16;
 output out17;
 output out18;
 output out19;
 output out2;
 output out20;
 output out21;
 output out22;
 output out23;
 output out24;
 output out25;
 output out26;
 output out27;
 output out28;
 output out29;
 output out3;
 output out30;
 output out31;
 output out32;
 output out33;
 output out34;
 output out35;
 output out36;
 output out37;
 output out38;
 output out39;
 output out4;
 output out40;
 output out41;
 output out42;
 output out43;
 output out44;
 output out45;
 output out46;
 output out47;
 output out48;
 output out49;
 output out5;
 output out50;
 output out51;
 output out52;
 output out53;
 output out54;
 output out55;
 output out56;
 output out57;
 output out58;
 output out59;
 output out6;
 output out60;
 output out61;
 output out7;
 output out8;
 output out9;
 input rst;

 wire net0;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net63;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net64;
 wire net640;
 wire net641;
 wire net642;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net65;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net66;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net67;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net68;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net69;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net7;
 wire net70;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net71;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net72;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net73;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net74;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net75;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net76;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net77;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net78;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net79;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net8;
 wire net80;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net81;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net82;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net83;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net643;
 wire net675;
 wire net699;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_0_net827;
 wire clknet_1_0__leaf_net827;
 wire clknet_1_1__leaf_net827;
 wire clknet_0_net597;
 wire clknet_1_0__leaf_net597;
 wire clknet_1_1__leaf_net597;
 wire clknet_0_net621;
 wire clknet_1_0__leaf_net621;
 wire clknet_1_1__leaf_net621;
 wire clknet_0_net644;
 wire clknet_1_0__leaf_net644;
 wire clknet_1_1__leaf_net644;
 wire clknet_0_net646;
 wire clknet_1_0__leaf_net646;
 wire clknet_1_1__leaf_net646;
 wire clknet_0_net826;
 wire clknet_1_0__leaf_net826;
 wire clknet_1_1__leaf_net826;
 wire clknet_0_net654;
 wire clknet_1_0__leaf_net654;
 wire clknet_1_1__leaf_net654;
 wire clknet_0_net653;
 wire clknet_1_0__leaf_net653;
 wire clknet_1_1__leaf_net653;
 wire clknet_0_net645;
 wire clknet_1_0__leaf_net645;
 wire clknet_1_1__leaf_net645;
 wire clknet_0_net655;
 wire clknet_1_0__leaf_net655;
 wire clknet_1_1__leaf_net655;
 wire clknet_0_net651;
 wire clknet_1_0__leaf_net651;
 wire clknet_1_1__leaf_net651;
 wire clknet_0_net625;
 wire clknet_1_0__leaf_net625;
 wire clknet_1_1__leaf_net625;
 wire clknet_0_net636;
 wire clknet_1_0__leaf_net636;
 wire clknet_1_1__leaf_net636;
 wire clknet_0_net623;
 wire clknet_1_0__leaf_net623;
 wire clknet_1_1__leaf_net623;
 wire clknet_0_net633;
 wire clknet_1_0__leaf_net633;
 wire clknet_1_1__leaf_net633;
 wire clknet_0_net629;
 wire clknet_1_0__leaf_net629;
 wire clknet_1_1__leaf_net629;
 wire clknet_0_net635;
 wire clknet_1_0__leaf_net635;
 wire clknet_1_1__leaf_net635;
 wire clknet_0_net634;
 wire clknet_1_0__leaf_net634;
 wire clknet_1_1__leaf_net634;
 wire clknet_0_net632;
 wire clknet_1_0__leaf_net632;
 wire clknet_1_1__leaf_net632;
 wire clknet_0_net631;
 wire clknet_1_0__leaf_net631;
 wire clknet_1_1__leaf_net631;
 wire clknet_0_net630;
 wire clknet_1_0__leaf_net630;
 wire clknet_1_1__leaf_net630;
 wire clknet_0_net626;
 wire clknet_1_0__leaf_net626;
 wire clknet_1_1__leaf_net626;
 wire clknet_0_net624;
 wire clknet_1_0__leaf_net624;
 wire clknet_1_1__leaf_net624;
 wire clknet_0_net622;
 wire clknet_1_0__leaf_net622;
 wire clknet_1_1__leaf_net622;
 wire clknet_0_net607;
 wire clknet_1_0__leaf_net607;
 wire clknet_1_1__leaf_net607;
 wire clknet_0_net609;
 wire clknet_1_0__leaf_net609;
 wire clknet_1_1__leaf_net609;
 wire clknet_0_net608;
 wire clknet_1_0__leaf_net608;
 wire clknet_1_1__leaf_net608;
 wire clknet_0_net600;
 wire clknet_1_0__leaf_net600;
 wire clknet_1_1__leaf_net600;
 wire clknet_0_net603;
 wire clknet_1_0__leaf_net603;
 wire clknet_1_1__leaf_net603;
 wire clknet_0_net604;
 wire clknet_1_0__leaf_net604;
 wire clknet_1_1__leaf_net604;
 wire clknet_0_net606;
 wire clknet_1_0__leaf_net606;
 wire clknet_1_1__leaf_net606;
 wire clknet_0_net468;
 wire clknet_1_0__leaf_net468;
 wire clknet_1_1__leaf_net468;
 wire clknet_0_net825;
 wire clknet_1_0__leaf_net825;
 wire clknet_1_1__leaf_net825;
 wire clknet_0_net238;
 wire clknet_1_0__leaf_net238;
 wire clknet_1_1__leaf_net238;
 wire clknet_0_net251;
 wire clknet_1_0__leaf_net251;
 wire clknet_1_1__leaf_net251;
 wire clknet_0_net239;
 wire clknet_1_0__leaf_net239;
 wire clknet_1_1__leaf_net239;
 wire clknet_0_net808;
 wire clknet_1_0__leaf_net808;
 wire clknet_1_1__leaf_net808;
 wire clknet_0_net541;
 wire clknet_1_0__leaf_net541;
 wire clknet_1_1__leaf_net541;
 wire clknet_0_net807;
 wire clknet_1_0__leaf_net807;
 wire clknet_1_1__leaf_net807;
 wire clknet_0_net806;
 wire clknet_1_0__leaf_net806;
 wire clknet_1_1__leaf_net806;
 wire clknet_0_net528;
 wire clknet_1_0__leaf_net528;
 wire clknet_1_1__leaf_net528;
 wire clknet_0_net788;
 wire clknet_1_0__leaf_net788;
 wire clknet_1_1__leaf_net788;
 wire clknet_0_net549;
 wire clknet_1_0__leaf_net549;
 wire clknet_1_1__leaf_net549;
 wire clknet_0_net567;
 wire clknet_1_0__leaf_net567;
 wire clknet_1_1__leaf_net567;
 wire clknet_0_net555;
 wire clknet_1_0__leaf_net555;
 wire clknet_1_1__leaf_net555;
 wire clknet_0_net563;
 wire clknet_1_0__leaf_net563;
 wire clknet_1_1__leaf_net563;
 wire clknet_0_net562;
 wire clknet_1_0__leaf_net562;
 wire clknet_1_1__leaf_net562;
 wire clknet_0_net566;
 wire clknet_1_0__leaf_net566;
 wire clknet_1_1__leaf_net566;
 wire clknet_0_net556;
 wire clknet_1_0__leaf_net556;
 wire clknet_1_1__leaf_net556;
 wire clknet_0_net560;
 wire clknet_1_0__leaf_net560;
 wire clknet_1_1__leaf_net560;
 wire clknet_0_net559;
 wire clknet_1_0__leaf_net559;
 wire clknet_1_1__leaf_net559;
 wire clknet_0_net557;
 wire clknet_1_0__leaf_net557;
 wire clknet_1_1__leaf_net557;
 wire clknet_0_net558;
 wire clknet_1_0__leaf_net558;
 wire clknet_1_1__leaf_net558;
 wire clknet_0_net561;
 wire clknet_1_0__leaf_net561;
 wire clknet_1_1__leaf_net561;
 wire clknet_0_net552;
 wire clknet_1_0__leaf_net552;
 wire clknet_1_1__leaf_net552;
 wire clknet_0_net554;
 wire clknet_1_0__leaf_net554;
 wire clknet_1_1__leaf_net554;
 wire clknet_0_net551;
 wire clknet_1_0__leaf_net551;
 wire clknet_1_1__leaf_net551;
 wire clknet_0_net550;
 wire clknet_1_0__leaf_net550;
 wire clknet_1_1__leaf_net550;
 wire clknet_0_net553;
 wire clknet_1_0__leaf_net553;
 wire clknet_1_1__leaf_net553;
 wire clknet_0_net439;
 wire clknet_1_0__leaf_net439;
 wire clknet_1_1__leaf_net439;
 wire clknet_0_net449;
 wire clknet_1_0__leaf_net449;
 wire clknet_1_1__leaf_net449;
 wire clknet_0_net450;
 wire clknet_1_0__leaf_net450;
 wire clknet_1_1__leaf_net450;
 wire clknet_0_net446;
 wire clknet_1_0__leaf_net446;
 wire clknet_1_1__leaf_net446;
 wire clknet_0_net444;
 wire clknet_1_0__leaf_net444;
 wire clknet_1_1__leaf_net444;
 wire clknet_0_net445;
 wire clknet_1_0__leaf_net445;
 wire clknet_1_1__leaf_net445;
 wire clknet_0_net447;
 wire clknet_1_0__leaf_net447;
 wire clknet_1_1__leaf_net447;
 wire clknet_0_net442;
 wire clknet_1_0__leaf_net442;
 wire clknet_1_1__leaf_net442;
 wire clknet_0_net443;
 wire clknet_1_0__leaf_net443;
 wire clknet_1_1__leaf_net443;
 wire clknet_0_net441;
 wire clknet_1_0__leaf_net441;
 wire clknet_1_1__leaf_net441;
 wire clknet_0_net440;
 wire clknet_1_0__leaf_net440;
 wire clknet_1_1__leaf_net440;
 wire clknet_0_net434;
 wire clknet_1_0__leaf_net434;
 wire clknet_1_1__leaf_net434;
 wire clknet_0_net436;
 wire clknet_1_0__leaf_net436;
 wire clknet_1_1__leaf_net436;
 wire clknet_0_net437;
 wire clknet_1_0__leaf_net437;
 wire clknet_1_1__leaf_net437;
 wire clknet_0_net438;
 wire clknet_1_0__leaf_net438;
 wire clknet_1_1__leaf_net438;
 wire clknet_0_net435;
 wire clknet_1_0__leaf_net435;
 wire clknet_1_1__leaf_net435;
 wire clknet_0_net346;
 wire clknet_1_0__leaf_net346;
 wire clknet_1_1__leaf_net346;
 wire clknet_0_net360;
 wire clknet_1_0__leaf_net360;
 wire clknet_1_1__leaf_net360;
 wire clknet_0_net363;
 wire clknet_1_0__leaf_net363;
 wire clknet_1_1__leaf_net363;
 wire clknet_0_net362;
 wire clknet_1_0__leaf_net362;
 wire clknet_1_1__leaf_net362;
 wire clknet_0_net361;
 wire clknet_1_0__leaf_net361;
 wire clknet_1_1__leaf_net361;
 wire clknet_0_net359;
 wire clknet_1_0__leaf_net359;
 wire clknet_1_1__leaf_net359;
 wire clknet_0_net572;
 wire clknet_1_0__leaf_net572;
 wire clknet_1_1__leaf_net572;
 wire clknet_0_net589;
 wire clknet_1_0__leaf_net589;
 wire clknet_1_1__leaf_net589;
 wire clknet_0_net591;
 wire clknet_1_0__leaf_net591;
 wire clknet_1_1__leaf_net591;
 wire clknet_0_net590;
 wire clknet_1_0__leaf_net590;
 wire clknet_1_1__leaf_net590;
 wire clknet_0_net576;
 wire clknet_1_0__leaf_net576;
 wire clknet_1_1__leaf_net576;
 wire clknet_0_net575;
 wire clknet_1_0__leaf_net575;
 wire clknet_1_1__leaf_net575;
 wire clknet_0_net574;
 wire clknet_1_0__leaf_net574;
 wire clknet_1_1__leaf_net574;
 wire clknet_0_net573;
 wire clknet_1_0__leaf_net573;
 wire clknet_1_1__leaf_net573;
 wire clknet_0_net460;
 wire clknet_1_0__leaf_net460;
 wire clknet_1_1__leaf_net460;
 wire clknet_0_net467;
 wire clknet_1_0__leaf_net467;
 wire clknet_1_1__leaf_net467;
 wire clknet_0_net463;
 wire clknet_1_0__leaf_net463;
 wire clknet_1_1__leaf_net463;
 wire clknet_0_net461;
 wire clknet_1_0__leaf_net461;
 wire clknet_1_1__leaf_net461;
 wire clknet_0_net462;
 wire clknet_1_0__leaf_net462;
 wire clknet_1_1__leaf_net462;
 wire clknet_0_net371;
 wire clknet_1_0__leaf_net371;
 wire clknet_1_1__leaf_net371;
 wire clknet_0_net380;
 wire clknet_1_0__leaf_net380;
 wire clknet_1_1__leaf_net380;
 wire clknet_0_net375;
 wire clknet_1_0__leaf_net375;
 wire clknet_1_1__leaf_net375;
 wire clknet_0_net373;
 wire clknet_1_0__leaf_net373;
 wire clknet_1_1__leaf_net373;
 wire clknet_0_net736;
 wire clknet_1_0__leaf_net736;
 wire clknet_1_1__leaf_net736;
 wire clknet_0_net668;
 wire clknet_1_0__leaf_net668;
 wire clknet_1_1__leaf_net668;
 wire clknet_0_net396;
 wire clknet_1_0__leaf_net396;
 wire clknet_1_1__leaf_net396;
 wire clknet_0_net403;
 wire clknet_1_0__leaf_net403;
 wire clknet_1_1__leaf_net403;
 wire clknet_0_net406;
 wire clknet_1_0__leaf_net406;
 wire clknet_1_1__leaf_net406;
 wire clknet_0_net411;
 wire clknet_1_0__leaf_net411;
 wire clknet_1_1__leaf_net411;
 wire clknet_0_net412;
 wire clknet_1_0__leaf_net412;
 wire clknet_1_1__leaf_net412;
 wire clknet_0_net410;
 wire clknet_1_0__leaf_net410;
 wire clknet_1_1__leaf_net410;
 wire clknet_0_net415;
 wire clknet_1_0__leaf_net415;
 wire clknet_1_1__leaf_net415;
 wire clknet_0_net408;
 wire clknet_1_0__leaf_net408;
 wire clknet_1_1__leaf_net408;
 wire clknet_0_net407;
 wire clknet_1_0__leaf_net407;
 wire clknet_1_1__leaf_net407;
 wire clknet_0_net401;
 wire clknet_1_0__leaf_net401;
 wire clknet_1_1__leaf_net401;
 wire clknet_0_net430;
 wire clknet_1_0__leaf_net430;
 wire clknet_1_1__leaf_net430;
 wire clknet_0_net404;
 wire clknet_1_0__leaf_net404;
 wire clknet_1_1__leaf_net404;
 wire clknet_0_net402;
 wire clknet_1_0__leaf_net402;
 wire clknet_1_1__leaf_net402;
 wire clknet_0_net400;
 wire clknet_1_0__leaf_net400;
 wire clknet_1_1__leaf_net400;
 wire clknet_0_net399;
 wire clknet_1_0__leaf_net399;
 wire clknet_1_1__leaf_net399;
 wire clknet_0_net398;
 wire clknet_1_0__leaf_net398;
 wire clknet_1_1__leaf_net398;
 wire clknet_0_net397;
 wire clknet_1_0__leaf_net397;
 wire clknet_1_1__leaf_net397;
 wire clknet_0_net394;
 wire clknet_1_0__leaf_net394;
 wire clknet_1_1__leaf_net394;
 wire clknet_0_net395;
 wire clknet_1_0__leaf_net395;
 wire clknet_1_1__leaf_net395;
 wire clknet_0_net299;
 wire clknet_1_0__leaf_net299;
 wire clknet_1_1__leaf_net299;
 wire clknet_0_net288;
 wire clknet_1_0__leaf_net288;
 wire clknet_1_1__leaf_net288;
 wire clknet_0_net297;
 wire clknet_1_0__leaf_net297;
 wire clknet_1_1__leaf_net297;
 wire clknet_0_net296;
 wire clknet_1_0__leaf_net296;
 wire clknet_1_1__leaf_net296;
 wire clknet_0_net294;
 wire clknet_1_0__leaf_net294;
 wire clknet_1_1__leaf_net294;
 wire clknet_0_net292;
 wire clknet_1_0__leaf_net292;
 wire clknet_1_1__leaf_net292;
 wire clknet_0_net295;
 wire clknet_1_0__leaf_net295;
 wire clknet_1_1__leaf_net295;
 wire clknet_0_net291;
 wire clknet_1_0__leaf_net291;
 wire clknet_1_1__leaf_net291;
 wire clknet_0_net289;
 wire clknet_1_0__leaf_net289;
 wire clknet_1_1__leaf_net289;
 wire clknet_0_net290;
 wire clknet_1_0__leaf_net290;
 wire clknet_1_1__leaf_net290;
 wire clknet_0_net910;
 wire clknet_1_0__leaf_net910;
 wire clknet_1_1__leaf_net910;
 wire clknet_0_net311;
 wire clknet_1_0__leaf_net311;
 wire clknet_1_1__leaf_net311;
 wire clknet_0_net305;
 wire clknet_1_0__leaf_net305;
 wire clknet_1_1__leaf_net305;
 wire clknet_0_net306;
 wire clknet_1_0__leaf_net306;
 wire clknet_1_1__leaf_net306;
 wire clknet_0_net312;
 wire clknet_1_0__leaf_net312;
 wire clknet_1_1__leaf_net312;
 wire clknet_0_net308;
 wire clknet_1_0__leaf_net308;
 wire clknet_1_1__leaf_net308;
 wire clknet_0_net314;
 wire clknet_1_0__leaf_net314;
 wire clknet_1_1__leaf_net314;
 wire clknet_0_net317;
 wire clknet_1_0__leaf_net317;
 wire clknet_1_1__leaf_net317;
 wire clknet_0_net303;
 wire clknet_1_0__leaf_net303;
 wire clknet_1_1__leaf_net303;
 wire clknet_0_net310;
 wire clknet_1_0__leaf_net310;
 wire clknet_1_1__leaf_net310;
 wire clknet_0_net307;
 wire clknet_1_0__leaf_net307;
 wire clknet_1_1__leaf_net307;
 wire clknet_0_net372;
 wire clknet_1_0__leaf_net372;
 wire clknet_1_1__leaf_net372;
 wire clknet_0_net386;
 wire clknet_1_0__leaf_net386;
 wire clknet_1_1__leaf_net386;
 wire clknet_0_net367;
 wire clknet_1_0__leaf_net367;
 wire clknet_1_1__leaf_net367;
 wire clknet_0_net381;
 wire clknet_1_0__leaf_net381;
 wire clknet_1_1__leaf_net381;
 wire clknet_0_net358;
 wire clknet_1_0__leaf_net358;
 wire clknet_1_1__leaf_net358;
 wire clknet_0_net357;
 wire clknet_1_0__leaf_net357;
 wire clknet_1_1__leaf_net357;
 wire clknet_0_net352;
 wire clknet_1_0__leaf_net352;
 wire clknet_1_1__leaf_net352;
 wire clknet_0_net351;
 wire clknet_1_0__leaf_net351;
 wire clknet_1_1__leaf_net351;
 wire clknet_0_net350;
 wire clknet_1_0__leaf_net350;
 wire clknet_1_1__leaf_net350;
 wire clknet_0_net354;
 wire clknet_1_0__leaf_net354;
 wire clknet_1_1__leaf_net354;
 wire clknet_0_net356;
 wire clknet_1_0__leaf_net356;
 wire clknet_1_1__leaf_net356;
 wire clknet_0_net353;
 wire clknet_1_0__leaf_net353;
 wire clknet_1_1__leaf_net353;
 wire clknet_0_net355;
 wire clknet_1_0__leaf_net355;
 wire clknet_1_1__leaf_net355;
 wire clknet_0_net349;
 wire clknet_1_0__leaf_net349;
 wire clknet_1_1__leaf_net349;
 wire clknet_0_net368;
 wire clknet_1_0__leaf_net368;
 wire clknet_1_1__leaf_net368;
 wire clknet_0_net376;
 wire clknet_1_0__leaf_net376;
 wire clknet_1_1__leaf_net376;
 wire clknet_0_net347;
 wire clknet_1_0__leaf_net347;
 wire clknet_1_1__leaf_net347;
 wire clknet_0_net787;
 wire clknet_1_0__leaf_net787;
 wire clknet_1_1__leaf_net787;
 wire clknet_0_net342;
 wire clknet_1_0__leaf_net342;
 wire clknet_1_1__leaf_net342;
 wire clknet_0_net786;
 wire clknet_1_0__leaf_net786;
 wire clknet_1_1__leaf_net786;
 wire clknet_0_net341;
 wire clknet_1_0__leaf_net341;
 wire clknet_1_1__leaf_net341;
 wire clknet_0_net769;
 wire clknet_1_0__leaf_net769;
 wire clknet_1_1__leaf_net769;
 wire clknet_0_net302;
 wire clknet_1_0__leaf_net302;
 wire clknet_1_1__leaf_net302;
 wire clknet_0_net737;
 wire clknet_1_0__leaf_net737;
 wire clknet_1_1__leaf_net737;
 wire clknet_0_net169;
 wire clknet_1_0__leaf_net169;
 wire clknet_1_1__leaf_net169;
 wire clknet_0_net176;
 wire clknet_1_0__leaf_net176;
 wire clknet_1_1__leaf_net176;
 wire clknet_0_net192;
 wire clknet_1_0__leaf_net192;
 wire clknet_1_1__leaf_net192;
 wire clknet_0_net166;
 wire clknet_1_0__leaf_net166;
 wire clknet_1_1__leaf_net166;
 wire clknet_0_net175;
 wire clknet_1_0__leaf_net175;
 wire clknet_1_1__leaf_net175;
 wire clknet_0_net180;
 wire clknet_1_0__leaf_net180;
 wire clknet_1_1__leaf_net180;
 wire clknet_0_net168;
 wire clknet_1_0__leaf_net168;
 wire clknet_1_1__leaf_net168;
 wire clknet_0_net768;
 wire clknet_1_0__leaf_net768;
 wire clknet_1_1__leaf_net768;
 wire clknet_0_net158;
 wire clknet_1_0__leaf_net158;
 wire clknet_1_1__leaf_net158;
 wire clknet_0_net157;
 wire clknet_1_0__leaf_net157;
 wire clknet_1_1__leaf_net157;
 wire clknet_0_net767;
 wire clknet_1_0__leaf_net767;
 wire clknet_1_1__leaf_net767;
 wire clknet_0_net256;
 wire clknet_1_0__leaf_net256;
 wire clknet_1_1__leaf_net256;
 wire clknet_0_net270;
 wire clknet_1_0__leaf_net270;
 wire clknet_1_1__leaf_net270;
 wire clknet_0_net257;
 wire clknet_1_0__leaf_net257;
 wire clknet_1_1__leaf_net257;
 wire clknet_0_net134;
 wire clknet_1_0__leaf_net134;
 wire clknet_1_1__leaf_net134;
 wire clknet_0_net133;
 wire clknet_1_0__leaf_net133;
 wire clknet_1_1__leaf_net133;
 wire clknet_0_net735;
 wire clknet_1_0__leaf_net735;
 wire clknet_1_1__leaf_net735;
 wire clknet_0_net118;
 wire clknet_1_0__leaf_net118;
 wire clknet_1_1__leaf_net118;
 wire clknet_0_net119;
 wire clknet_1_0__leaf_net119;
 wire clknet_1_1__leaf_net119;
 wire clknet_0_net117;
 wire clknet_1_0__leaf_net117;
 wire clknet_1_1__leaf_net117;
 wire clknet_0_net128;
 wire clknet_1_0__leaf_net128;
 wire clknet_1_1__leaf_net128;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;

 sky130_fd_sc_hd__and3_1 c100 (.A(net34),
    .B(net36),
    .C(net29),
    .X(net38));
 sky130_fd_sc_hd__and3_1 c101 (.A(net35),
    .B(net27),
    .C(net38),
    .X(net39));
 sky130_fd_sc_hd__or4bb_1 c102 (.A(net31),
    .B(net37),
    .C_N(net36),
    .D_N(net919),
    .X(net40));
 sky130_fd_sc_hd__and3_1 c103 (.A(net40),
    .B(net919),
    .C(net28),
    .X(net41));
 sky130_fd_sc_hd__or4bb_1 c104 (.A(net37),
    .B(net31),
    .C_N(net41),
    .D_N(net28),
    .X(net42));
 sky130_fd_sc_hd__mux4_1 c105 (.A0(net42),
    .A1(net38),
    .A2(net39),
    .A3(net37),
    .S0(net27),
    .S1(net29),
    .X(net43));
 sky130_fd_sc_hd__mux4_1 c106 (.A0(net32),
    .A1(net42),
    .A2(net38),
    .A3(net30),
    .S0(net40),
    .S1(net761),
    .X(net44));
 sky130_fd_sc_hd__mux4_1 c107 (.A0(net39),
    .A1(net41),
    .A2(net42),
    .A3(net27),
    .S0(net36),
    .S1(net761),
    .X(net45));
 sky130_fd_sc_hd__a2111o_1 c108 (.A1(net30),
    .A2(net27),
    .B1(net35),
    .C1(clknet_1_1__leaf_net735),
    .D1(net760),
    .X(net46));
 sky130_fd_sc_hd__mux4_1 c109 (.A0(net38),
    .A1(net46),
    .A2(net31),
    .A3(net42),
    .S0(net37),
    .S1(net760),
    .X(net47));
 sky130_fd_sc_hd__buf_1 c110 (.A(net742),
    .X(net48));
 sky130_fd_sc_hd__and2_0 c111 (.A(net932),
    .B(net741),
    .X(net49));
 sky130_fd_sc_hd__and3_1 c112 (.A(net28),
    .B(net49),
    .C(net932),
    .X(net50));
 sky130_fd_sc_hd__and2_1 c113 (.A(net49),
    .B(net932),
    .X(net51));
 sky130_fd_sc_hd__and2_2 c114 (.A(net930),
    .B(net932),
    .X(net52));
 sky130_fd_sc_hd__and2_0 c115 (.A(net930),
    .B(net932),
    .X(net53));
 sky130_fd_sc_hd__or4bb_2 c116 (.A(net50),
    .B(net53),
    .C_N(net930),
    .D_N(net932),
    .X(net54));
 sky130_fd_sc_hd__or4bb_1 c117 (.A(net49),
    .B(net54),
    .C_N(net52),
    .D_N(net930),
    .X(net55));
 sky130_fd_sc_hd__and3_1 c118 (.A(net55),
    .B(net930),
    .C(net50),
    .X(net56));
 sky130_fd_sc_hd__and3_1 c119 (.A(net52),
    .B(net930),
    .C(net932),
    .X(net57));
 sky130_fd_sc_hd__and3_1 c120 (.A(net54),
    .B(net932),
    .C(net52),
    .X(net58));
 sky130_fd_sc_hd__or4bb_2 c121 (.A(net55),
    .B(net57),
    .C_N(net58),
    .D_N(net930),
    .X(net59));
 sky130_fd_sc_hd__a2111o_1 c122 (.A1(net53),
    .A2(net58),
    .B1(net930),
    .C1(net52),
    .D1(net59),
    .X(net60));
 sky130_fd_sc_hd__or4bb_2 c123 (.A(net48),
    .B(net52),
    .C_N(net57),
    .D_N(net54),
    .X(net61));
 sky130_fd_sc_hd__or4bb_2 c124 (.A(net58),
    .B(net930),
    .C_N(net61),
    .D_N(net54),
    .X(net62));
 sky130_fd_sc_hd__a2111o_1 c125 (.A1(net56),
    .A2(net55),
    .B1(net54),
    .C1(net52),
    .D1(net61),
    .X(net63));
 sky130_fd_sc_hd__mux4_1 c126 (.A0(net54),
    .A1(net56),
    .A2(net61),
    .A3(net63),
    .S0(net932),
    .S1(net52),
    .X(net64));
 sky130_fd_sc_hd__mux4_1 c127 (.A0(net60),
    .A1(net61),
    .A2(net56),
    .A3(net51),
    .S0(net62),
    .S1(net36),
    .X(net65));
 sky130_fd_sc_hd__a2111o_1 c128 (.A1(net57),
    .A2(net63),
    .B1(net60),
    .C1(net62),
    .D1(net48),
    .X(net66));
 sky130_fd_sc_hd__a2111o_1 c129 (.A1(net64),
    .A2(net62),
    .B1(net59),
    .C1(net51),
    .D1(net63),
    .X(net67));
 sky130_fd_sc_hd__a2111o_1 c130 (.A1(net63),
    .A2(net62),
    .B1(net66),
    .C1(net930),
    .D1(net718),
    .X(net68));
 sky130_fd_sc_hd__mux4_1 c131 (.A0(net66),
    .A1(net64),
    .A2(net62),
    .A3(net932),
    .S0(net65),
    .S1(net964),
    .X(net69));
 sky130_fd_sc_hd__and2_1 c132 (.A(net890),
    .B(net887),
    .X(net70));
 sky130_fd_sc_hd__and3_1 c133 (.A(net876),
    .B(net840),
    .C(net845),
    .X(net71));
 sky130_fd_sc_hd__and3_1 c134 (.A(net71),
    .B(net854),
    .C(net843),
    .X(net72));
 sky130_fd_sc_hd__and3_1 c135 (.A(net70),
    .B(net675),
    .C(net699),
    .X(net73));
 sky130_fd_sc_hd__or4bb_4 c136 (.A(net73),
    .B(net838),
    .C_N(net72),
    .D_N(net835),
    .X(net74));
 sky130_fd_sc_hd__or4bb_1 c137 (.A(net71),
    .B(net836),
    .C_N(net72),
    .D_N(net74),
    .X(net75));
 sky130_fd_sc_hd__or4bb_1 c138 (.A(net75),
    .B(net891),
    .C_N(net844),
    .D_N(net74),
    .X(net76));
 sky130_fd_sc_hd__and3_2 c139 (.A(net74),
    .B(net926),
    .C(net841),
    .X(net77));
 sky130_fd_sc_hd__or4bb_2 c140 (.A(net74),
    .B(net77),
    .C_N(net70),
    .D_N(net927),
    .X(net78));
 sky130_fd_sc_hd__a2111o_1 c141 (.A1(net78),
    .A2(net892),
    .B1(net75),
    .C1(net77),
    .D1(net926),
    .X(net79));
 sky130_fd_sc_hd__a2111o_4 c142 (.A1(net79),
    .A2(net74),
    .B1(net77),
    .C1(net78),
    .D1(net926),
    .X(net80));
 sky130_fd_sc_hd__a2111o_1 c143 (.A1(net80),
    .A2(net78),
    .B1(net865),
    .C1(net77),
    .D1(net926),
    .X(net81));
 sky130_fd_sc_hd__mux4_1 c144 (.A0(net77),
    .A1(net837),
    .A2(net80),
    .A3(net81),
    .S0(net926),
    .S1(net74),
    .X(net82));
 sky130_fd_sc_hd__mux4_1 c145 (.A0(net82),
    .A1(net80),
    .A2(net842),
    .A3(net74),
    .S0(net926),
    .S1(net77),
    .X(net83));
 sky130_fd_sc_hd__a2111o_1 c146 (.A1(net71),
    .A2(net77),
    .B1(net74),
    .C1(net80),
    .D1(net927),
    .X(net84));
 sky130_fd_sc_hd__mux4_1 c147 (.A0(net81),
    .A1(net78),
    .A2(net834),
    .A3(net83),
    .S0(net926),
    .S1(net74),
    .X(net85));
 sky130_fd_sc_hd__a2111o_1 c148 (.A1(net85),
    .A2(net80),
    .B1(net82),
    .C1(net74),
    .D1(net926),
    .X(net86));
 sky130_fd_sc_hd__mux4_1 c149 (.A0(net72),
    .A1(net75),
    .A2(net86),
    .A3(net84),
    .S0(net78),
    .S1(net80),
    .X(net87));
 sky130_fd_sc_hd__mux4_1 c150 (.A0(net87),
    .A1(net86),
    .A2(net643),
    .A3(net79),
    .S0(net80),
    .S1(net926),
    .X(net88));
 sky130_fd_sc_hd__mux4_1 c151 (.A0(net83),
    .A1(net82),
    .A2(net86),
    .A3(net80),
    .S0(net926),
    .S1(net763),
    .X(net89));
 sky130_fd_sc_hd__mux4_1 c152 (.A0(net89),
    .A1(net927),
    .A2(net839),
    .A3(net79),
    .S0(net80),
    .S1(net963),
    .X(net90));
 sky130_fd_sc_hd__mux4_1 c153 (.A0(net89),
    .A1(net927),
    .A2(net77),
    .A3(net80),
    .S0(net754),
    .S1(net762),
    .X(net91));
 sky130_fd_sc_hd__and2_1 c154 (.A(net864),
    .B(net848),
    .X(net92));
 sky130_fd_sc_hd__and2_1 c155 (.A(net855),
    .B(net92),
    .X(net93));
 sky130_fd_sc_hd__and2_1 c156 (.A(net93),
    .B(net860),
    .X(net94));
 sky130_fd_sc_hd__and3_1 c157 (.A(net93),
    .B(net867),
    .C(net931),
    .X(net95));
 sky130_fd_sc_hd__or4bb_4 c158 (.A(net931),
    .B(net851),
    .C_N(net856),
    .D_N(net92),
    .X(net96));
 sky130_fd_sc_hd__and3_1 c159 (.A(net73),
    .B(net96),
    .C(net95),
    .X(net97));
 sky130_fd_sc_hd__a2111o_1 c160 (.A1(net859),
    .A2(net93),
    .B1(net97),
    .C1(net931),
    .D1(net92),
    .X(net98));
 sky130_fd_sc_hd__and3_1 c161 (.A(net97),
    .B(net96),
    .C(net93),
    .X(net99));
 sky130_fd_sc_hd__a2111o_2 c162 (.A1(net98),
    .A2(net92),
    .B1(net928),
    .C1(net96),
    .D1(net931),
    .X(net100));
 sky130_fd_sc_hd__and3_2 c163 (.A(net928),
    .B(net862),
    .C(net99),
    .X(net101));
 sky130_fd_sc_hd__a2111o_1 c164 (.A1(net99),
    .A2(net101),
    .B1(net931),
    .C1(net100),
    .D1(net84),
    .X(net102));
 sky130_fd_sc_hd__a2111o_4 c165 (.A1(net101),
    .A2(net846),
    .B1(net96),
    .C1(net931),
    .D1(net102),
    .X(net103));
 sky130_fd_sc_hd__mux4_2 c166 (.A0(net100),
    .A1(net101),
    .A2(net847),
    .A3(net103),
    .S0(net98),
    .S1(net931),
    .X(net104));
 sky130_fd_sc_hd__mux4_2 c167 (.A0(net102),
    .A1(net104),
    .A2(net100),
    .A3(net96),
    .S0(net103),
    .S1(net101),
    .X(net105));
 sky130_fd_sc_hd__mux4_2 c168 (.A0(net105),
    .A1(net96),
    .A2(net104),
    .A3(net850),
    .S0(net103),
    .S1(net101),
    .X(net106));
 sky130_fd_sc_hd__mux4_1 c169 (.A0(net86),
    .A1(net103),
    .A2(net931),
    .A3(net101),
    .S0(net100),
    .S1(net106),
    .X(net107));
 sky130_fd_sc_hd__mux4_2 c170 (.A0(net103),
    .A1(net95),
    .A2(net105),
    .A3(net92),
    .S0(net93),
    .S1(net100),
    .X(net108));
 sky130_fd_sc_hd__mux4_1 c171 (.A0(net92),
    .A1(net103),
    .A2(net108),
    .A3(net101),
    .S0(net105),
    .S1(net104),
    .X(net109));
 sky130_fd_sc_hd__mux4_1 c172 (.A0(net108),
    .A1(net105),
    .A2(net103),
    .A3(net931),
    .S0(net101),
    .X(net110));
 sky130_fd_sc_hd__mux4_1 c173 (.A0(net92),
    .A1(net853),
    .A2(net105),
    .A3(net108),
    .S0(net103),
    .S1(net959),
    .X(net111));
 sky130_fd_sc_hd__mux4_1 c174 (.A0(net95),
    .A1(net108),
    .A2(net931),
    .A3(net103),
    .S0(net713),
    .S1(net961),
    .X(net112));
 sky130_fd_sc_hd__mux4_1 c175 (.A0(net108),
    .A1(net101),
    .A2(net94),
    .A3(net750),
    .S0(net764),
    .S1(net961),
    .X(net113));
 sky130_fd_sc_hd__and2_1 c176 (.A(net104),
    .B(net766),
    .X(net114));
 sky130_fd_sc_hd__and2_1 c177 (.A(net871),
    .B(net114),
    .X(net115));
 sky130_fd_sc_hd__and3_4 c178 (.A(net114),
    .B(net104),
    .C(net766),
    .X(net116));
 sky130_fd_sc_hd__buf_1 c179 (.A(clknet_1_0__leaf_net735),
    .X(net117));
 sky130_fd_sc_hd__buf_1 c180 (.A(clknet_1_0__leaf_net735),
    .X(net118));
 sky130_fd_sc_hd__and3_1 c181 (.A(net114),
    .B(clknet_1_0__leaf_net118),
    .C(net96),
    .X(net119));
 sky130_fd_sc_hd__clkbuf_1 c182 (.A(net828),
    .X(net120));
 sky130_fd_sc_hd__buf_1 c183 (.A(net755),
    .X(net121));
 sky130_fd_sc_hd__buf_1 c184 (.A(net755),
    .X(net122));
 sky130_fd_sc_hd__sdfrbp_1 c185 (.CLK(clknet_4_2_0_clk),
    .D(net121),
    .RESET_B(net115),
    .SCD(net122),
    .SCE(clknet_1_0__leaf_net118),
    .Q(net124),
    .Q_N(net123));
 sky130_fd_sc_hd__sdfrbp_1 c186 (.CLK(clknet_4_0_0_clk),
    .D(net104),
    .RESET_B(net122),
    .SCD(clknet_1_0__leaf_net118),
    .SCE(net106),
    .Q(net126),
    .Q_N(net125));
 sky130_fd_sc_hd__sdfrtn_1 c187 (.CLK_N(clknet_4_2_0_clk),
    .D(clknet_1_1__leaf_net119),
    .RESET_B(net947),
    .SCD(net125),
    .SCE(net121),
    .Q(net127));
 sky130_fd_sc_hd__and3_1 c188 (.A(net126),
    .B(clknet_1_0__leaf_net117),
    .C(net123),
    .X(net128));
 sky130_fd_sc_hd__sdfbbn_1 c189 (.CLK_N(clknet_4_2_0_clk),
    .D(clknet_1_0__leaf_net128),
    .RESET_B(clknet_1_1__leaf_net117),
    .SCD(clknet_1_1__leaf_net118),
    .SCE(clknet_1_0__leaf_net119),
    .SET_B(net116),
    .Q(net130),
    .Q_N(net129));
 sky130_fd_sc_hd__sdfrtp_1 c190 (.CLK(clknet_4_2_0_clk),
    .D(net122),
    .RESET_B(net945),
    .SCD(net127),
    .SCE(net115),
    .Q(net131));
 sky130_fd_sc_hd__mux4_1 c191 (.A0(clknet_1_0__leaf_net117),
    .A1(net131),
    .A2(net124),
    .A3(clknet_1_1__leaf_net118),
    .S0(net125),
    .S1(net116),
    .X(net132));
 sky130_fd_sc_hd__and3_1 c192 (.A(net121),
    .B(net131),
    .C(clknet_1_0__leaf_net767),
    .X(net133));
 sky130_fd_sc_hd__mux4_1 c193 (.A0(net127),
    .A1(net130),
    .A2(clknet_1_1__leaf_net128),
    .A3(clknet_1_1__leaf_net118),
    .S0(clknet_1_1__leaf_net133),
    .S1(clknet_1_1__leaf_net767),
    .X(net134));
 sky130_fd_sc_hd__mux4_1 c194 (.A0(net120),
    .A1(clknet_1_0__leaf_net133),
    .A2(clknet_1_0__leaf_net119),
    .A3(net127),
    .S0(clknet_1_0__leaf_net134),
    .S1(clknet_1_0__leaf_net767),
    .X(net135));
 sky130_fd_sc_hd__a2111o_1 c195 (.A1(clknet_1_1__leaf_net134),
    .A2(clknet_1_0__leaf_net133),
    .B1(net131),
    .C1(net116),
    .X(net136));
 sky130_fd_sc_hd__mux4_1 c196 (.A0(clknet_1_1__leaf_net118),
    .A1(clknet_1_0__leaf_net128),
    .A2(net129),
    .A3(net127),
    .S0(net700),
    .S1(clknet_1_1__leaf_net767),
    .X(net137));
 sky130_fd_sc_hd__a2111o_1 c197 (.A1(net137),
    .A2(clknet_1_1__leaf_net128),
    .B1(net131),
    .C1(clknet_1_1__leaf_net118),
    .D1(net701),
    .X(net138));
 sky130_fd_sc_hd__buf_1 c198 (.A(net724),
    .X(net139));
 sky130_fd_sc_hd__buf_6 c199 (.A(net724),
    .X(net140));
 sky130_fd_sc_hd__and2_4 c200 (.A(net140),
    .B(net130),
    .X(net141));
 sky130_fd_sc_hd__and2_0 c201 (.A(net141),
    .B(net139),
    .X(net142));
 sky130_fd_sc_hd__and2_4 c202 (.A(net141),
    .B(net124),
    .X(net143));
 sky130_fd_sc_hd__and2_4 c203 (.A(net143),
    .B(net140),
    .X(net144));
 sky130_fd_sc_hd__and3_1 c204 (.A(net925),
    .B(net143),
    .C(net139),
    .X(net145));
 sky130_fd_sc_hd__and3_1 c205 (.A(net145),
    .B(net143),
    .C(net925),
    .X(net146));
 sky130_fd_sc_hd__and3_4 c206 (.A(net146),
    .B(net143),
    .C(net925),
    .X(net147));
 sky130_fd_sc_hd__or4bb_4 c207 (.A(net139),
    .B(net925),
    .C_N(net143),
    .D_N(net147),
    .X(net148));
 sky130_fd_sc_hd__and3_1 c208 (.A(net147),
    .B(net920),
    .C(net143),
    .X(net149));
 sky130_fd_sc_hd__and3_1 c209 (.A(net146),
    .B(net925),
    .C(net920),
    .X(net150));
 sky130_fd_sc_hd__a2111o_2 c210 (.A1(net140),
    .A2(net150),
    .B1(net147),
    .C1(net942),
    .D1(net143),
    .X(net151));
 sky130_fd_sc_hd__a2111o_1 c211 (.A1(net149),
    .A2(net147),
    .B1(net151),
    .C1(net937),
    .D1(net942),
    .X(net152));
 sky130_fd_sc_hd__mux4_1 c212 (.A0(net942),
    .A1(net150),
    .A2(net152),
    .A3(net151),
    .S0(net936),
    .S1(net929),
    .X(net153));
 sky130_fd_sc_hd__mux4_1 c213 (.A0(net152),
    .A1(net151),
    .A2(net153),
    .A3(net941),
    .S0(net116),
    .S1(net935),
    .X(net154));
 sky130_fd_sc_hd__a2111o_1 c214 (.A1(net153),
    .A2(net152),
    .B1(net940),
    .C1(net151),
    .D1(net150),
    .X(net155));
 sky130_fd_sc_hd__mux4_2 c215 (.A0(net142),
    .A1(net155),
    .A2(net147),
    .A3(net144),
    .S0(net970),
    .S1(net151),
    .X(net156));
 sky130_fd_sc_hd__a2111o_1 c216 (.A1(net156),
    .A2(net155),
    .B1(net147),
    .C1(net151),
    .D1(clknet_1_0__leaf_net768),
    .X(net157));
 sky130_fd_sc_hd__mux4_1 c217 (.A0(net145),
    .A1(clknet_1_0__leaf_net157),
    .A2(net156),
    .A3(net151),
    .S0(net149),
    .S1(clknet_1_0__leaf_net768),
    .X(net158));
 sky130_fd_sc_hd__mux4_1 c218 (.A0(clknet_1_0__leaf_net157),
    .A1(net142),
    .A2(net155),
    .A3(clknet_1_0__leaf_net158),
    .S0(net156),
    .S1(clknet_1_1__leaf_net768),
    .X(net159));
 sky130_fd_sc_hd__sdfbbn_1 c219 (.CLK_N(clknet_4_2_0_clk),
    .D(net151),
    .RESET_B(clknet_1_1__leaf_net158),
    .SCD(clknet_1_1__leaf_net157),
    .SCE(net156),
    .SET_B(net724),
    .Q(net161),
    .Q_N(net160));
 sky130_fd_sc_hd__and2_2 c220 (.A(net36),
    .B(net938),
    .X(net162));
 sky130_fd_sc_hd__and2_0 c221 (.A(net162),
    .B(net761),
    .X(net163));
 sky130_fd_sc_hd__and2_0 c222 (.A(net163),
    .B(net162),
    .X(net164));
 sky130_fd_sc_hd__and2_1 c223 (.A(net162),
    .B(net938),
    .X(net165));
 sky130_fd_sc_hd__buf_1 c224 (.A(clknet_1_1__leaf_net737),
    .X(net166));
 sky130_fd_sc_hd__and3_2 c225 (.A(net929),
    .B(net162),
    .C(net165),
    .X(net167));
 sky130_fd_sc_hd__and2_0 c226 (.A(net165),
    .B(clknet_1_0__leaf_net166),
    .X(net168));
 sky130_fd_sc_hd__buf_1 c227 (.A(clknet_1_1__leaf_net737),
    .X(net169));
 sky130_fd_sc_hd__buf_1 c228 (.A(net742),
    .X(net170));
 sky130_fd_sc_hd__clkbuf_2 c229 (.A(net752),
    .X(net171));
 sky130_fd_sc_hd__clkbuf_2 c230 (.A(net756),
    .X(net172));
 sky130_fd_sc_hd__mux4_1 c231 (.A0(net171),
    .A1(clknet_1_1__leaf_net169),
    .A2(clknet_1_0__leaf_net168),
    .A3(net162),
    .S0(net165),
    .S1(net167),
    .X(net173));
 sky130_fd_sc_hd__and3_1 c232 (.A(net172),
    .B(net171),
    .C(net165),
    .X(net174));
 sky130_fd_sc_hd__or4bb_1 c233 (.A(clknet_1_1__leaf_net166),
    .B(net172),
    .C_N(net171),
    .D_N(clknet_1_1__leaf_net769),
    .X(net175));
 sky130_fd_sc_hd__a2111o_1 c234 (.A1(clknet_1_0__leaf_net169),
    .A2(clknet_1_1__leaf_net175),
    .B1(net172),
    .C1(net162),
    .D1(net171),
    .X(net176));
 sky130_fd_sc_hd__mux4_1 c235 (.A0(net170),
    .A1(net162),
    .A2(net167),
    .A3(net171),
    .S0(clknet_1_1__leaf_net175),
    .S1(net172),
    .X(net177));
 sky130_fd_sc_hd__mux4_1 c236 (.A0(net41),
    .A1(clknet_1_0__leaf_net175),
    .A2(net167),
    .A3(net148),
    .S0(clknet_1_0__leaf_net769),
    .S1(net771),
    .X(net178));
 sky130_fd_sc_hd__mux4_1 c237 (.A0(clknet_1_1__leaf_net175),
    .A1(net174),
    .A2(net171),
    .A3(net172),
    .S0(net770),
    .S1(net773),
    .X(net179));
 sky130_fd_sc_hd__mux4_1 c238 (.A0(clknet_1_0__leaf_net175),
    .A1(net171),
    .A2(net162),
    .A3(net740),
    .S0(net771),
    .S1(net773),
    .X(net180));
 sky130_fd_sc_hd__mux4_1 c239 (.A0(net174),
    .A1(clknet_1_0__leaf_net176),
    .A2(net172),
    .A3(clknet_1_1__leaf_net175),
    .S0(clknet_1_0__leaf_net769),
    .S1(net773),
    .X(net181));
 sky130_fd_sc_hd__mux4_1 c240 (.A0(clknet_1_0__leaf_net180),
    .A1(clknet_1_0__leaf_net175),
    .A2(net161),
    .A3(clknet_1_0__leaf_net737),
    .S0(net771),
    .S1(net772),
    .X(net182));
 sky130_fd_sc_hd__mux4_1 c241 (.A0(clknet_1_1__leaf_net180),
    .A1(net182),
    .A2(clknet_1_0__leaf_net175),
    .A3(clknet_1_0__leaf_net737),
    .S0(net770),
    .S1(net773),
    .X(net183));
 sky130_fd_sc_hd__clkbuf_1 c242 (.A(net662),
    .X(net184));
 sky130_fd_sc_hd__and2_0 c243 (.A(net184),
    .B(net772),
    .X(net185));
 sky130_fd_sc_hd__and3_1 c244 (.A(net61),
    .B(net185),
    .C(net772),
    .X(net186));
 sky130_fd_sc_hd__buf_1 c245 (.A(net662),
    .X(net187));
 sky130_fd_sc_hd__and2_1 c246 (.A(net186),
    .B(net52),
    .X(net188));
 sky130_fd_sc_hd__and2_0 c247 (.A(net185),
    .B(net187),
    .X(net189));
 sky130_fd_sc_hd__and3_1 c248 (.A(net187),
    .B(net186),
    .C(net923),
    .X(net190));
 sky130_fd_sc_hd__and3_1 c249 (.A(net924),
    .B(net190),
    .C(net188),
    .X(net191));
 sky130_fd_sc_hd__and3_1 c250 (.A(clknet_1_1__leaf_net176),
    .B(net184),
    .C(net923),
    .X(net192));
 sky130_fd_sc_hd__and2_2 c251 (.A(net184),
    .B(net923),
    .X(net193));
 sky130_fd_sc_hd__or4bb_1 c252 (.A(net193),
    .B(net185),
    .C_N(net52),
    .D_N(net923),
    .X(net194));
 sky130_fd_sc_hd__sdfrtp_1 c253 (.CLK(clknet_4_10_0_clk),
    .D(net52),
    .RESET_B(clknet_1_0__leaf_net192),
    .SCD(net193),
    .SCE(net923),
    .Q(net906));
 sky130_fd_sc_hd__or4bb_1 c254 (.A(net194),
    .B(net193),
    .C_N(net906),
    .D_N(net923),
    .X(net195));
 sky130_fd_sc_hd__a2111o_1 c255 (.A1(net195),
    .A2(net188),
    .B1(net194),
    .C1(net193),
    .D1(net923),
    .X(net196));
 sky130_fd_sc_hd__sdfbbp_1 c256 (.CLK(clknet_4_10_0_clk),
    .D(clknet_1_1__leaf_net192),
    .RESET_B(net193),
    .SCD(net194),
    .SCE(net923),
    .SET_B(net196),
    .Q(net198),
    .Q_N(net197));
 sky130_fd_sc_hd__a2111o_1 c257 (.A1(net196),
    .A2(net191),
    .B1(net956),
    .C1(net193),
    .D1(net924),
    .X(net199));
 sky130_fd_sc_hd__mux4_2 c258 (.A0(net906),
    .A1(net193),
    .A2(net195),
    .A3(net923),
    .S0(net187),
    .S1(net707),
    .X(net200));
 sky130_fd_sc_hd__mux4_1 c259 (.A0(net191),
    .A1(net200),
    .A2(net195),
    .A3(net924),
    .S0(net193),
    .S1(net706),
    .X(net201));
 sky130_fd_sc_hd__mux4_1 c260 (.A0(net188),
    .A1(net200),
    .A2(net191),
    .A3(net923),
    .S0(net742),
    .S1(net962),
    .X(net202));
 sky130_fd_sc_hd__mux4_1 c261 (.A0(net59),
    .A1(net200),
    .A2(net193),
    .A3(net190),
    .S0(net197),
    .S1(net775),
    .X(net203));
 sky130_fd_sc_hd__mux4_1 c262 (.A0(net203),
    .A1(net196),
    .A2(net200),
    .A3(net924),
    .S0(net193),
    .S1(net775),
    .X(net204));
 sky130_fd_sc_hd__mux4_1 c263 (.A0(net198),
    .A1(net200),
    .A2(net924),
    .A3(net203),
    .S0(net707),
    .S1(net776),
    .X(net205));
 sky130_fd_sc_hd__and2_1 c264 (.A(net73),
    .B(net928),
    .X(net206));
 sky130_fd_sc_hd__and2_1 c265 (.A(net922),
    .B(net84),
    .X(net207));
 sky130_fd_sc_hd__and2_2 c266 (.A(net207),
    .B(net922),
    .X(net208));
 sky130_fd_sc_hd__or4bb_1 c267 (.A(net922),
    .B(net208),
    .C_N(net207),
    .D_N(net754),
    .X(net209));
 sky130_fd_sc_hd__and2_1 c268 (.A(net207),
    .B(net208),
    .X(net210));
 sky130_fd_sc_hd__and3_2 c269 (.A(net210),
    .B(net922),
    .C(net927),
    .X(net211));
 sky130_fd_sc_hd__and3_1 c270 (.A(net922),
    .B(net208),
    .C(net210),
    .X(net212));
 sky130_fd_sc_hd__and3_1 c271 (.A(net211),
    .B(net212),
    .C(net208),
    .X(net213));
 sky130_fd_sc_hd__buf_1 c272 (.X(net214));
 sky130_fd_sc_hd__and3_1 c273 (.A(net84),
    .B(net211),
    .C(net208),
    .X(net215));
 sky130_fd_sc_hd__clkbuf_1 c274 (.A(net674),
    .X(net216));
 sky130_fd_sc_hd__and2_1 c275 (.A(net208),
    .B(net216),
    .X(net217));
 sky130_fd_sc_hd__buf_1 c276 (.A(clknet_1_0__leaf_net825),
    .X(net218));
 sky130_fd_sc_hd__and2_1 c277 (.A(net217),
    .B(net208),
    .X(net219));
 sky130_fd_sc_hd__mux4_1 c278 (.A0(net219),
    .A1(net217),
    .A2(net213),
    .A3(net212),
    .S0(net922),
    .S1(net211),
    .X(net220));
 sky130_fd_sc_hd__a2111o_1 c279 (.A1(net212),
    .A2(net219),
    .B1(net213),
    .C1(net211),
    .D1(net208),
    .X(net221));
 sky130_fd_sc_hd__sdfbbn_1 c280 (.CLK_N(clknet_4_0_0_clk),
    .D(net215),
    .RESET_B(net217),
    .SCD(net219),
    .SCE(net212),
    .SET_B(net210),
    .Q(net223),
    .Q_N(net222));
 sky130_fd_sc_hd__and3_1 c281 (.A(net223),
    .B(net219),
    .C(net217),
    .X(net224));
 sky130_fd_sc_hd__a2111o_1 c282 (.A1(net218),
    .A2(net224),
    .B1(net222),
    .C1(net213),
    .D1(net730),
    .X(net225));
 sky130_fd_sc_hd__a2111o_1 c283 (.A1(net224),
    .A2(net210),
    .B1(net219),
    .C1(net730),
    .D1(net739),
    .X(net226));
 sky130_fd_sc_hd__mux4_1 c284 (.A0(net207),
    .A1(net223),
    .A2(net224),
    .A3(net219),
    .S0(net211),
    .X(net227));
 sky130_fd_sc_hd__sdfbbn_1 c285 (.CLK_N(clknet_4_0_0_clk),
    .D(net224),
    .RESET_B(net211),
    .SCD(net208),
    .SCE(net222),
    .SET_B(net759),
    .Q(net229),
    .Q_N(net228));
 sky130_fd_sc_hd__and3_1 c286 (.A(net229),
    .B(net96),
    .C(net104),
    .X(net230));
 sky130_fd_sc_hd__and2_1 c287 (.A(net915),
    .B(net104),
    .X(net231));
 sky130_fd_sc_hd__buf_1 c288 (.A(net951),
    .X(net232));
 sky130_fd_sc_hd__dlymetal6s2s_1 c289 (.A(net744),
    .X(net233));
 sky130_fd_sc_hd__and2_1 c290 (.A(net922),
    .B(net915),
    .X(net234));
 sky130_fd_sc_hd__dfbbn_1 c291 (.CLK_N(clknet_4_1_0_clk),
    .D(net231),
    .RESET_B(net233),
    .SET_B(net915),
    .Q(net236),
    .Q_N(net235));
 sky130_fd_sc_hd__sdfrtp_1 c292 (.CLK(clknet_4_1_0_clk),
    .D(net234),
    .RESET_B(net866),
    .SCD(net233),
    .SCE(net916),
    .Q(net237));
 sky130_fd_sc_hd__buf_1 c293 (.A(clknet_1_1__leaf_net825),
    .X(net238));
 sky130_fd_sc_hd__and2_0 c294 (.A(net916),
    .B(clknet_1_1__leaf_net238),
    .X(net239));
 sky130_fd_sc_hd__sdfsbp_1 c295 (.CLK(clknet_4_1_0_clk),
    .D(net233),
    .SCD(net232),
    .SCE(clknet_1_0__leaf_net239),
    .SET_B(net916),
    .Q(net241),
    .Q_N(net240));
 sky130_fd_sc_hd__sdfsbp_1 c296 (.CLK(clknet_4_1_0_clk),
    .D(net954),
    .SCD(net231),
    .SCE(net949),
    .SET_B(net916),
    .Q(net243),
    .Q_N(net242));
 sky130_fd_sc_hd__sdfstp_1 c297 (.CLK(clknet_4_1_0_clk),
    .D(net232),
    .SCD(net954),
    .SCE(net234),
    .SET_B(net916),
    .Q(net244));
 sky130_fd_sc_hd__sdfbbp_1 c298 (.CLK(clknet_4_1_0_clk),
    .D(clknet_1_0__leaf_net239),
    .RESET_B(net233),
    .SCD(net960),
    .SCE(net916),
    .SET_B(net949),
    .Q(net246),
    .Q_N(net245));
 sky130_fd_sc_hd__mux4_1 c299 (.A0(net241),
    .A1(net237),
    .A2(net246),
    .A3(net242),
    .S0(clknet_1_1__leaf_net239),
    .S1(net916),
    .X(net247));
 sky130_fd_sc_hd__mux4_1 c300 (.A0(net244),
    .A1(clknet_1_0__leaf_net238),
    .A2(net245),
    .A3(net234),
    .S0(net916),
    .S1(net778),
    .X(net248));
 sky130_fd_sc_hd__a2111o_1 c301 (.A1(net246),
    .A2(net235),
    .B1(net915),
    .C1(net778),
    .D1(net779),
    .X(net249));
 sky130_fd_sc_hd__mux4_1 c302 (.A0(net243),
    .A1(net249),
    .A2(net234),
    .A3(net233),
    .S0(net915),
    .S1(net779),
    .X(net250));
 sky130_fd_sc_hd__a2111o_1 c303 (.A1(clknet_1_0__leaf_net238),
    .A2(net244),
    .B1(net915),
    .C1(net779),
    .D1(net780),
    .X(net251));
 sky130_fd_sc_hd__mux4_1 c304 (.A0(net236),
    .A1(net241),
    .A2(net915),
    .A3(net778),
    .S0(net779),
    .S1(net780),
    .X(net252));
 sky130_fd_sc_hd__mux4_1 c305 (.A0(net252),
    .A1(net241),
    .A2(net249),
    .A3(clknet_1_0__leaf_net251),
    .S0(net779),
    .S1(net780),
    .X(net253));
 sky130_fd_sc_hd__mux4_1 c306 (.A0(clknet_1_0__leaf_net251),
    .A1(net922),
    .A2(net915),
    .A3(net778),
    .S0(net779),
    .S1(net780),
    .X(net254));
 sky130_fd_sc_hd__a2111o_1 c307 (.A1(net915),
    .A2(net738),
    .B1(net778),
    .C1(net779),
    .D1(net780),
    .X(net255));
 sky130_fd_sc_hd__and2_0 c308 (.A(net138),
    .B(net104),
    .X(net256));
 sky130_fd_sc_hd__and2_0 c309 (.A(clknet_1_0__leaf_net256),
    .B(net104),
    .X(net257));
 sky130_fd_sc_hd__clkbuf_2 c310 (.A(net678),
    .X(net258));
 sky130_fd_sc_hd__clkbuf_1 c311 (.A(net678),
    .X(net259));
 sky130_fd_sc_hd__clkbuf_2 c312 (.A(net829),
    .X(net260));
 sky130_fd_sc_hd__buf_1 c313 (.X(net261));
 sky130_fd_sc_hd__and2_1 c314 (.A(net258),
    .B(net261),
    .X(net262));
 sky130_fd_sc_hd__and2_0 c315 (.A(net259),
    .B(net261),
    .X(net263));
 sky130_fd_sc_hd__buf_1 c316 (.A(net683),
    .X(net264));
 sky130_fd_sc_hd__and2_0 c317 (.A(clknet_1_0__leaf_net256),
    .B(net264),
    .X(net265));
 sky130_fd_sc_hd__sdfstp_1 c318 (.CLK(clknet_4_3_0_clk),
    .D(clknet_1_1__leaf_net251),
    .SCD(net264),
    .SCE(clknet_1_0__leaf_net257),
    .SET_B(clknet_1_0__leaf_net256),
    .Q(net266));
 sky130_fd_sc_hd__and3_2 c319 (.A(net262),
    .B(net266),
    .C(net228),
    .X(net267));
 sky130_fd_sc_hd__sdfbbn_1 c320 (.CLK_N(clknet_4_3_0_clk),
    .D(net265),
    .RESET_B(net266),
    .SCD(net264),
    .SCE(net262),
    .SET_B(net258),
    .Q(net269),
    .Q_N(net268));
 sky130_fd_sc_hd__mux4_1 c321 (.A0(net267),
    .A1(net262),
    .A2(clknet_1_1__leaf_net256),
    .A3(net266),
    .S0(net258),
    .S1(net261),
    .X(net270));
 sky130_fd_sc_hd__mux4_1 c322 (.A0(net264),
    .A1(net269),
    .A2(clknet_1_1__leaf_net257),
    .A3(net262),
    .S0(net258),
    .S1(net267),
    .X(net271));
 sky130_fd_sc_hd__mux4_1 c323 (.A0(net260),
    .A1(clknet_1_0__leaf_net256),
    .A2(net268),
    .A3(net267),
    .S0(clknet_1_0__leaf_net270),
    .S1(net710),
    .X(net272));
 sky130_fd_sc_hd__mux4_1 c324 (.A0(net266),
    .A1(net261),
    .A2(net267),
    .A3(net268),
    .S0(clknet_1_0__leaf_net270),
    .S1(net782),
    .X(net273));
 sky130_fd_sc_hd__mux4_1 c325 (.A0(net269),
    .A1(net260),
    .A2(net267),
    .A3(clknet_1_1__leaf_net256),
    .S0(clknet_1_0__leaf_net270),
    .S1(net266),
    .X(net274));
 sky130_fd_sc_hd__mux4_1 c326 (.A0(clknet_1_0__leaf_net270),
    .A1(net266),
    .A2(net267),
    .A3(net258),
    .S0(clknet_1_1__leaf_net256),
    .S1(net743),
    .X(net275));
 sky130_fd_sc_hd__mux4_1 c327 (.A0(net263),
    .A1(net269),
    .A2(clknet_1_0__leaf_net270),
    .A3(net267),
    .S0(clknet_1_1__leaf_net256),
    .S1(net781),
    .X(net276));
 sky130_fd_sc_hd__a2111o_1 c328 (.A1(clknet_1_0__leaf_net270),
    .A2(net264),
    .B1(net262),
    .C1(net709),
    .D1(net783),
    .X(net277));
 sky130_fd_sc_hd__mux4_1 c329 (.A0(net258),
    .A1(net261),
    .A2(clknet_1_1__leaf_net270),
    .A3(net266),
    .S0(net747),
    .S1(net784),
    .X(net278));
 sky130_fd_sc_hd__clkbuf_1 c330 (.A(net673),
    .X(net279));
 sky130_fd_sc_hd__and2_1 c331 (.A(net279),
    .B(net161),
    .X(net280));
 sky130_fd_sc_hd__clkbuf_1 c332 (.A(net673),
    .X(net281));
 sky130_fd_sc_hd__and2_1 c333 (.A(net280),
    .B(net281),
    .X(net282));
 sky130_fd_sc_hd__and3_4 c334 (.A(net920),
    .B(net280),
    .C(net282),
    .X(net283));
 sky130_fd_sc_hd__and2_2 c335 (.A(net282),
    .B(net280),
    .X(net284));
 sky130_fd_sc_hd__and2_1 c336 (.A(net282),
    .B(net284),
    .X(net285));
 sky130_fd_sc_hd__and3_1 c337 (.A(net260),
    .B(net284),
    .C(net282),
    .X(net286));
 sky130_fd_sc_hd__and3_1 c338 (.A(net284),
    .B(net280),
    .C(net748),
    .X(net287));
 sky130_fd_sc_hd__buf_1 c339 (.A(clknet_1_0__leaf_net736),
    .X(net288));
 sky130_fd_sc_hd__mux4_2 c340 (.A0(net281),
    .A1(clknet_1_0__leaf_net288),
    .A2(net286),
    .A3(net280),
    .S0(net283),
    .S1(net282),
    .X(net289));
 sky130_fd_sc_hd__or4bb_4 c341 (.A(net287),
    .B(clknet_1_0__leaf_net289),
    .C_N(net283),
    .D_N(net284),
    .X(net290));
 sky130_fd_sc_hd__a2111o_1 c342 (.A1(clknet_1_0__leaf_net288),
    .A2(net285),
    .B1(clknet_1_1__leaf_net289),
    .C1(clknet_1_0__leaf_net290),
    .D1(net282),
    .X(net291));
 sky130_fd_sc_hd__mux4_2 c343 (.A0(net279),
    .A1(net287),
    .A2(clknet_1_0__leaf_net290),
    .A3(clknet_1_0__leaf_net289),
    .S0(clknet_1_0__leaf_net288),
    .S1(net280),
    .X(net292));
 sky130_fd_sc_hd__a2111o_1 c344 (.A1(clknet_1_1__leaf_net292),
    .A2(net283),
    .B1(clknet_1_0__leaf_net290),
    .C1(clknet_1_0__leaf_net291),
    .D1(clknet_1_1__leaf_net270),
    .X(net293));
 sky130_fd_sc_hd__and3_1 c345 (.A(net284),
    .B(clknet_1_1__leaf_net288),
    .C(clknet_1_0__leaf_net291),
    .X(net294));
 sky130_fd_sc_hd__mux4_2 c346 (.A0(clknet_1_1__leaf_net289),
    .A1(net285),
    .A2(clknet_1_0__leaf_net291),
    .A3(net280),
    .S0(clknet_1_0__leaf_net292),
    .S1(net732),
    .X(net295));
 sky130_fd_sc_hd__mux4_2 c347 (.A0(net285),
    .A1(clknet_1_0__leaf_net295),
    .A2(clknet_1_1__leaf_net288),
    .A3(clknet_1_1__leaf_net291),
    .S0(net284),
    .S1(clknet_1_0__leaf_net294),
    .X(net296));
 sky130_fd_sc_hd__a2111o_1 c348 (.A1(clknet_1_0__leaf_net296),
    .A2(clknet_1_1__leaf_net291),
    .B1(net286),
    .C1(clknet_1_1__leaf_net288),
    .D1(net970),
    .X(net297));
 sky130_fd_sc_hd__mux4_1 c349 (.A0(net280),
    .A1(clknet_1_0__leaf_net290),
    .A2(net283),
    .A3(clknet_1_1__leaf_net270),
    .S0(clknet_1_1__leaf_net291),
    .S1(clknet_1_0__leaf_net288),
    .X(net298));
 sky130_fd_sc_hd__mux4_2 c350 (.A0(clknet_1_1__leaf_net291),
    .A1(clknet_1_1__leaf_net295),
    .A2(clknet_1_0__leaf_net297),
    .A3(net285),
    .S0(clknet_1_1__leaf_net288),
    .S1(clknet_1_1__leaf_net736),
    .X(net299));
 sky130_fd_sc_hd__mux4_2 c351 (.A0(clknet_1_1__leaf_net297),
    .A1(clknet_1_1__leaf_net294),
    .A2(clknet_1_1__leaf_net296),
    .A3(clknet_1_0__leaf_net299),
    .S0(net284),
    .S1(clknet_1_1__leaf_net736),
    .X(net300));
 sky130_fd_sc_hd__clkbuf_2 c352 (.A(net669),
    .X(net301));
 sky130_fd_sc_hd__and2_0 c353 (.A(net301),
    .B(clknet_1_1__leaf_net769),
    .X(net302));
 sky130_fd_sc_hd__and2_0 c354 (.A(clknet_1_1__leaf_net290),
    .B(net740),
    .X(net303));
 sky130_fd_sc_hd__buf_1 c355 (.A(net669),
    .X(net304));
 sky130_fd_sc_hd__and3_1 c356 (.A(clknet_1_1__leaf_net290),
    .B(net301),
    .C(net304),
    .X(net305));
 sky130_fd_sc_hd__and3_1 c357 (.A(clknet_1_0__leaf_net302),
    .B(clknet_1_0__leaf_net303),
    .C(clknet_1_0__leaf_net305),
    .X(net306));
 sky130_fd_sc_hd__and3_1 c358 (.A(net304),
    .B(clknet_1_1__leaf_net303),
    .C(net301),
    .X(net307));
 sky130_fd_sc_hd__and3_1 c359 (.A(clknet_1_0__leaf_net306),
    .B(clknet_1_1__leaf_net307),
    .C(net304),
    .X(net308));
 sky130_fd_sc_hd__and3_1 c360 (.A(clknet_1_0__leaf_net308),
    .B(clknet_1_0__leaf_net303),
    .C(clknet_1_0__leaf_net307),
    .X(net309));
 sky130_fd_sc_hd__and3_1 c361 (.A(net301),
    .B(net304),
    .C(clknet_1_1__leaf_net303),
    .X(net310));
 sky130_fd_sc_hd__a2111o_1 c362 (.A1(clknet_1_0__leaf_net305),
    .A2(clknet_1_1__leaf_net308),
    .B1(net304),
    .C1(clknet_1_1__leaf_net290),
    .D1(clknet_1_0__leaf_net306),
    .X(net311));
 sky130_fd_sc_hd__or4bb_1 c363 (.A(net309),
    .B(clknet_1_1__leaf_net310),
    .C_N(clknet_1_1__leaf_net306),
    .D_N(net304),
    .X(net312));
 sky130_fd_sc_hd__mux4_1 c364 (.A0(clknet_1_0__leaf_net311),
    .A1(clknet_1_1__leaf_net307),
    .A2(clknet_1_0__leaf_net312),
    .A3(net304),
    .S0(clknet_1_1__leaf_net303),
    .S1(clknet_1_1__leaf_net305),
    .X(net313));
 sky130_fd_sc_hd__mux4_1 c365 (.A0(clknet_1_0__leaf_net302),
    .A1(clknet_1_0__leaf_net307),
    .A2(clknet_1_0__leaf_net308),
    .A3(clknet_1_0__leaf_net303),
    .S0(clknet_1_0__leaf_net310),
    .S1(net908),
    .X(net314));
 sky130_fd_sc_hd__sdfbbn_1 c366 (.CLK_N(clknet_4_8_0_clk),
    .D(clknet_1_0__leaf_net310),
    .RESET_B(clknet_1_1__leaf_net312),
    .SCD(clknet_1_0__leaf_net314),
    .SCE(clknet_1_1__leaf_net306),
    .SET_B(net301),
    .Q(net316),
    .Q_N(net315));
 sky130_fd_sc_hd__and3_1 c367 (.A(net283),
    .B(clknet_1_0__leaf_net314),
    .C(net316),
    .X(net317));
 sky130_fd_sc_hd__mux4_1 c368 (.A0(clknet_1_1__leaf_net303),
    .A1(clknet_1_0__leaf_net314),
    .A2(clknet_1_1__leaf_net310),
    .A3(clknet_1_0__leaf_net317),
    .S0(clknet_1_0__leaf_net312),
    .S1(net908),
    .X(net318));
 sky130_fd_sc_hd__a2111o_1 c369 (.A1(clknet_1_1__leaf_net317),
    .A2(clknet_1_1__leaf_net312),
    .B1(clknet_1_1__leaf_net314),
    .C1(net301),
    .D1(net785),
    .X(net319));
 sky130_fd_sc_hd__mux4_1 c370 (.A0(clknet_1_1__leaf_net312),
    .A1(clknet_1_0__leaf_net311),
    .A2(clknet_1_1__leaf_net314),
    .A3(clknet_1_1__leaf_net317),
    .S0(net908),
    .S1(net785),
    .X(net320));
 sky130_fd_sc_hd__a2111o_1 c371 (.A1(clknet_1_1__leaf_net314),
    .A2(net315),
    .B1(clknet_1_0__leaf_net317),
    .C1(net705),
    .D1(net785),
    .X(net321));
 sky130_fd_sc_hd__a2111o_1 c372 (.A1(net301),
    .A2(clknet_1_1__leaf_net311),
    .B1(net705),
    .C1(net752),
    .D1(net785),
    .X(net322));
 sky130_fd_sc_hd__mux4_1 c373 (.A0(net316),
    .A1(net322),
    .A2(clknet_1_1__leaf_net314),
    .A3(net705),
    .S0(net752),
    .S1(net785),
    .X(net323));
 sky130_fd_sc_hd__or4bb_1 c392 (.A(net906),
    .B(net776),
    .C_N(net908),
    .D_N(net899),
    .X(net912));
 sky130_fd_sc_hd__sdfstp_1 c393 (.CLK(clknet_4_10_0_clk),
    .D(net912),
    .SCD(net167),
    .SCE(net776),
    .SET_B(net777),
    .Q(net911));
 sky130_fd_sc_hd__mux4_1 c394 (.A0(net911),
    .A1(net912),
    .A2(clknet_1_1__leaf_net290),
    .A3(net776),
    .S0(net777),
    .S1(net908),
    .X(net910));
 sky130_fd_sc_hd__a2111o_1 c395 (.A1(net190),
    .A2(clknet_1_0__leaf_net910),
    .B1(net912),
    .C1(net911),
    .D1(net899),
    .X(net913));
 sky130_fd_sc_hd__and2_1 c396 (.A(net206),
    .B(net758),
    .X(net324));
 sky130_fd_sc_hd__and2_0 c397 (.A(net921),
    .B(net928),
    .X(net325));
 sky130_fd_sc_hd__and2_1 c398 (.A(net921),
    .B(net206),
    .X(net326));
 sky130_fd_sc_hd__and3_1 c399 (.A(net921),
    .B(net326),
    .C(net325),
    .X(net327));
 sky130_fd_sc_hd__and2_1 c400 (.A(net326),
    .B(net327),
    .X(net328));
 sky130_fd_sc_hd__and3_1 c401 (.A(net327),
    .B(net328),
    .C(net921),
    .X(net329));
 sky130_fd_sc_hd__and3_1 c402 (.A(net329),
    .B(net327),
    .C(net922),
    .X(net330));
 sky130_fd_sc_hd__and3_1 c403 (.A(net326),
    .B(net921),
    .C(net329),
    .X(net331));
 sky130_fd_sc_hd__and3_1 c404 (.A(net331),
    .B(net330),
    .C(net328),
    .X(net332));
 sky130_fd_sc_hd__or4bb_2 c405 (.A(net328),
    .B(net331),
    .C_N(net325),
    .D_N(net921),
    .X(net333));
 sky130_fd_sc_hd__and3_1 c406 (.A(net332),
    .B(net333),
    .C(net328),
    .X(net334));
 sky130_fd_sc_hd__and2_1 c407 (.A(net330),
    .B(net333),
    .X(net335));
 sky130_fd_sc_hd__and3_1 c408 (.A(net334),
    .B(net328),
    .C(net921),
    .X(net336));
 sky130_fd_sc_hd__a2111o_1 c409 (.A1(net326),
    .A2(net336),
    .B1(net328),
    .C1(net921),
    .D1(net329),
    .X(net337));
 sky130_fd_sc_hd__mux4_1 c410 (.A0(net325),
    .A1(net330),
    .A2(net327),
    .A3(net331),
    .S0(net921),
    .S1(net336),
    .X(net338));
 sky130_fd_sc_hd__mux4_1 c411 (.A0(net336),
    .A1(net333),
    .A2(net326),
    .A3(net327),
    .S0(net921),
    .S1(clknet_1_1__leaf_net786),
    .X(net339));
 sky130_fd_sc_hd__mux4_1 c412 (.A0(net335),
    .A1(net333),
    .A2(net327),
    .A3(net336),
    .S0(clknet_1_1__leaf_net786),
    .S1(clknet_1_1__leaf_net787),
    .X(net340));
 sky130_fd_sc_hd__a2111o_1 c413 (.A1(net335),
    .A2(net330),
    .B1(net324),
    .C1(net728),
    .D1(clknet_1_0__leaf_net786),
    .X(net341));
 sky130_fd_sc_hd__or4bb_1 c414 (.A(net333),
    .B(net330),
    .C_N(clknet_1_0__leaf_net786),
    .D_N(clknet_1_0__leaf_net787),
    .X(net342));
 sky130_fd_sc_hd__mux4_1 c415 (.A0(clknet_1_0__leaf_net341),
    .A1(net336),
    .A2(clknet_1_0__leaf_net342),
    .A3(net332),
    .S0(clknet_1_0__leaf_net786),
    .S1(clknet_1_0__leaf_net788),
    .X(net343));
 sky130_fd_sc_hd__or4bb_1 c416 (.A(clknet_1_0__leaf_net342),
    .B(clknet_1_0__leaf_net341),
    .C_N(net728),
    .D_N(clknet_1_0__leaf_net787),
    .X(net344));
 sky130_fd_sc_hd__mux4_1 c417 (.A0(net335),
    .A1(clknet_1_1__leaf_net341),
    .A2(net332),
    .A3(net330),
    .S0(clknet_1_1__leaf_net342),
    .S1(net744),
    .X(net345));
 sky130_fd_sc_hd__and2_0 c418 (.A(clknet_1_0__leaf_net788),
    .B(net790),
    .X(net346));
 sky130_fd_sc_hd__and2_0 c419 (.A(net324),
    .B(clknet_1_1__leaf_net346),
    .X(net347));
 sky130_fd_sc_hd__buf_1 c420 (.A(net745),
    .X(net348));
 sky130_fd_sc_hd__and2_0 c421 (.A(clknet_1_0__leaf_net346),
    .B(net348),
    .X(net349));
 sky130_fd_sc_hd__and2_0 c422 (.A(clknet_1_0__leaf_net346),
    .B(net348),
    .X(net350));
 sky130_fd_sc_hd__and2_0 c423 (.A(clknet_1_0__leaf_net349),
    .B(clknet_1_0__leaf_net346),
    .X(net351));
 sky130_fd_sc_hd__and2_0 c424 (.A(clknet_1_0__leaf_net350),
    .B(clknet_1_1__leaf_net346),
    .X(net352));
 sky130_fd_sc_hd__and2_0 c425 (.A(clknet_1_0__leaf_net347),
    .B(clknet_1_1__leaf_net350),
    .X(net353));
 sky130_fd_sc_hd__and2_0 c426 (.A(clknet_1_0__leaf_net353),
    .B(clknet_1_0__leaf_net350),
    .X(net354));
 sky130_fd_sc_hd__and2_0 c427 (.A(net348),
    .B(clknet_1_0__leaf_net353),
    .X(net355));
 sky130_fd_sc_hd__and3_1 c428 (.A(clknet_1_1__leaf_net354),
    .B(clknet_1_0__leaf_net353),
    .C(net348),
    .X(net356));
 sky130_fd_sc_hd__a2111o_1 c429 (.A1(clknet_1_0__leaf_net352),
    .A2(clknet_1_0__leaf_net356),
    .B1(net348),
    .C1(clknet_1_0__leaf_net353),
    .D1(clknet_1_1__leaf_net346),
    .X(net357));
 sky130_fd_sc_hd__a2111o_1 c430 (.A1(clknet_1_0__leaf_net354),
    .A2(clknet_1_0__leaf_net355),
    .B1(clknet_1_0__leaf_net353),
    .C1(net348),
    .D1(clknet_1_0__leaf_net346),
    .X(net358));
 sky130_fd_sc_hd__a2111o_1 c431 (.A1(clknet_1_1__leaf_net355),
    .A2(clknet_1_0__leaf_net350),
    .B1(clknet_1_0__leaf_net358),
    .C1(clknet_1_0__leaf_net353),
    .D1(clknet_1_1__leaf_net346),
    .X(net359));
 sky130_fd_sc_hd__a2111o_1 c432 (.A1(clknet_1_1__leaf_net347),
    .A2(clknet_1_1__leaf_net359),
    .B1(clknet_1_0__leaf_net356),
    .C1(clknet_1_1__leaf_net346),
    .D1(clknet_1_1__leaf_net358),
    .X(net360));
 sky130_fd_sc_hd__mux4_1 c433 (.A0(clknet_1_1__leaf_net357),
    .A1(clknet_1_1__leaf_net359),
    .A2(clknet_1_0__leaf_net360),
    .A3(clknet_1_1__leaf_net358),
    .S0(clknet_1_0__leaf_net356),
    .S1(clknet_1_0__leaf_net353),
    .X(net361));
 sky130_fd_sc_hd__a2111o_1 c434 (.A1(clknet_1_0__leaf_net360),
    .A2(clknet_1_1__leaf_net350),
    .B1(clknet_1_0__leaf_net359),
    .C1(clknet_1_1__leaf_net356),
    .D1(clknet_1_1__leaf_net361),
    .X(net362));
 sky130_fd_sc_hd__a2111o_1 c435 (.A1(clknet_1_0__leaf_net361),
    .A2(clknet_1_0__leaf_net359),
    .B1(clknet_1_0__leaf_net357),
    .C1(clknet_1_1__leaf_net352),
    .D1(clknet_1_0__leaf_net360),
    .X(net363));
 sky130_fd_sc_hd__mux4_1 c436 (.A0(clknet_1_1__leaf_net356),
    .A1(clknet_1_1__leaf_net358),
    .A2(clknet_1_1__leaf_net359),
    .A3(clknet_1_1__leaf_net360),
    .S0(clknet_1_1__leaf_net350),
    .S1(clknet_1_0__leaf_net362),
    .X(net364));
 sky130_fd_sc_hd__mux4_1 c437 (.A0(clknet_1_1__leaf_net351),
    .A1(clknet_1_0__leaf_net363),
    .A2(clknet_1_1__leaf_net360),
    .A3(clknet_1_1__leaf_net356),
    .S0(clknet_1_0__leaf_net359),
    .X(net365));
 sky130_fd_sc_hd__a2111o_1 c438 (.A1(clknet_1_1__leaf_net362),
    .A2(clknet_1_1__leaf_net360),
    .B1(clknet_1_1__leaf_net359),
    .C1(clknet_1_0__leaf_net358),
    .D1(net716),
    .X(net366));
 sky130_fd_sc_hd__a2111o_1 c439 (.A1(clknet_1_0__leaf_net358),
    .A2(clknet_1_0__leaf_net351),
    .B1(clknet_1_0__leaf_net359),
    .C1(net717),
    .D1(net745),
    .X(net367));
 sky130_fd_sc_hd__and2_0 c440 (.A(clknet_1_1__leaf_net349),
    .B(net260),
    .X(net368));
 sky130_fd_sc_hd__clkbuf_2 c441 (.A(net824),
    .X(net369));
 sky130_fd_sc_hd__and2_0 c442 (.A(clknet_1_1__leaf_net367),
    .B(clknet_1_0__leaf_net368),
    .X(net370));
 sky130_fd_sc_hd__and3_1 c443 (.A(net369),
    .B(clknet_1_0__leaf_net368),
    .C(clknet_1_0__leaf_net359),
    .X(net371));
 sky130_fd_sc_hd__and3_1 c444 (.A(clknet_1_0__leaf_net371),
    .B(clknet_1_1__leaf_net353),
    .C(clknet_1_1__leaf_net368),
    .X(net372));
 sky130_fd_sc_hd__or4bb_1 c445 (.A(clknet_1_0__leaf_net371),
    .B(clknet_1_1__leaf_net368),
    .C_N(net369),
    .D_N(clknet_1_0__leaf_net372),
    .X(net373));
 sky130_fd_sc_hd__buf_1 c446 (.A(net824),
    .X(net374));
 sky130_fd_sc_hd__and3_1 c447 (.A(net374),
    .B(clknet_1_0__leaf_net371),
    .C(clknet_1_0__leaf_net372),
    .X(net375));
 sky130_fd_sc_hd__and3_1 c448 (.A(clknet_1_1__leaf_net368),
    .B(net374),
    .C(net369),
    .X(net376));
 sky130_fd_sc_hd__sedfxbp_1 c449 (.CLK(clknet_4_4_0_clk),
    .D(clknet_1_0__leaf_net375),
    .DE(clknet_1_0__leaf_net373),
    .SCD(clknet_1_0__leaf_net372),
    .SCE(clknet_1_0__leaf_net371),
    .Q(net378),
    .Q_N(net377));
 sky130_fd_sc_hd__a2111o_1 c450 (.A1(clknet_1_0__leaf_net376),
    .A2(clknet_1_1__leaf_net375),
    .B1(clknet_1_1__leaf_net368),
    .C1(net377),
    .D1(clknet_1_0__leaf_net373),
    .X(net379));
 sky130_fd_sc_hd__or4bb_1 c451 (.A(clknet_1_1__leaf_net353),
    .B(clknet_1_0__leaf_net371),
    .C_N(net374),
    .D_N(net377),
    .X(net380));
 sky130_fd_sc_hd__a2111o_1 c452 (.A1(net370),
    .A2(net374),
    .B1(net369),
    .C1(clknet_1_1__leaf_net353),
    .D1(net720),
    .X(net381));
 sky130_fd_sc_hd__sdfbbp_1 c453 (.CLK(clknet_4_3_0_clk),
    .D(clknet_1_0__leaf_net380),
    .RESET_B(net966),
    .SCD(clknet_1_0__leaf_net373),
    .SCE(clknet_1_0__leaf_net372),
    .SET_B(net952),
    .Q(net383),
    .Q_N(net382));
 sky130_fd_sc_hd__sdfbbn_1 c454 (.CLK_N(clknet_4_6_0_clk),
    .D(clknet_1_0__leaf_net381),
    .RESET_B(net943),
    .SCD(net377),
    .SCE(clknet_1_0__leaf_net372),
    .SET_B(clknet_1_0__leaf_net376),
    .Q(net385),
    .Q_N(net384));
 sky130_fd_sc_hd__or4bb_1 c455 (.A(clknet_1_1__leaf_net372),
    .B(net378),
    .C_N(net382),
    .D_N(clknet_1_1__leaf_net376),
    .X(net386));
 sky130_fd_sc_hd__sdfbbn_1 c456 (.CLK_N(clknet_4_6_0_clk),
    .D(clknet_1_1__leaf_net380),
    .RESET_B(clknet_1_0__leaf_net386),
    .SCD(net378),
    .SCE(clknet_1_1__leaf_net353),
    .SET_B(net745),
    .Q(net388),
    .Q_N(net387));
 sky130_fd_sc_hd__mux4_1 c457 (.A0(clknet_1_1__leaf_net386),
    .A1(net384),
    .A2(net382),
    .A3(net387),
    .S0(clknet_1_1__leaf_net371),
    .S1(net369),
    .X(net389));
 sky130_fd_sc_hd__mux4_1 c458 (.A0(net378),
    .A1(clknet_1_1__leaf_net386),
    .A2(clknet_1_1__leaf_net376),
    .A3(net260),
    .S0(net387),
    .S1(net719),
    .X(net390));
 sky130_fd_sc_hd__mux4_1 c459 (.A0(net385),
    .A1(net388),
    .A2(clknet_1_1__leaf_net371),
    .A3(net369),
    .S0(clknet_1_1__leaf_net386),
    .S1(net791),
    .X(net391));
 sky130_fd_sc_hd__mux4_1 c460 (.A0(net388),
    .A1(net943),
    .A2(clknet_1_1__leaf_net381),
    .A3(net378),
    .S0(clknet_1_0__leaf_net386),
    .S1(net793),
    .X(net392));
 sky130_fd_sc_hd__mux4_1 c461 (.A0(clknet_1_1__leaf_net372),
    .A1(clknet_1_0__leaf_net386),
    .A2(net369),
    .A3(net377),
    .S0(net743),
    .S1(net794),
    .X(net393));
 sky130_fd_sc_hd__buf_1 c462 (.A(clknet_1_1__leaf_net668),
    .X(net394));
 sky130_fd_sc_hd__and2_0 c463 (.A(clknet_1_0__leaf_net394),
    .B(net283),
    .X(net395));
 sky130_fd_sc_hd__buf_1 c464 (.A(clknet_1_0__leaf_net668),
    .X(net396));
 sky130_fd_sc_hd__and2_0 c465 (.A(clknet_1_0__leaf_net396),
    .B(net792),
    .X(net397));
 sky130_fd_sc_hd__and2_0 c466 (.A(clknet_1_1__leaf_net397),
    .B(clknet_1_0__leaf_net396),
    .X(net398));
 sky130_fd_sc_hd__and2_0 c467 (.A(clknet_1_1__leaf_net398),
    .B(clknet_1_1__leaf_net396),
    .X(net399));
 sky130_fd_sc_hd__and3_1 c468 (.A(clknet_1_0__leaf_net396),
    .B(clknet_1_0__leaf_net397),
    .C(net920),
    .X(net400));
 sky130_fd_sc_hd__and2_0 c469 (.A(clknet_1_0__leaf_net400),
    .B(clknet_1_1__leaf_net396),
    .X(net401));
 sky130_fd_sc_hd__and2_0 c470 (.A(clknet_1_0__leaf_net398),
    .B(clknet_1_1__leaf_net401),
    .X(net402));
 sky130_fd_sc_hd__a2111o_1 c471 (.A1(clknet_1_0__leaf_net402),
    .A2(clknet_1_1__leaf_net396),
    .B1(clknet_1_1__leaf_net400),
    .C1(clknet_1_1__leaf_net401),
    .D1(clknet_1_0__leaf_net399),
    .X(net403));
 sky130_fd_sc_hd__and3_1 c472 (.A(clknet_1_1__leaf_net399),
    .B(clknet_1_1__leaf_net401),
    .C(clknet_1_0__leaf_net402),
    .X(net404));
 sky130_fd_sc_hd__or4bb_1 c473 (.A(clknet_1_0__leaf_net403),
    .B(clknet_1_0__leaf_net394),
    .C_N(clknet_1_1__leaf_net401),
    .D_N(clknet_1_1__leaf_net402),
    .X(net405));
 sky130_fd_sc_hd__or4bb_1 c474 (.A(clknet_1_1__leaf_net404),
    .B(clknet_1_0__leaf_net402),
    .C_N(clknet_1_0__leaf_net403),
    .D_N(clknet_1_1__leaf_net401),
    .X(net406));
 sky130_fd_sc_hd__or4bb_1 c475 (.A(clknet_1_1__leaf_net406),
    .B(clknet_1_1__leaf_net404),
    .C_N(clknet_1_1__leaf_net400),
    .D_N(clknet_1_0__leaf_net401),
    .X(net407));
 sky130_fd_sc_hd__or4bb_1 c476 (.A(clknet_1_1__leaf_net394),
    .B(clknet_1_0__leaf_net406),
    .C_N(clknet_1_0__leaf_net400),
    .D_N(clknet_1_1__leaf_net401),
    .X(net408));
 sky130_fd_sc_hd__or4bb_1 c477 (.A(clknet_1_1__leaf_net408),
    .B(clknet_1_0__leaf_net401),
    .C_N(clknet_1_1__leaf_net406),
    .D_N(clknet_1_0__leaf_net404),
    .X(net409));
 sky130_fd_sc_hd__mux4_1 c478 (.A0(net405),
    .A1(clknet_1_0__leaf_net404),
    .A2(clknet_1_0__leaf_net408),
    .A3(clknet_1_0__leaf_net406),
    .S0(clknet_1_0__leaf_net401),
    .S1(clknet_1_1__leaf_net395),
    .X(net410));
 sky130_fd_sc_hd__mux4_1 c479 (.A0(clknet_1_1__leaf_net400),
    .A1(clknet_1_0__leaf_net407),
    .A2(clknet_1_1__leaf_net406),
    .A3(clknet_1_1__leaf_net408),
    .S0(clknet_1_1__leaf_net402),
    .S1(clknet_1_0__leaf_net401),
    .X(net411));
 sky130_fd_sc_hd__mux4_1 c480 (.A0(net409),
    .A1(clknet_1_1__leaf_net411),
    .A2(clknet_1_1__leaf_net408),
    .A3(clknet_1_1__leaf_net402),
    .S0(clknet_1_1__leaf_net401),
    .S1(clknet_1_0__leaf_net410),
    .X(net412));
 sky130_fd_sc_hd__mux4_1 c481 (.A0(clknet_1_0__leaf_net411),
    .A1(clknet_1_0__leaf_net406),
    .A2(clknet_1_0__leaf_net408),
    .A3(clknet_1_1__leaf_net394),
    .S0(clknet_1_0__leaf_net412),
    .S1(net733),
    .X(net413));
 sky130_fd_sc_hd__mux4_1 c482 (.A0(clknet_1_1__leaf_net412),
    .A1(clknet_1_0__leaf_net404),
    .A2(clknet_1_0__leaf_net408),
    .A3(clknet_1_1__leaf_net403),
    .S0(clknet_1_0__leaf_net401),
    .X(net414));
 sky130_fd_sc_hd__a2111o_1 c483 (.A1(clknet_1_1__leaf_net410),
    .A2(clknet_1_1__leaf_net407),
    .B1(clknet_1_1__leaf_net404),
    .C1(clknet_1_1__leaf_net408),
    .D1(net729),
    .X(net415));
 sky130_fd_sc_hd__and2_2 c484 (.A(net729),
    .B(net899),
    .X(net416));
 sky130_fd_sc_hd__buf_1 c485 (.A(net726),
    .X(net417));
 sky130_fd_sc_hd__and2_1 c486 (.A(net417),
    .B(net729),
    .X(net418));
 sky130_fd_sc_hd__and2_0 c487 (.A(net417),
    .B(net416),
    .X(net419));
 sky130_fd_sc_hd__and3_1 c488 (.A(net418),
    .B(net417),
    .C(net729),
    .X(net420));
 sky130_fd_sc_hd__and3_1 c489 (.A(net416),
    .B(net420),
    .C(net908),
    .X(net900));
 sky130_fd_sc_hd__and2_2 c490 (.A(net420),
    .B(net416),
    .X(net907));
 sky130_fd_sc_hd__or4bb_1 c491 (.A(net907),
    .B(net420),
    .C_N(net900),
    .D_N(net418),
    .X(net421));
 sky130_fd_sc_hd__and3_1 c492 (.A(net421),
    .B(net416),
    .C(net907),
    .X(net422));
 sky130_fd_sc_hd__and2_1 c493 (.A(net907),
    .B(net418),
    .X(net423));
 sky130_fd_sc_hd__and3_1 c494 (.A(net418),
    .B(net907),
    .C(net422),
    .X(net424));
 sky130_fd_sc_hd__or4bb_2 c495 (.A(net417),
    .B(net424),
    .C_N(net422),
    .D_N(net907),
    .X(net425));
 sky130_fd_sc_hd__a2111o_2 c496 (.A1(net424),
    .A2(net425),
    .B1(net417),
    .C1(net907),
    .D1(net423),
    .X(net904));
 sky130_fd_sc_hd__or4bb_2 c497 (.A(net422),
    .B(net904),
    .C_N(net424),
    .D_N(net418),
    .X(net426));
 sky130_fd_sc_hd__or4bb_2 c498 (.A(net420),
    .B(net904),
    .C_N(net426),
    .D_N(net423),
    .X(net427));
 sky130_fd_sc_hd__mux4_2 c499 (.A0(net904),
    .A1(net427),
    .A2(net907),
    .A3(net426),
    .S0(net425),
    .S1(net900),
    .X(net428));
 sky130_fd_sc_hd__mux4_2 c500 (.A0(net426),
    .A1(net428),
    .A2(net424),
    .A3(net425),
    .S0(net418),
    .S1(net907),
    .X(net903));
 sky130_fd_sc_hd__mux4_1 c501 (.A0(net423),
    .A1(net428),
    .A2(net427),
    .A3(net426),
    .S0(net903),
    .S1(net904),
    .X(net429));
 sky130_fd_sc_hd__mux4_1 c502 (.A0(net419),
    .A1(net429),
    .A2(net427),
    .A3(net428),
    .S0(clknet_1_1__leaf_net401),
    .S1(net903),
    .X(net430));
 sky130_fd_sc_hd__mux4_1 c503 (.A0(net167),
    .A1(clknet_1_1__leaf_net430),
    .A2(net903),
    .A3(net429),
    .S0(net428),
    .S1(net427),
    .X(net431));
 sky130_fd_sc_hd__mux4_1 c504 (.A0(net422),
    .A1(net426),
    .A2(net429),
    .A3(clknet_1_0__leaf_net430),
    .S0(net904),
    .S1(net726),
    .X(net432));
 sky130_fd_sc_hd__mux4_1 c505 (.A0(net425),
    .A1(net432),
    .A2(clknet_1_0__leaf_net430),
    .A3(net429),
    .S0(net426),
    .S1(net726),
    .X(net433));
 sky130_fd_sc_hd__and2_0 c528 (.A(net928),
    .B(clknet_1_0__leaf_net788),
    .X(net434));
 sky130_fd_sc_hd__and2_0 c529 (.A(clknet_1_0__leaf_net434),
    .B(net789),
    .X(net435));
 sky130_fd_sc_hd__and2_0 c530 (.A(clknet_1_0__leaf_net435),
    .B(clknet_1_1__leaf_net434),
    .X(net436));
 sky130_fd_sc_hd__and2_0 c531 (.A(clknet_1_1__leaf_net436),
    .B(clknet_1_1__leaf_net435),
    .X(net437));
 sky130_fd_sc_hd__and2_0 c532 (.A(clknet_1_0__leaf_net437),
    .B(clknet_1_1__leaf_net435),
    .X(net438));
 sky130_fd_sc_hd__and3_1 c533 (.A(clknet_1_0__leaf_net435),
    .B(clknet_1_0__leaf_net436),
    .C(clknet_1_1__leaf_net788),
    .X(net439));
 sky130_fd_sc_hd__and3_1 c534 (.A(clknet_1_1__leaf_net436),
    .B(clknet_1_1__leaf_net439),
    .C(clknet_1_1__leaf_net435),
    .X(net440));
 sky130_fd_sc_hd__and3_1 c535 (.A(clknet_1_0__leaf_net438),
    .B(clknet_1_0__leaf_net440),
    .C(clknet_1_0__leaf_net439),
    .X(net441));
 sky130_fd_sc_hd__and3_1 c536 (.A(clknet_1_1__leaf_net439),
    .B(clknet_1_0__leaf_net437),
    .C(clknet_1_1__leaf_net435),
    .X(net442));
 sky130_fd_sc_hd__and3_1 c537 (.A(clknet_1_0__leaf_net441),
    .B(clknet_1_0__leaf_net442),
    .C(net790),
    .X(net443));
 sky130_fd_sc_hd__and3_1 c538 (.A(clknet_1_0__leaf_net440),
    .B(clknet_1_0__leaf_net443),
    .C(clknet_1_1__leaf_net439),
    .X(net444));
 sky130_fd_sc_hd__and3_1 c539 (.A(clknet_1_1__leaf_net441),
    .B(clknet_1_0__leaf_net443),
    .C(clknet_1_0__leaf_net444),
    .X(net445));
 sky130_fd_sc_hd__mux4_1 c540 (.A0(clknet_1_1__leaf_net434),
    .A1(clknet_1_0__leaf_net445),
    .A2(clknet_1_0__leaf_net442),
    .A3(clknet_1_0__leaf_net439),
    .S0(clknet_1_0__leaf_net441),
    .S1(clknet_1_0__leaf_net444),
    .X(net446));
 sky130_fd_sc_hd__a2111o_1 c541 (.A1(clknet_1_0__leaf_net442),
    .A2(clknet_1_0__leaf_net436),
    .B1(clknet_1_0__leaf_net445),
    .C1(clknet_1_0__leaf_net435),
    .D1(clknet_1_0__leaf_net434),
    .X(net447));
 sky130_fd_sc_hd__or4bb_1 c542 (.A(clknet_1_0__leaf_net447),
    .B(clknet_1_0__leaf_net442),
    .C_N(clknet_1_0__leaf_net444),
    .D_N(clknet_1_0__leaf_net435),
    .X(net448));
 sky130_fd_sc_hd__a2111o_1 c543 (.A1(clknet_1_1__leaf_net444),
    .A2(clknet_1_1__leaf_net435),
    .B1(clknet_1_0__leaf_net439),
    .C1(clknet_1_0__leaf_net442),
    .D1(clknet_1_0__leaf_net438),
    .X(net449));
 sky130_fd_sc_hd__a2111o_1 c544 (.A1(clknet_1_1__leaf_net449),
    .A2(clknet_1_1__leaf_net442),
    .B1(clknet_1_1__leaf_net444),
    .C1(clknet_1_1__leaf_net437),
    .D1(net715),
    .X(net450));
 sky130_fd_sc_hd__mux4_1 c545 (.A0(clknet_1_0__leaf_net450),
    .A1(clknet_1_0__leaf_net449),
    .A2(clknet_1_1__leaf_net444),
    .A3(clknet_1_1__leaf_net440),
    .S0(clknet_1_1__leaf_net435),
    .S1(clknet_1_0__leaf_net442),
    .X(net451));
 sky130_fd_sc_hd__mux4_1 c546 (.A0(clknet_1_1__leaf_net443),
    .A1(clknet_1_1__leaf_net445),
    .A2(clknet_1_0__leaf_net450),
    .A3(clknet_1_0__leaf_net449),
    .S0(clknet_1_1__leaf_net442),
    .S1(net796),
    .X(net452));
 sky130_fd_sc_hd__mux4_1 c547 (.A0(clknet_1_0__leaf_net446),
    .A1(clknet_1_1__leaf_net447),
    .A2(clknet_1_1__leaf_net450),
    .A3(net714),
    .S0(net796),
    .S1(net797),
    .X(net453));
 sky130_fd_sc_hd__mux4_1 c548 (.A0(clknet_1_1__leaf_net438),
    .A1(clknet_1_1__leaf_net444),
    .A2(clknet_1_1__leaf_net442),
    .A3(net796),
    .S0(net797),
    .S1(net933),
    .X(net454));
 sky130_fd_sc_hd__mux4_1 c549 (.A0(net454),
    .A1(clknet_1_1__leaf_net446),
    .A2(clknet_1_0__leaf_net444),
    .A3(clknet_1_1__leaf_net442),
    .S0(net796),
    .S1(net797),
    .X(net455));
 sky130_fd_sc_hd__and2_1 c550 (.A(net715),
    .B(net933),
    .X(net456));
 sky130_fd_sc_hd__and2_1 c551 (.A(net456),
    .B(net933),
    .X(net457));
 sky130_fd_sc_hd__and2_1 c552 (.A(net457),
    .B(net456),
    .X(net458));
 sky130_fd_sc_hd__and3_1 c553 (.A(net456),
    .B(net457),
    .C(net933),
    .X(net459));
 sky130_fd_sc_hd__or4bb_1 c554 (.A(net458),
    .B(net459),
    .C_N(net457),
    .D_N(clknet_1_1__leaf_net359),
    .X(net460));
 sky130_fd_sc_hd__and2_0 c555 (.A(net458),
    .B(clknet_1_0__leaf_net460),
    .X(net461));
 sky130_fd_sc_hd__and3_1 c556 (.A(clknet_1_0__leaf_net461),
    .B(net459),
    .C(net456),
    .X(net462));
 sky130_fd_sc_hd__and3_1 c557 (.A(net459),
    .B(clknet_1_0__leaf_net460),
    .C(clknet_1_0__leaf_net461),
    .X(net463));
 sky130_fd_sc_hd__sdfbbp_1 c558 (.CLK(clknet_4_5_0_clk),
    .D(clknet_1_0__leaf_net463),
    .RESET_B(clknet_1_0__leaf_net461),
    .SCD(clknet_1_0__leaf_net460),
    .SCE(net456),
    .SET_B(clknet_1_1__leaf_net359),
    .Q(net465),
    .Q_N(net464));
 sky130_fd_sc_hd__a2111o_1 c559 (.A1(clknet_1_1__leaf_net359),
    .A2(net465),
    .B1(clknet_1_0__leaf_net462),
    .C1(net457),
    .D1(net459),
    .X(net466));
 sky130_fd_sc_hd__and3_1 c560 (.A(clknet_1_1__leaf_net460),
    .B(clknet_1_1__leaf_net461),
    .C(net722),
    .X(net467));
 sky130_fd_sc_hd__buf_1 c561 (.A(clknet_1_0__leaf_net827),
    .X(net468));
 sky130_fd_sc_hd__mux4_1 c562 (.A0(clknet_1_1__leaf_net463),
    .A1(net458),
    .A2(clknet_1_1__leaf_net461),
    .A3(clknet_1_1__leaf_net460),
    .S0(clknet_1_1__leaf_net467),
    .S1(clknet_1_0__leaf_net359),
    .X(net469));
 sky130_fd_sc_hd__sdfbbn_1 c563 (.CLK_N(clknet_4_4_0_clk),
    .D(net457),
    .RESET_B(clknet_1_0__leaf_net467),
    .SCD(net458),
    .SCE(clknet_1_0__leaf_net463),
    .SET_B(clknet_1_0__leaf_net468),
    .Q(net471),
    .Q_N(net470));
 sky130_fd_sc_hd__sedfxbp_1 c564 (.CLK(clknet_4_5_0_clk),
    .D(net471),
    .DE(clknet_1_0__leaf_net467),
    .SCD(clknet_1_0__leaf_net460),
    .SCE(clknet_1_0__leaf_net468),
    .Q(net473),
    .Q_N(net472));
 sky130_fd_sc_hd__sdfbbn_1 c565 (.CLK_N(clknet_4_6_0_clk),
    .D(net473),
    .RESET_B(clknet_1_1__leaf_net468),
    .SCD(clknet_1_1__leaf_net467),
    .SCE(clknet_1_1__leaf_net461),
    .SET_B(net944),
    .Q(net475),
    .Q_N(net474));
 sky130_fd_sc_hd__sdfbbp_1 c566 (.CLK(clknet_4_5_0_clk),
    .D(clknet_1_0__leaf_net468),
    .RESET_B(net473),
    .SCD(net475),
    .SCE(clknet_1_0__leaf_net460),
    .SET_B(clknet_1_0__leaf_net467),
    .Q(net477),
    .Q_N(net476));
 sky130_fd_sc_hd__mux4_1 c567 (.A0(clknet_1_1__leaf_net363),
    .A1(net477),
    .A2(net470),
    .A3(net456),
    .S0(clknet_1_0__leaf_net468),
    .S1(net944),
    .X(net478));
 sky130_fd_sc_hd__mux4_1 c568 (.A0(net465),
    .A1(net458),
    .A2(clknet_1_1__leaf_net467),
    .A3(clknet_1_1__leaf_net463),
    .S0(net722),
    .S1(net800),
    .X(net479));
 sky130_fd_sc_hd__mux4_1 c569 (.A0(net471),
    .A1(net476),
    .A2(net458),
    .A3(net472),
    .S0(net722),
    .S1(net802),
    .X(net480));
 sky130_fd_sc_hd__mux4_1 c570 (.A0(clknet_1_1__leaf_net462),
    .A1(net480),
    .A2(clknet_1_0__leaf_net467),
    .A3(net470),
    .S0(net476),
    .S1(net722),
    .X(net481));
 sky130_fd_sc_hd__mux4_1 c571 (.A0(net477),
    .A1(clknet_1_1__leaf_net467),
    .A2(net480),
    .A3(clknet_1_1__leaf_net460),
    .S0(clknet_1_1__leaf_net788),
    .S1(net803),
    .X(net482));
 sky130_fd_sc_hd__clkbuf_1 c572 (.A(net704),
    .X(net483));
 sky130_fd_sc_hd__buf_1 c573 (.A(net704),
    .X(net484));
 sky130_fd_sc_hd__and2_1 c574 (.A(net484),
    .B(net803),
    .X(net485));
 sky130_fd_sc_hd__and2_2 c575 (.A(net485),
    .B(net484),
    .X(net486));
 sky130_fd_sc_hd__and2_1 c576 (.A(net486),
    .B(net800),
    .X(net487));
 sky130_fd_sc_hd__buf_1 c577 (.A(net830),
    .X(net488));
 sky130_fd_sc_hd__and3_1 c578 (.A(net486),
    .B(net487),
    .C(net795),
    .X(net489));
 sky130_fd_sc_hd__and2_0 c579 (.A(net487),
    .B(net489),
    .X(net490));
 sky130_fd_sc_hd__and3_1 c580 (.A(net484),
    .B(net485),
    .C(net486),
    .X(net491));
 sky130_fd_sc_hd__or4bb_2 c581 (.A(net489),
    .B(net485),
    .C_N(net488),
    .D_N(net804),
    .X(net492));
 sky130_fd_sc_hd__and3_1 c582 (.A(net486),
    .B(net489),
    .C(net491),
    .X(net493));
 sky130_fd_sc_hd__or4bb_2 c583 (.A(net493),
    .B(net485),
    .C_N(net486),
    .D_N(net492),
    .X(net494));
 sky130_fd_sc_hd__and3_1 c584 (.A(net489),
    .B(net492),
    .C(net494),
    .X(net495));
 sky130_fd_sc_hd__and3_1 c585 (.A(net488),
    .B(net486),
    .C(net490),
    .X(net496));
 sky130_fd_sc_hd__and3_1 c586 (.A(net494),
    .B(net488),
    .C(net495),
    .X(net497));
 sky130_fd_sc_hd__mux4_1 c587 (.A0(net491),
    .A1(net488),
    .A2(net496),
    .A3(net486),
    .S0(net492),
    .S1(net484),
    .X(net498));
 sky130_fd_sc_hd__a2111o_1 c588 (.A1(net498),
    .A2(net491),
    .B1(net494),
    .C1(net496),
    .D1(clknet_1_1__leaf_net270),
    .X(net499));
 sky130_fd_sc_hd__mux4_1 c589 (.A0(net483),
    .A1(net491),
    .A2(net484),
    .A3(net495),
    .S0(net494),
    .S1(net803),
    .X(net500));
 sky130_fd_sc_hd__or4bb_1 c590 (.A(net495),
    .B(net496),
    .C_N(net498),
    .D_N(net704),
    .X(net501));
 sky130_fd_sc_hd__mux4_1 c591 (.A0(net501),
    .A1(net492),
    .A2(net495),
    .A3(net498),
    .S0(net489),
    .S1(net486),
    .X(net502));
 sky130_fd_sc_hd__mux4_1 c592 (.A0(net497),
    .A1(net496),
    .A2(net501),
    .A3(net502),
    .S0(net486),
    .S1(net487),
    .X(net503));
 sky130_fd_sc_hd__mux4_1 c593 (.A0(net492),
    .A1(net502),
    .A2(net495),
    .A3(net494),
    .S0(net501),
    .S1(net798),
    .X(net504));
 sky130_fd_sc_hd__clkbuf_2 c594 (.A(net680),
    .X(net505));
 sky130_fd_sc_hd__and2_1 c595 (.A(net505),
    .B(net283),
    .X(net506));
 sky130_fd_sc_hd__and3_1 c596 (.A(net500),
    .B(net505),
    .C(net917),
    .X(net507));
 sky130_fd_sc_hd__and3_1 c597 (.A(net507),
    .B(net917),
    .C(net729),
    .X(net508));
 sky130_fd_sc_hd__and2_1 c598 (.A(net508),
    .B(net917),
    .X(net509));
 sky130_fd_sc_hd__clkbuf_1 c599 (.A(net679),
    .X(net510));
 sky130_fd_sc_hd__or4bb_2 c600 (.A(net509),
    .B(net507),
    .C_N(net505),
    .D_N(net917),
    .X(net511));
 sky130_fd_sc_hd__and3_2 c601 (.A(net510),
    .B(net505),
    .C(net511),
    .X(net512));
 sky130_fd_sc_hd__a2111o_2 c602 (.A1(net512),
    .A2(net505),
    .B1(net917),
    .C1(net511),
    .D1(net729),
    .X(net513));
 sky130_fd_sc_hd__sdfbbn_1 c603 (.CLK_N(clknet_4_12_0_clk),
    .D(net513),
    .RESET_B(net512),
    .SCD(net505),
    .SCE(clknet_1_1__leaf_net415),
    .SET_B(net917),
    .Q(net515),
    .Q_N(net514));
 sky130_fd_sc_hd__sdfbbn_1 c604 (.CLK_N(clknet_4_14_0_clk),
    .D(net511),
    .RESET_B(net513),
    .SCD(net515),
    .SCE(net512),
    .SET_B(net918),
    .Q(net517),
    .Q_N(net516));
 sky130_fd_sc_hd__mux4_1 c605 (.A0(net507),
    .A1(net512),
    .A2(net508),
    .A3(net505),
    .S0(net513),
    .S1(net917),
    .X(net518));
 sky130_fd_sc_hd__a2111o_2 c606 (.A1(net505),
    .A2(net517),
    .B1(net515),
    .C1(net512),
    .D1(net918),
    .X(net519));
 sky130_fd_sc_hd__a2111o_1 c607 (.A1(net512),
    .A2(net511),
    .B1(net508),
    .C1(net519),
    .D1(net948),
    .X(net520));
 sky130_fd_sc_hd__sdfbbp_1 c608 (.CLK(clknet_4_13_0_clk),
    .D(net519),
    .RESET_B(net514),
    .SCD(net512),
    .SCE(net712),
    .SET_B(net948),
    .Q(net522),
    .Q_N(net521));
 sky130_fd_sc_hd__sdfbbn_1 c609 (.CLK_N(clknet_4_12_0_clk),
    .D(net508),
    .RESET_B(net522),
    .SCD(net512),
    .SCE(net519),
    .SET_B(net513),
    .Q(net524),
    .Q_N(net523));
 sky130_fd_sc_hd__mux4_1 c610 (.A0(net517),
    .A1(net522),
    .A2(net513),
    .A3(net519),
    .S0(net512),
    .S1(net523),
    .X(net525));
 sky130_fd_sc_hd__sdfbbn_1 c611 (.CLK_N(clknet_4_15_0_clk),
    .D(net955),
    .RESET_B(net519),
    .SCD(net521),
    .SCE(net729),
    .SET_B(clknet_1_0__leaf_net806),
    .Q(net527),
    .Q_N(net526));
 sky130_fd_sc_hd__mux4_1 c612 (.A0(net526),
    .A1(net511),
    .A2(net505),
    .A3(net509),
    .S0(net524),
    .S1(clknet_1_1__leaf_net806),
    .X(net528));
 sky130_fd_sc_hd__mux4_1 c613 (.A0(net527),
    .A1(clknet_1_0__leaf_net528),
    .A2(net918),
    .A3(net516),
    .S0(net519),
    .S1(clknet_1_0__leaf_net806),
    .X(net529));
 sky130_fd_sc_hd__mux4_1 c614 (.A0(clknet_1_0__leaf_net528),
    .A1(net511),
    .A2(net712),
    .A3(net805),
    .S0(clknet_1_1__leaf_net806),
    .S1(clknet_1_0__leaf_net807),
    .X(net530));
 sky130_fd_sc_hd__mux4_1 c615 (.A0(net509),
    .A1(net530),
    .A2(clknet_1_1__leaf_net528),
    .A3(net511),
    .S0(clknet_1_1__leaf_net806),
    .S1(clknet_1_1__leaf_net807),
    .X(net531));
 sky130_fd_sc_hd__and3_2 c616 (.A(net900),
    .B(net918),
    .C(net908),
    .X(net896));
 sky130_fd_sc_hd__and3_1 c617 (.A(net504),
    .B(net712),
    .C(net902),
    .X(net893));
 sky130_fd_sc_hd__and2_2 c618 (.A(net893),
    .B(net918),
    .X(net894));
 sky130_fd_sc_hd__and3_2 c619 (.A(net893),
    .B(net515),
    .C(net894),
    .X(net532));
 sky130_fd_sc_hd__mux4_1 c62 (.A0(net879),
    .A1(net878),
    .A2(net872),
    .A3(net877),
    .S0(net875),
    .S1(net881),
    .X(net0));
 sky130_fd_sc_hd__or4bb_1 c620 (.A(net532),
    .B(net893),
    .C_N(net894),
    .D_N(net514),
    .X(net897));
 sky130_fd_sc_hd__and3_2 c621 (.A(net897),
    .B(net896),
    .C(net899),
    .X(net898));
 sky130_fd_sc_hd__sedfxtp_2 c622 (.CLK(clknet_4_15_0_clk),
    .D(net898),
    .DE(net532),
    .SCD(net893),
    .SCE(net918),
    .Q(net533));
 sky130_fd_sc_hd__or4bb_1 c623 (.A(net934),
    .B(net532),
    .C_N(net894),
    .D_N(net902),
    .X(net534));
 sky130_fd_sc_hd__or4bb_2 c624 (.A(net897),
    .B(net534),
    .C_N(net896),
    .D_N(net934),
    .X(net535));
 sky130_fd_sc_hd__a2111o_1 c625 (.A1(net532),
    .A2(net535),
    .B1(net934),
    .C1(net898),
    .D1(net896),
    .X(net536));
 sky130_fd_sc_hd__sdfbbp_1 c626 (.CLK(clknet_4_15_0_clk),
    .D(net534),
    .RESET_B(net896),
    .SCD(net532),
    .SCE(net898),
    .SET_B(net958),
    .Q(net538),
    .Q_N(net537));
 sky130_fd_sc_hd__a2111o_1 c627 (.A1(net533),
    .A2(net532),
    .B1(net537),
    .C1(net894),
    .D1(net711),
    .X(net539));
 sky130_fd_sc_hd__mux4_1 c628 (.A0(net894),
    .A1(net534),
    .A2(net539),
    .A3(net535),
    .S0(net934),
    .S1(net704),
    .X(net540));
 sky130_fd_sc_hd__a2111o_1 c629 (.A1(net896),
    .A2(net934),
    .B1(net894),
    .C1(net539),
    .D1(clknet_1_0__leaf_net808),
    .X(net541));
 sky130_fd_sc_hd__mux4_1 c63 (.A0(net888),
    .A1(net886),
    .A2(net883),
    .A3(net885),
    .S0(net0),
    .S1(net875),
    .X(net1));
 sky130_fd_sc_hd__mux4_1 c630 (.A0(net539),
    .A1(net538),
    .A2(clknet_1_0__leaf_net541),
    .A3(net934),
    .S0(net894),
    .S1(clknet_1_0__leaf_net808),
    .X(net542));
 sky130_fd_sc_hd__mux4_1 c631 (.A0(net539),
    .A1(net934),
    .A2(net894),
    .A3(net535),
    .S0(clknet_1_0__leaf_net808),
    .S1(net895),
    .X(net543));
 sky130_fd_sc_hd__mux4_1 c632 (.A0(net538),
    .A1(clknet_1_1__leaf_net541),
    .A2(net535),
    .A3(net539),
    .S0(net533),
    .S1(net810),
    .X(net544));
 sky130_fd_sc_hd__mux4_1 c633 (.A0(net898),
    .A1(net515),
    .A2(net934),
    .A3(clknet_1_1__leaf_net808),
    .S0(net810),
    .S1(net811),
    .X(net545));
 sky130_fd_sc_hd__mux4_1 c634 (.A0(net535),
    .A1(clknet_1_1__leaf_net401),
    .A2(clknet_1_0__leaf_net541),
    .A3(net934),
    .S0(clknet_1_0__leaf_net808),
    .S1(net810),
    .X(net546));
 sky130_fd_sc_hd__mux4_1 c635 (.A0(net897),
    .A1(net533),
    .A2(net532),
    .A3(net534),
    .S0(net813),
    .S1(net950),
    .X(net547));
 sky130_fd_sc_hd__mux4_1 c636 (.A0(net515),
    .A1(net547),
    .A2(clknet_1_1__leaf_net541),
    .A3(net809),
    .S0(net812),
    .S1(net813),
    .X(net548));
 sky130_fd_sc_hd__sdfbbn_1 c637 (.CLK_N(clknet_4_14_0_clk),
    .D(net547),
    .RESET_B(net898),
    .SCD(net711),
    .SCE(net967),
    .SET_B(net950),
    .Q(net914),
    .Q_N(net905));
 sky130_fd_sc_hd__mux4_1 c64 (.A0(net873),
    .A1(net880),
    .A2(net3),
    .A3(net1),
    .S0(net874),
    .S1(net882),
    .X(net2));
 sky130_fd_sc_hd__mux4_1 c65 (.A0(net863),
    .A1(net852),
    .A2(net857),
    .A3(net858),
    .S0(net849),
    .S1(net868),
    .X(net3));
 sky130_fd_sc_hd__and2_1 c66 (.A(net889),
    .B(net871),
    .X(net4));
 sky130_fd_sc_hd__and2_0 c660 (.A(clknet_1_1__leaf_net788),
    .B(net933),
    .X(net549));
 sky130_fd_sc_hd__and2_0 c661 (.A(clknet_1_0__leaf_net549),
    .B(net933),
    .X(net550));
 sky130_fd_sc_hd__and2_0 c662 (.A(clknet_1_0__leaf_net550),
    .B(clknet_1_0__leaf_net549),
    .X(net551));
 sky130_fd_sc_hd__and2_0 c663 (.A(clknet_1_0__leaf_net549),
    .B(net933),
    .X(net552));
 sky130_fd_sc_hd__and3_1 c664 (.A(clknet_1_0__leaf_net550),
    .B(net324),
    .C(net933),
    .X(net553));
 sky130_fd_sc_hd__and2_0 c665 (.A(clknet_1_0__leaf_net553),
    .B(clknet_1_0__leaf_net552),
    .X(net554));
 sky130_fd_sc_hd__and3_1 c666 (.A(clknet_1_0__leaf_net554),
    .B(clknet_1_0__leaf_net551),
    .C(clknet_1_1__leaf_net549),
    .X(net555));
 sky130_fd_sc_hd__and2_0 c667 (.A(clknet_1_0__leaf_net555),
    .B(clknet_1_1__leaf_net553),
    .X(net556));
 sky130_fd_sc_hd__and2_0 c668 (.A(clknet_1_0__leaf_net556),
    .B(clknet_1_1__leaf_net550),
    .X(net557));
 sky130_fd_sc_hd__and2_0 c669 (.A(clknet_1_1__leaf_net553),
    .B(clknet_1_0__leaf_net557),
    .X(net558));
 sky130_fd_sc_hd__and2_1 c67 (.A(net870),
    .B(net4),
    .X(net5));
 sky130_fd_sc_hd__and3_1 c670 (.A(clknet_1_0__leaf_net554),
    .B(clknet_1_1__leaf_net558),
    .C(clknet_1_0__leaf_net556),
    .X(net559));
 sky130_fd_sc_hd__and3_1 c671 (.A(clknet_1_1__leaf_net556),
    .B(clknet_1_1__leaf_net554),
    .C(clknet_1_0__leaf_net557),
    .X(net560));
 sky130_fd_sc_hd__and3_1 c672 (.A(clknet_1_1__leaf_net552),
    .B(clknet_1_0__leaf_net558),
    .C(clknet_1_0__leaf_net553),
    .X(net561));
 sky130_fd_sc_hd__and3_1 c673 (.A(clknet_1_1__leaf_net551),
    .B(clknet_1_0__leaf_net555),
    .C(clknet_1_0__leaf_net554),
    .X(net562));
 sky130_fd_sc_hd__a2111o_1 c674 (.A1(clknet_1_0__leaf_net560),
    .A2(clknet_1_0__leaf_net562),
    .B1(clknet_1_1__leaf_net554),
    .C1(clknet_1_0__leaf_net559),
    .D1(clknet_1_1__leaf_net555),
    .X(net563));
 sky130_fd_sc_hd__buf_1 c675 (.A(net831),
    .X(net564));
 sky130_fd_sc_hd__mux4_1 c676 (.A0(clknet_1_0__leaf_net563),
    .A1(clknet_1_1__leaf_net555),
    .A2(net564),
    .A3(clknet_1_0__leaf_net562),
    .S0(clknet_1_0__leaf_net561),
    .S1(clknet_1_1__leaf_net556),
    .X(net565));
 sky130_fd_sc_hd__and3_1 c677 (.A(net564),
    .B(clknet_1_1__leaf_net562),
    .C(net815),
    .X(net566));
 sky130_fd_sc_hd__mux4_1 c678 (.A0(clknet_1_1__leaf_net562),
    .A1(clknet_1_0__leaf_net566),
    .A2(clknet_1_0__leaf_net561),
    .A3(clknet_1_1__leaf_net557),
    .S0(clknet_1_1__leaf_net554),
    .S1(clknet_1_1__leaf_net549),
    .X(net567));
 sky130_fd_sc_hd__mux4_1 c679 (.A0(clknet_1_1__leaf_net549),
    .A1(clknet_1_0__leaf_net567),
    .A2(clknet_1_1__leaf_net560),
    .A3(clknet_1_1__leaf_net566),
    .S0(clknet_1_1__leaf_net561),
    .S1(net815),
    .X(net568));
 sky130_fd_sc_hd__and2_1 c68 (.A(net4),
    .B(net5),
    .X(net6));
 sky130_fd_sc_hd__mux4_1 c680 (.A0(clknet_1_1__leaf_net559),
    .A1(clknet_1_0__leaf_net566),
    .A2(clknet_1_1__leaf_net567),
    .A3(net564),
    .S0(net753),
    .S1(net815),
    .X(net569));
 sky130_fd_sc_hd__mux4_1 c681 (.A0(clknet_1_1__leaf_net561),
    .A1(clknet_1_0__leaf_net567),
    .A2(clknet_1_0__leaf_net560),
    .A3(clknet_1_1__leaf_net557),
    .S1(net753),
    .X(net570));
 sky130_fd_sc_hd__and2_2 c682 (.A(net475),
    .B(net698),
    .X(net571));
 sky130_fd_sc_hd__and2_0 c683 (.A(net571),
    .B(clknet_1_1__leaf_net359),
    .X(net572));
 sky130_fd_sc_hd__and3_1 c684 (.A(clknet_1_0__leaf_net572),
    .B(net571),
    .C(net475),
    .X(net573));
 sky130_fd_sc_hd__and3_1 c685 (.A(clknet_1_0__leaf_net573),
    .B(clknet_1_0__leaf_net572),
    .C(net571),
    .X(net574));
 sky130_fd_sc_hd__and2_0 c686 (.A(clknet_1_0__leaf_net572),
    .B(clknet_1_0__leaf_net573),
    .X(net575));
 sky130_fd_sc_hd__and3_1 c687 (.A(clknet_1_0__leaf_net572),
    .B(net571),
    .C(net804),
    .X(net576));
 sky130_fd_sc_hd__buf_1 c688 (.A(net672),
    .X(net577));
 sky130_fd_sc_hd__or4bb_1 c689 (.A(net571),
    .B(net577),
    .C_N(clknet_1_0__leaf_net572),
    .D_N(clknet_1_0__leaf_net575),
    .X(net578));
 sky130_fd_sc_hd__and2_0 c69 (.A(net5),
    .B(net861),
    .X(net7));
 sky130_fd_sc_hd__buf_1 c690 (.A(net671),
    .X(net579));
 sky130_fd_sc_hd__dlymetal6s2s_1 c691 (.X(net580));
 sky130_fd_sc_hd__buf_1 c692 (.A(net691),
    .X(net581));
 sky130_fd_sc_hd__sdfbbn_1 c693 (.CLK_N(clknet_4_7_0_clk),
    .D(net580),
    .RESET_B(clknet_1_0__leaf_net575),
    .SCD(net581),
    .SCE(net571),
    .SET_B(clknet_1_1__leaf_net572),
    .Q(net583),
    .Q_N(net582));
 sky130_fd_sc_hd__and3_1 c694 (.A(net571),
    .B(net580),
    .C(net579),
    .X(net584));
 sky130_fd_sc_hd__sdfbbp_1 c695 (.CLK(clknet_4_7_0_clk),
    .D(clknet_1_1__leaf_net574),
    .RESET_B(net584),
    .SCD(net580),
    .SCE(net579),
    .SET_B(clknet_1_0__leaf_net575),
    .Q(net586),
    .Q_N(net585));
 sky130_fd_sc_hd__and3_1 c696 (.A(net583),
    .B(net586),
    .C(net584),
    .X(net587));
 sky130_fd_sc_hd__and3_1 c697 (.A(net579),
    .B(net586),
    .C(net581),
    .X(net588));
 sky130_fd_sc_hd__mux4_1 c698 (.A0(net588),
    .A1(net582),
    .A2(net580),
    .A3(clknet_1_1__leaf_net572),
    .S0(net585),
    .S1(net571),
    .X(net589));
 sky130_fd_sc_hd__mux4_1 c699 (.A0(net587),
    .A1(net588),
    .A2(net580),
    .A3(net579),
    .S0(clknet_1_0__leaf_net589),
    .S1(net734),
    .X(net590));
 sky130_fd_sc_hd__and3_1 c70 (.A(net884),
    .B(net6),
    .C(net5),
    .X(net8));
 sky130_fd_sc_hd__mux4_1 c700 (.A0(clknet_1_1__leaf_net576),
    .A1(clknet_1_0__leaf_net589),
    .A2(net586),
    .A3(net580),
    .S0(net734),
    .S1(net815),
    .X(net591));
 sky130_fd_sc_hd__mux4_1 c701 (.A0(clknet_1_0__leaf_net590),
    .A1(net588),
    .A2(clknet_1_1__leaf_net591),
    .A3(net580),
    .S0(net585),
    .S1(net815),
    .X(net592));
 sky130_fd_sc_hd__mux4_1 c702 (.A0(clknet_1_0__leaf_net591),
    .A1(net581),
    .A2(clknet_1_1__leaf_net589),
    .A3(clknet_1_1__leaf_net590),
    .S0(net585),
    .S1(net816),
    .X(net593));
 sky130_fd_sc_hd__mux4_1 c703 (.A0(net584),
    .A1(net587),
    .A2(clknet_1_0__leaf_net591),
    .A3(net579),
    .S0(net734),
    .S1(net816),
    .X(net594));
 sky130_fd_sc_hd__and2_1 c704 (.A(net490),
    .B(net803),
    .X(net595));
 sky130_fd_sc_hd__dlymetal6s2s_1 c705 (.A(net670),
    .X(net596));
 sky130_fd_sc_hd__buf_1 c706 (.A(clknet_1_1__leaf_net827),
    .X(net597));
 sky130_fd_sc_hd__clkbuf_1 c707 (.A(net670),
    .X(net598));
 sky130_fd_sc_hd__and2_2 c708 (.A(net596),
    .B(net598),
    .X(net599));
 sky130_fd_sc_hd__and3_1 c709 (.A(clknet_1_0__leaf_net597),
    .B(net596),
    .C(net798),
    .X(net600));
 sky130_fd_sc_hd__and3_1 c71 (.A(net6),
    .B(net4),
    .C(net929),
    .X(net9));
 sky130_fd_sc_hd__sdfbbn_1 c710 (.CLK_N(clknet_4_7_0_clk),
    .D(net577),
    .RESET_B(clknet_1_1__leaf_net575),
    .SCD(net599),
    .SCE(net933),
    .SET_B(net817),
    .Q(net602),
    .Q_N(net601));
 sky130_fd_sc_hd__and3_1 c711 (.A(net503),
    .B(net602),
    .C(clknet_1_1__leaf_net600),
    .X(net603));
 sky130_fd_sc_hd__and3_1 c712 (.A(clknet_1_0__leaf_net603),
    .B(net596),
    .C(net474),
    .X(net604));
 sky130_fd_sc_hd__and2_0 c713 (.A(clknet_1_0__leaf_net597),
    .B(clknet_1_0__leaf_net600),
    .X(net605));
 sky130_fd_sc_hd__and3_1 c714 (.A(clknet_1_0__leaf_net604),
    .B(net601),
    .C(net599),
    .X(net606));
 sky130_fd_sc_hd__a2111o_1 c715 (.A1(net605),
    .A2(net595),
    .B1(clknet_1_0__leaf_net606),
    .C1(net599),
    .D1(net601),
    .X(net607));
 sky130_fd_sc_hd__mux4_1 c716 (.A0(clknet_1_0__leaf_net604),
    .A1(clknet_1_0__leaf_net606),
    .A2(net595),
    .A3(clknet_1_0__leaf_net607),
    .S0(net577),
    .S1(net817),
    .X(net608));
 sky130_fd_sc_hd__and3_1 c717 (.A(clknet_1_0__leaf_net606),
    .B(clknet_1_1__leaf_net607),
    .C(net599),
    .X(net609));
 sky130_fd_sc_hd__sdfbbn_1 c718 (.CLK_N(clknet_4_13_0_clk),
    .D(clknet_1_1__leaf_net608),
    .RESET_B(net599),
    .SCD(clknet_1_0__leaf_net609),
    .SCE(clknet_1_1__leaf_net604),
    .SET_B(clknet_1_1__leaf_net606),
    .Q(net611),
    .Q_N(net610));
 sky130_fd_sc_hd__sdfbbp_1 c719 (.CLK(clknet_4_13_0_clk),
    .D(clknet_1_1__leaf_net607),
    .RESET_B(clknet_1_1__leaf_net608),
    .SCD(net610),
    .SCE(clknet_1_1__leaf_net609),
    .SET_B(net599),
    .Q(net613),
    .Q_N(net612));
 sky130_fd_sc_hd__and3_2 c72 (.A(net6),
    .B(net9),
    .C(net929),
    .X(net10));
 sky130_fd_sc_hd__sdfbbn_1 c720 (.CLK_N(clknet_4_13_0_clk),
    .D(clknet_1_0__leaf_net600),
    .RESET_B(net611),
    .SCD(clknet_1_0__leaf_net606),
    .SCE(clknet_1_0__leaf_net607),
    .SET_B(clknet_1_1__leaf_net373),
    .Q(net615),
    .Q_N(net614));
 sky130_fd_sc_hd__a2111o_1 c721 (.A1(net615),
    .A2(clknet_1_1__leaf_net606),
    .B1(net611),
    .C1(clknet_1_0__leaf_net608),
    .D1(clknet_1_0__leaf_net609),
    .X(net616));
 sky130_fd_sc_hd__mux4_1 c722 (.A0(net602),
    .A1(clknet_1_1__leaf_net603),
    .A2(clknet_1_0__leaf_net608),
    .A3(net599),
    .S0(clknet_1_1__leaf_net606),
    .S1(net615),
    .X(net617));
 sky130_fd_sc_hd__mux4_1 c723 (.A0(clknet_1_1__leaf_net609),
    .A1(net611),
    .A2(net613),
    .A3(clknet_1_1__leaf_net604),
    .S0(clknet_1_1__leaf_net606),
    .S1(net818),
    .X(net618));
 sky130_fd_sc_hd__a2111o_1 c724 (.A1(net612),
    .A2(clknet_1_1__leaf_net597),
    .B1(net610),
    .C1(net753),
    .D1(net819),
    .X(net619));
 sky130_fd_sc_hd__mux4_1 c725 (.A0(net613),
    .A1(net619),
    .A2(net614),
    .A3(net610),
    .S0(net753),
    .S1(net819),
    .X(net620));
 sky130_fd_sc_hd__and2_0 c726 (.A(net620),
    .B(net514),
    .X(net621));
 sky130_fd_sc_hd__and2_0 c727 (.A(clknet_1_0__leaf_net621),
    .B(net599),
    .X(net622));
 sky130_fd_sc_hd__and3_1 c728 (.A(clknet_1_1__leaf_net622),
    .B(clknet_1_1__leaf_net621),
    .C(net917),
    .X(net623));
 sky130_fd_sc_hd__and2_0 c729 (.A(clknet_1_0__leaf_net622),
    .B(clknet_1_0__leaf_net623),
    .X(net624));
 sky130_fd_sc_hd__or4bb_2 c73 (.A(net9),
    .B(net6),
    .C_N(net10),
    .D_N(net929),
    .X(net11));
 sky130_fd_sc_hd__and3_1 c730 (.A(net917),
    .B(clknet_1_0__leaf_net624),
    .C(clknet_1_0__leaf_net621),
    .X(net625));
 sky130_fd_sc_hd__and2_0 c731 (.A(clknet_1_0__leaf_net623),
    .B(clknet_1_0__leaf_net624),
    .X(net626));
 sky130_fd_sc_hd__sdfbbn_1 c732 (.CLK_N(clknet_4_12_0_clk),
    .D(clknet_1_1__leaf_net625),
    .RESET_B(clknet_1_1__leaf_net626),
    .SCD(clknet_1_0__leaf_net624),
    .SCE(clknet_1_1__leaf_net575),
    .SET_B(clknet_1_0__leaf_net401),
    .Q(net628),
    .Q_N(net627));
 sky130_fd_sc_hd__or4bb_1 c733 (.A(clknet_1_1__leaf_net622),
    .B(net627),
    .C_N(clknet_1_1__leaf_net623),
    .D_N(net598),
    .X(net629));
 sky130_fd_sc_hd__mux4_1 c734 (.A0(net598),
    .A1(clknet_1_1__leaf_net622),
    .A2(clknet_1_1__leaf_net629),
    .A3(net627),
    .S0(clknet_1_1__leaf_net626),
    .S1(net729),
    .X(net630));
 sky130_fd_sc_hd__and3_1 c735 (.A(clknet_1_1__leaf_net624),
    .B(clknet_1_0__leaf_net629),
    .C(clknet_1_0__leaf_net626),
    .X(net631));
 sky130_fd_sc_hd__mux4_1 c736 (.A0(clknet_1_0__leaf_net626),
    .A1(net628),
    .A2(clknet_1_1__leaf_net630),
    .A3(net514),
    .S0(clknet_1_1__leaf_net624),
    .S1(clknet_1_1__leaf_net629),
    .X(net632));
 sky130_fd_sc_hd__and3_1 c737 (.A(clknet_1_1__leaf_net632),
    .B(clknet_1_0__leaf_net622),
    .C(clknet_1_1__leaf_net623),
    .X(net633));
 sky130_fd_sc_hd__or4bb_1 c738 (.A(clknet_1_0__leaf_net630),
    .B(clknet_1_1__leaf_net631),
    .C_N(clknet_1_1__leaf_net624),
    .D_N(clknet_1_1__leaf_net629),
    .X(net634));
 sky130_fd_sc_hd__mux4_1 c739 (.A0(net628),
    .A1(clknet_1_1__leaf_net626),
    .A2(clknet_1_1__leaf_net631),
    .A3(clknet_1_1__leaf_net634),
    .S0(clknet_1_1__leaf_net629),
    .S1(clknet_1_1__leaf_net622),
    .X(net635));
 sky130_fd_sc_hd__and3_1 c74 (.A(net10),
    .B(net11),
    .C(net9),
    .X(net12));
 sky130_fd_sc_hd__mux4_1 c740 (.A0(clknet_1_0__leaf_net629),
    .A1(clknet_1_1__leaf_net631),
    .A2(clknet_1_0__leaf_net632),
    .A3(clknet_1_0__leaf_net634),
    .S0(clknet_1_0__leaf_net625),
    .S1(clknet_1_1__leaf_net626),
    .X(net636));
 sky130_fd_sc_hd__clkbuf_1 c741 (.A(net833),
    .X(net637));
 sky130_fd_sc_hd__mux4_1 c742 (.A0(clknet_1_0__leaf_net636),
    .A1(clknet_1_0__leaf_net634),
    .A2(net637),
    .A3(clknet_1_1__leaf_net626),
    .S0(clknet_1_0__leaf_net624),
    .S1(clknet_1_0__leaf_net631),
    .X(net638));
 sky130_fd_sc_hd__sedfxtp_1 c743 (.CLK(clknet_4_9_0_clk),
    .D(clknet_1_0__leaf_net401),
    .DE(clknet_1_0__leaf_net634),
    .SCD(clknet_1_0__leaf_net636),
    .SCE(net965),
    .Q(net639));
 sky130_fd_sc_hd__mux4_1 c744 (.A0(net637),
    .A1(net639),
    .A2(clknet_1_1__leaf_net633),
    .A3(clknet_1_1__leaf_net636),
    .S0(clknet_1_0__leaf_net629),
    .S1(clknet_1_1__leaf_net634),
    .X(net640));
 sky130_fd_sc_hd__mux4_1 c745 (.A0(clknet_1_0__leaf_net633),
    .A1(clknet_1_1__leaf_net636),
    .A2(clknet_1_0__leaf_net631),
    .A3(clknet_1_0__leaf_net629),
    .S0(clknet_1_0__leaf_net626),
    .S1(net822),
    .X(net641));
 sky130_fd_sc_hd__a2111o_1 c746 (.A1(clknet_1_1__leaf_net634),
    .A2(net639),
    .B1(clknet_1_0__leaf_net636),
    .C1(net821),
    .D1(net822),
    .X(net642));
 sky130_fd_sc_hd__mux4_1 c747 (.A0(clknet_1_0__leaf_net631),
    .A1(clknet_1_1__leaf_net636),
    .A2(clknet_1_0__leaf_net622),
    .A3(clknet_1_1__leaf_net634),
    .S1(net823),
    .X(net703));
 sky130_fd_sc_hd__and3_1 c748 (.A(clknet_1_1__leaf_net621),
    .B(net904),
    .C(clknet_1_0__leaf_net626),
    .X(net644));
 sky130_fd_sc_hd__and2_0 c749 (.A(clknet_1_0__leaf_net644),
    .B(clknet_1_0__leaf_net626),
    .X(net645));
 sky130_fd_sc_hd__and3_2 c75 (.A(net7),
    .B(net9),
    .C(net11),
    .X(net13));
 sky130_fd_sc_hd__and3_1 c750 (.A(clknet_1_1__leaf_net644),
    .B(clknet_1_1__leaf_net645),
    .C(net895),
    .X(net646));
 sky130_fd_sc_hd__buf_1 c751 (.A(net757),
    .X(net647));
 sky130_fd_sc_hd__clkbuf_1 c752 (.A(net957),
    .X(net648));
 sky130_fd_sc_hd__dlymetal6s2s_1 c753 (.A(net756),
    .X(net649));
 sky130_fd_sc_hd__clkbuf_1 c754 (.A(net695),
    .X(net650));
 sky130_fd_sc_hd__and3_1 c755 (.A(net647),
    .B(clknet_1_1__leaf_net645),
    .C(net649),
    .X(net651));
 sky130_fd_sc_hd__buf_1 c756 (.A(net696),
    .X(net652));
 sky130_fd_sc_hd__buf_1 c757 (.A(clknet_1_1__leaf_net826),
    .X(net653));
 sky130_fd_sc_hd__buf_1 c758 (.A(clknet_1_0__leaf_net826),
    .X(net654));
 sky130_fd_sc_hd__a2111o_1 c759 (.A1(net650),
    .A2(net649),
    .B1(net647),
    .C1(net652),
    .D1(clknet_1_0__leaf_net645),
    .X(net655));
 sky130_fd_sc_hd__and3_2 c76 (.A(net4),
    .B(net2),
    .C(net13),
    .X(net14));
 sky130_fd_sc_hd__mux4_1 c760 (.A0(net652),
    .A1(clknet_1_1__leaf_net654),
    .A2(clknet_1_0__leaf_net645),
    .A3(clknet_1_1__leaf_net646),
    .S0(clknet_1_1__leaf_net655),
    .S1(net650),
    .X(net656));
 sky130_fd_sc_hd__sdfbbp_1 c761 (.CLK(clknet_4_11_0_clk),
    .D(clknet_1_0__leaf_net653),
    .RESET_B(clknet_1_0__leaf_net655),
    .SCD(net649),
    .SCE(clknet_1_0__leaf_net646),
    .SET_B(clknet_1_0__leaf_net654),
    .Q(net658),
    .Q_N(net657));
 sky130_fd_sc_hd__mux4_1 c762 (.A0(clknet_1_0__leaf_net653),
    .A1(net658),
    .A2(clknet_1_1__leaf_net646),
    .A3(net649),
    .S0(net652),
    .X(net659));
 sky130_fd_sc_hd__mux4_1 c763 (.A0(net658),
    .A1(clknet_1_1__leaf_net646),
    .A2(clknet_1_0__leaf_net645),
    .A3(net649),
    .S0(clknet_1_0__leaf_net655),
    .S1(net751),
    .X(net660));
 sky130_fd_sc_hd__mux4_1 c764 (.A0(clknet_1_1__leaf_net646),
    .A1(clknet_1_0__leaf_net651),
    .A2(net657),
    .A3(net647),
    .S0(clknet_1_0__leaf_net645),
    .S1(net751),
    .X(net661));
 sky130_fd_sc_hd__a2111o_1 c77 (.A1(net11),
    .A2(net12),
    .B1(net10),
    .C1(net13),
    .D1(net14),
    .X(net15));
 sky130_fd_sc_hd__and3_1 c78 (.A(net5),
    .B(net13),
    .C(net14),
    .X(net16));
 sky130_fd_sc_hd__or4bb_2 c79 (.A(net16),
    .B(net929),
    .C_N(net14),
    .D_N(net13),
    .X(net17));
 sky130_fd_sc_hd__a2111o_1 c80 (.A1(net13),
    .A2(net17),
    .B1(net10),
    .C1(net14),
    .D1(net929),
    .X(net18));
 sky130_fd_sc_hd__a2111o_1 c81 (.A1(net18),
    .A2(net929),
    .B1(net17),
    .C1(net13),
    .D1(net14),
    .X(net19));
 sky130_fd_sc_hd__mux4_1 c82 (.A0(net14),
    .A1(net17),
    .A2(net7),
    .A3(net19),
    .S0(net18),
    .S1(net13),
    .X(net20));
 sky130_fd_sc_hd__mux4_1 c83 (.A0(net15),
    .A1(net20),
    .A2(net18),
    .A3(net19),
    .S0(net929),
    .S1(net17),
    .X(net21));
 sky130_fd_sc_hd__mux4_1 c84 (.A0(net20),
    .A1(net17),
    .A2(net18),
    .A3(net12),
    .S0(net14),
    .S1(net21),
    .X(net22));
 sky130_fd_sc_hd__mux4_1 c85 (.A0(net21),
    .A1(net15),
    .A2(net18),
    .A3(net8),
    .S0(net11),
    .X(net23));
 sky130_fd_sc_hd__a2111o_1 c86 (.A1(net19),
    .A2(net13),
    .B1(net14),
    .C1(net17),
    .D1(net702),
    .X(net24));
 sky130_fd_sc_hd__mux4_1 c87 (.A0(net24),
    .A1(net19),
    .A2(net16),
    .A3(net20),
    .S0(net13),
    .S1(net702),
    .X(net25));
 sky130_fd_sc_hd__and2_1 c88 (.A(net10),
    .B(net929),
    .X(net26));
 sky130_fd_sc_hd__and2_2 c89 (.A(net26),
    .B(net10),
    .X(net27));
 sky130_fd_sc_hd__and2_1 c90 (.A(net27),
    .B(net26),
    .X(net28));
 sky130_fd_sc_hd__and2_1 c91 (.A(net26),
    .B(net27),
    .X(net29));
 sky130_fd_sc_hd__and3_1 c92 (.A(net28),
    .B(net26),
    .C(net919),
    .X(net30));
 sky130_fd_sc_hd__and3_1 c93 (.A(net919),
    .B(net27),
    .C(net28),
    .X(net31));
 sky130_fd_sc_hd__and3_1 c94 (.A(net26),
    .B(net919),
    .C(net10),
    .X(net32));
 sky130_fd_sc_hd__and3_1 c95 (.A(net31),
    .B(net919),
    .C(net28),
    .X(net33));
 sky130_fd_sc_hd__and2_0 c96 (.A(net27),
    .B(net919),
    .X(net34));
 sky130_fd_sc_hd__and2_1 c97 (.A(net919),
    .B(net30),
    .X(net35));
 sky130_fd_sc_hd__and3_1 c98 (.A(net33),
    .B(net35),
    .C(net919),
    .X(net36));
 sky130_fd_sc_hd__mux4_2 c99 (.A0(net30),
    .A1(net35),
    .A2(net31),
    .A3(net33),
    .S0(net919),
    .S1(net27),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_1 merge765 (.A(net752),
    .X(net662));
 sky130_fd_sc_hd__mux4_1 merge766 (.A0(clknet_1_0__leaf_net368),
    .A1(clknet_1_0__leaf_net270),
    .A2(clknet_1_0__leaf_net373),
    .A3(net369),
    .S0(clknet_1_0__leaf_net367),
    .S1(net749),
    .X(net663));
 sky130_fd_sc_hd__or4bb_1 merge767 (.A(net10),
    .B(net25),
    .C_N(net139),
    .D_N(net116),
    .X(net664));
 sky130_fd_sc_hd__or4bb_1 merge768 (.A(net474),
    .B(clknet_1_1__leaf_net373),
    .C_N(net933),
    .D_N(net801),
    .X(net665));
 sky130_fd_sc_hd__or4bb_1 merge769 (.A(net231),
    .B(net916),
    .C_N(net106),
    .D_N(net232),
    .X(net666));
 sky130_fd_sc_hd__or4bb_1 merge770 (.A(net116),
    .B(net869),
    .C_N(net114),
    .D_N(net870),
    .X(net667));
 sky130_fd_sc_hd__buf_1 merge771 (.A(clknet_1_0__leaf_net736),
    .X(net668));
 sky130_fd_sc_hd__sedfxtp_1 merge772 (.CLK(clknet_4_9_0_clk),
    .D(net167),
    .DE(clknet_1_1__leaf_net299),
    .SCD(clknet_1_1__leaf_net302),
    .SCE(net733),
    .Q(net669));
 sky130_fd_sc_hd__clkbuf_1 merge773 (.A(net832),
    .X(net670));
 sky130_fd_sc_hd__sdfrbp_1 merge774 (.CLK(clknet_4_7_0_clk),
    .D(clknet_1_0__leaf_net574),
    .RESET_B(clknet_1_0__leaf_net576),
    .SCD(clknet_1_0__leaf_net575),
    .SCE(net815),
    .Q(net672),
    .Q_N(net671));
 sky130_fd_sc_hd__clkbuf_1 merge775 (.A(net745),
    .X(net673));
 sky130_fd_sc_hd__sdfbbn_1 merge776 (.CLK_N(clknet_4_0_0_clk),
    .D(net213),
    .RESET_B(net210),
    .SCD(net922),
    .SET_B(net215),
    .Q(net214),
    .Q_N(net674));
 sky130_fd_sc_hd__or4bb_1 merge777 (.A(clknet_1_1__leaf_net645),
    .B(clknet_1_0__leaf_net644),
    .C_N(clknet_1_0__leaf_net646),
    .D_N(net823),
    .X(net676));
 sky130_fd_sc_hd__or4bb_1 merge778 (.A(net164),
    .B(net163),
    .C_N(clknet_1_0__leaf_net168),
    .D_N(net167),
    .X(net677));
 sky130_fd_sc_hd__dlymetal6s2s_1 merge779 (.A(net726),
    .X(net678));
 sky130_fd_sc_hd__sdfrbp_1 merge780 (.CLK(clknet_4_12_0_clk),
    .D(clknet_1_0__leaf_net415),
    .RESET_B(net946),
    .SCD(net508),
    .SCE(net917),
    .Q(net680),
    .Q_N(net679));
 sky130_fd_sc_hd__or4bb_1 merge781 (.A(net25),
    .B(clknet_1_0__leaf_net168),
    .C_N(net160),
    .D_N(net741),
    .X(net681));
 sky130_fd_sc_hd__mux4_1 merge782 (.A0(net209),
    .A1(net210),
    .A2(net213),
    .A3(net96),
    .S0(net915),
    .S1(net234),
    .X(net682));
 sky130_fd_sc_hd__sdfrtn_1 merge783 (.CLK_N(clknet_4_3_0_clk),
    .RESET_B(clknet_1_0__leaf_net257),
    .SCD(net116),
    .SCE(net260),
    .Q(net261));
 sky130_fd_sc_hd__a2111o_1 merge784 (.A1(clknet_1_0__leaf_net346),
    .A2(clknet_1_1__leaf_net251),
    .B1(net160),
    .C1(clknet_1_0__leaf_net270),
    .D1(net970),
    .X(net684));
 sky130_fd_sc_hd__mux4_1 merge785 (.A0(clknet_1_1__leaf_net635),
    .A1(clknet_1_1__leaf_net653),
    .A2(net649),
    .A3(net905),
    .S0(net652),
    .S1(clknet_1_1__leaf_net646),
    .X(net685));
 sky130_fd_sc_hd__a2111o_1 merge786 (.A1(net416),
    .A2(clknet_1_0__leaf_net373),
    .B1(clknet_1_1__leaf_net257),
    .C1(clknet_1_1__leaf_net256),
    .D1(net258),
    .X(net686));
 sky130_fd_sc_hd__mux4_1 merge787 (.A0(clknet_1_1__leaf_net467),
    .A1(clknet_1_1__leaf_net463),
    .A2(clknet_1_1__leaf_net460),
    .A3(net595),
    .S0(clknet_1_0__leaf_net575),
    .S1(net596),
    .X(net687));
 sky130_fd_sc_hd__mux4_1 merge788 (.A0(net65),
    .A1(net186),
    .A2(net164),
    .A3(net165),
    .S0(clknet_1_0__leaf_net168),
    .S1(net772),
    .X(net688));
 sky130_fd_sc_hd__mux4_1 merge789 (.A0(net255),
    .A1(clknet_1_0__leaf_net256),
    .A2(net96),
    .A3(clknet_1_1__leaf_net119),
    .S0(net116),
    .S1(clknet_1_0__leaf_net118),
    .X(net689));
 sky130_fd_sc_hd__mux4_1 merge790 (.A0(clknet_1_1__leaf_net561),
    .A1(clknet_1_1__leaf_net563),
    .A2(clknet_1_1__leaf_net560),
    .A3(clknet_1_1__leaf_net373),
    .S0(net485),
    .S1(net487),
    .X(net690));
 sky130_fd_sc_hd__sdfrtp_1 merge791 (.CLK(clknet_4_7_0_clk),
    .D(clknet_1_1__leaf_net573),
    .RESET_B(clknet_1_0__leaf_net575),
    .SCD(net579),
    .Q(net580));
 sky130_fd_sc_hd__mux4_1 merge792 (.A0(net286),
    .A1(net284),
    .A2(clknet_1_1__leaf_net270),
    .A3(clknet_1_0__leaf_net373),
    .S0(clknet_1_0__leaf_net395),
    .S1(net795),
    .X(net692));
 sky130_fd_sc_hd__or4bb_1 merge793 (.A(net120),
    .B(clknet_1_0__leaf_net118),
    .C_N(net116),
    .D_N(net115),
    .X(net693));
 sky130_fd_sc_hd__mux4_1 merge794 (.A0(net599),
    .A1(clknet_1_0__leaf_net634),
    .A2(clknet_1_0__leaf_net635),
    .A3(net595),
    .S0(clknet_1_1__leaf_net575),
    .S1(net596),
    .X(net694));
 sky130_fd_sc_hd__sdfbbn_1 merge795 (.CLK_N(clknet_4_11_0_clk),
    .D(net648),
    .RESET_B(net649),
    .SCD(clknet_1_1__leaf_net651),
    .SCE(clknet_1_1__leaf_net645),
    .SET_B(clknet_1_0__leaf_net646),
    .Q(net696),
    .Q_N(net695));
 sky130_fd_sc_hd__mux4_1 merge796 (.A0(clknet_1_1__leaf_net626),
    .A1(clknet_1_0__leaf_net646),
    .A2(net170),
    .A3(clknet_1_1__leaf_net168),
    .S0(net171),
    .S1(net703),
    .X(net697));
 sky130_fd_sc_hd__dfrbp_1 merge797 (.CLK(clknet_4_7_0_clk),
    .D(net569),
    .Q(net570),
    .Q_N(net698));
 sky130_fd_sc_hd__dfrbp_1 merge798 (.CLK(clknet_4_2_0_clk),
    .D(net135),
    .Q(net136),
    .Q_N(net700));
 sky130_fd_sc_hd__dfrtn_1 merge799 (.CLK_N(clknet_4_8_0_clk),
    .D(net22),
    .Q(net23));
 sky130_fd_sc_hd__dfrtp_1 merge800 (.CLK(clknet_4_11_0_clk),
    .D(net642),
    .Q(net703));
 sky130_fd_sc_hd__dfrtp_1 merge801 (.CLK(clknet_4_12_0_clk),
    .D(net499),
    .RESET_B(net665),
    .Q(net704));
 sky130_fd_sc_hd__dfrtp_1 merge802 (.CLK(clknet_4_10_0_clk),
    .D(net319),
    .RESET_B(net320),
    .Q(net705));
 sky130_fd_sc_hd__dfsbp_1 merge803 (.CLK(clknet_4_10_0_clk),
    .D(net202),
    .SET_B(net199),
    .Q(net707),
    .Q_N(net706));
 sky130_fd_sc_hd__and2_0 merge804 (.A(net253),
    .B(net254),
    .X(net708));
 sky130_fd_sc_hd__dfsbp_1 merge805 (.CLK(clknet_4_3_0_clk),
    .D(net271),
    .SET_B(net273),
    .Q(net710),
    .Q_N(net709));
 sky130_fd_sc_hd__dfstp_1 merge806 (.CLK(clknet_4_15_0_clk),
    .D(net548),
    .SET_B(net536),
    .Q(net711));
 sky130_fd_sc_hd__dfstp_1 merge807 (.CLK(clknet_4_13_0_clk),
    .D(net531),
    .SET_B(net520),
    .Q(net712));
 sky130_fd_sc_hd__dfstp_1 merge808 (.CLK(clknet_4_0_0_clk),
    .D(net107),
    .Q(net110));
 sky130_fd_sc_hd__dlrbn_1 merge809 (.D(net455),
    .GATE_N(clknet_4_4_0_clk),
    .RESET_B(net448),
    .Q(net715),
    .Q_N(net714));
 sky130_fd_sc_hd__dlrbn_1 merge810 (.D(net364),
    .GATE_N(clknet_4_4_0_clk),
    .Q(net365),
    .Q_N(net716));
 sky130_fd_sc_hd__dlrbp_1 merge811 (.D(net67),
    .GATE(clknet_4_10_0_clk),
    .RESET_B(net69),
    .Q(net718),
    .Q_N(net909));
 sky130_fd_sc_hd__dlrbp_1 merge812 (.D(net379),
    .GATE(clknet_4_6_0_clk),
    .RESET_B(net389),
    .Q(net720),
    .Q_N(net719));
 sky130_fd_sc_hd__and2_0 merge813 (.A(net618),
    .B(net616),
    .X(net721));
 sky130_fd_sc_hd__dlrtn_1 merge814 (.D(net466),
    .GATE_N(clknet_4_4_0_clk),
    .RESET_B(net478),
    .Q(net722));
 sky130_fd_sc_hd__and2_0 merge815 (.A(net179),
    .B(net183),
    .X(net723));
 sky130_fd_sc_hd__dlrtn_2 merge816 (.D(net159),
    .GATE_N(clknet_4_8_0_clk),
    .RESET_B(net664),
    .Q(net724));
 sky130_fd_sc_hd__and2_0 merge817 (.A(net90),
    .B(net91),
    .X(net725));
 sky130_fd_sc_hd__dlrtn_1 merge818 (.D(net431),
    .GATE_N(clknet_4_11_0_clk),
    .RESET_B(net686),
    .Q(net726));
 sky130_fd_sc_hd__and2_0 merge819 (.A(net661),
    .B(net656),
    .X(net727));
 sky130_fd_sc_hd__dlrtp_1 merge820 (.D(net337),
    .GATE(clknet_4_1_0_clk),
    .RESET_B(net343),
    .Q(net728));
 sky130_fd_sc_hd__dlrtp_1 merge821 (.GATE(clknet_4_9_0_clk),
    .RESET_B(net413),
    .Q(net414));
 sky130_fd_sc_hd__dlrtp_1 merge822 (.D(net220),
    .GATE(clknet_4_0_0_clk),
    .RESET_B(net221),
    .Q(net730));
 sky130_fd_sc_hd__and2_0 merge823 (.A(net44),
    .B(net45),
    .X(net731));
 sky130_fd_sc_hd__edfxbp_1 merge824 (.CLK(clknet_4_9_0_clk),
    .D(net300),
    .DE(net293),
    .Q(net733),
    .Q_N(net732));
 sky130_fd_sc_hd__edfxtp_1 merge825 (.CLK(clknet_4_13_0_clk),
    .D(net593),
    .DE(net578),
    .Q(net734));
 sky130_fd_sc_hd__sdlclkp_1 merge826 (.CLK(clknet_4_2_0_clk),
    .GATE(net731),
    .SCE(net667),
    .GCLK(net735));
 sky130_fd_sc_hd__sdlclkp_2 merge827 (.CLK(clknet_4_9_0_clk),
    .GATE(net298),
    .SCE(net692),
    .GCLK(net736));
 sky130_fd_sc_hd__sdlclkp_4 merge828 (.CLK(clknet_4_8_0_clk),
    .GATE(net181),
    .SCE(net677),
    .GCLK(net737));
 sky130_fd_sc_hd__dfrbp_1 merge829 (.CLK(clknet_4_0_0_clk),
    .D(net225),
    .RESET_B(net708),
    .Q(net739),
    .Q_N(net738));
 sky130_fd_sc_hd__dfrbp_1 merge830 (.CLK(clknet_4_8_0_clk),
    .D(net47),
    .RESET_B(net723),
    .Q(net741),
    .Q_N(net740));
 sky130_fd_sc_hd__dfrtn_1 merge831 (.CLK_N(clknet_4_8_0_clk),
    .D(net68),
    .RESET_B(net681),
    .Q(net742));
 sky130_fd_sc_hd__dfrtp_1 merge832 (.CLK(clknet_4_3_0_clk),
    .D(net274),
    .RESET_B(net392),
    .Q(net743));
 sky130_fd_sc_hd__dfrtp_1 merge833 (.CLK(clknet_4_1_0_clk),
    .D(net344),
    .RESET_B(net666),
    .Q(net744));
 sky130_fd_sc_hd__dfrtp_2 merge834 (.CLK(clknet_4_3_0_clk),
    .D(net366),
    .RESET_B(net684),
    .Q(net745));
 sky130_fd_sc_hd__and2_0 merge835 (.A(net727),
    .B(net660),
    .X(net746));
 sky130_fd_sc_hd__dfsbp_1 merge836 (.CLK(clknet_4_3_0_clk),
    .D(net275),
    .SET_B(net277),
    .Q(net748),
    .Q_N(net747));
 sky130_fd_sc_hd__dfsbp_1 merge837 (.CLK(clknet_4_1_0_clk),
    .D(net112),
    .SET_B(net278),
    .Q(net750),
    .Q_N(net749));
 sky130_fd_sc_hd__dfstp_1 merge838 (.CLK(clknet_4_11_0_clk),
    .SET_B(net746),
    .Q(net659));
 sky130_fd_sc_hd__dfstp_1 merge839 (.CLK(clknet_4_10_0_clk),
    .D(net321),
    .SET_B(net688),
    .Q(net752));
 sky130_fd_sc_hd__dfstp_1 merge840 (.CLK(clknet_4_7_0_clk),
    .D(net721),
    .SET_B(net568),
    .Q(net753));
 sky130_fd_sc_hd__dlrbn_1 merge841 (.D(net693),
    .GATE_N(clknet_4_2_0_clk),
    .RESET_B(net725),
    .Q(net755),
    .Q_N(net754));
 sky130_fd_sc_hd__dlrbn_1 merge842 (.D(net676),
    .GATE_N(clknet_4_11_0_clk),
    .RESET_B(net697),
    .Q(net757),
    .Q_N(net756));
 sky130_fd_sc_hd__dlrbp_1 merge843 (.D(net226),
    .GATE(clknet_4_0_0_clk),
    .Q(net227),
    .Q_N(net758));
 sky130_fd_sc_hd__dfxbp_1 s844 (.CLK(clknet_4_8_0_clk),
    .D(net43),
    .Q(net761),
    .Q_N(net760));
 sky130_fd_sc_hd__dfxbp_1 s845 (.CLK(clknet_4_0_0_clk),
    .D(net88),
    .Q(net763),
    .Q_N(net762));
 sky130_fd_sc_hd__dfxtp_1 s846 (.CLK(clknet_4_1_0_clk),
    .D(net109),
    .Q(net764));
 sky130_fd_sc_hd__dfxtp_1 s847 (.CLK(clknet_4_1_0_clk),
    .D(net111),
    .Q(net765));
 sky130_fd_sc_hd__dfxtp_1 s848 (.CLK(clknet_4_1_0_clk),
    .D(net113),
    .Q(net766));
 sky130_fd_sc_hd__dlclkp_1 s849 (.CLK(clknet_4_2_0_clk),
    .GATE(net132),
    .GCLK(net767));
 sky130_fd_sc_hd__dlclkp_2 s850 (.CLK(clknet_4_2_0_clk),
    .GATE(net154),
    .GCLK(net768));
 sky130_fd_sc_hd__dlclkp_4 s851 (.CLK(clknet_4_10_0_clk),
    .GATE(net173),
    .GCLK(net769));
 sky130_fd_sc_hd__dlxbn_1 s852 (.D(net177),
    .GATE_N(clknet_4_8_0_clk),
    .Q(net771),
    .Q_N(net770));
 sky130_fd_sc_hd__dlxbn_1 s853 (.D(net178),
    .GATE_N(clknet_4_8_0_clk),
    .Q(net773),
    .Q_N(net772));
 sky130_fd_sc_hd__dlxbp_1 s854 (.D(net201),
    .GATE(clknet_4_10_0_clk),
    .Q(net775),
    .Q_N(net774));
 sky130_fd_sc_hd__dlxtn_1 s855 (.D(net204),
    .GATE_N(clknet_4_10_0_clk),
    .Q(net776));
 sky130_fd_sc_hd__dlxtn_1 s856 (.D(net205),
    .GATE_N(clknet_4_10_0_clk),
    .Q(net777));
 sky130_fd_sc_hd__dlxtn_1 s857 (.D(net247),
    .GATE_N(clknet_4_1_0_clk),
    .Q(net778));
 sky130_fd_sc_hd__dlxtp_1 s858 (.D(net248),
    .GATE(clknet_4_1_0_clk),
    .Q(net779));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s859 (.D(net250),
    .SLEEP_B(clknet_4_1_0_clk),
    .Q(net780));
 sky130_fd_sc_hd__dfxbp_1 s860 (.CLK(clknet_4_3_0_clk),
    .D(net272),
    .Q(net782),
    .Q_N(net781));
 sky130_fd_sc_hd__dfxbp_1 s861 (.CLK(clknet_4_3_0_clk),
    .D(net276),
    .Q(net784),
    .Q_N(net783));
 sky130_fd_sc_hd__dfxtp_2 s862 (.CLK(clknet_4_9_0_clk),
    .D(net313),
    .Q(net908));
 sky130_fd_sc_hd__dfxtp_1 s863 (.CLK(clknet_4_11_0_clk),
    .D(net318),
    .Q(net785));
 sky130_fd_sc_hd__dfxtp_1 s864 (.CLK(clknet_4_10_0_clk),
    .D(net323),
    .Q(net899));
 sky130_fd_sc_hd__dlclkp_1 s865 (.CLK(clknet_4_4_0_clk),
    .GATE(net338),
    .GCLK(net786));
 sky130_fd_sc_hd__dlclkp_2 s866 (.CLK(clknet_4_4_0_clk),
    .GATE(net339),
    .GCLK(net787));
 sky130_fd_sc_hd__dlclkp_4 s867 (.CLK(clknet_4_4_0_clk),
    .GATE(net340),
    .GCLK(net788));
 sky130_fd_sc_hd__dlxbn_1 s868 (.D(net345),
    .GATE_N(clknet_4_4_0_clk),
    .Q(net790),
    .Q_N(net789));
 sky130_fd_sc_hd__dlxbn_1 s869 (.D(net390),
    .GATE_N(clknet_4_12_0_clk),
    .Q(net792),
    .Q_N(net791));
 sky130_fd_sc_hd__dlxbp_1 s870 (.D(net391),
    .GATE(clknet_4_9_0_clk),
    .Q(net794),
    .Q_N(net793));
 sky130_fd_sc_hd__dlxtn_1 s871 (.D(net393),
    .GATE_N(clknet_4_9_0_clk),
    .Q(net795));
 sky130_fd_sc_hd__dlxtn_1 s872 (.D(net433),
    .GATE_N(clknet_4_14_0_clk),
    .Q(net902));
 sky130_fd_sc_hd__dlxtn_1 s873 (.D(net451),
    .GATE_N(clknet_4_5_0_clk),
    .Q(net796));
 sky130_fd_sc_hd__dlxtp_1 s874 (.D(net452),
    .GATE(clknet_4_5_0_clk),
    .Q(net797));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s875 (.D(net453),
    .SLEEP_B(clknet_4_4_0_clk),
    .Q(net798));
 sky130_fd_sc_hd__dfxbp_1 s876 (.CLK(clknet_4_6_0_clk),
    .D(net469),
    .Q(net800),
    .Q_N(net799));
 sky130_fd_sc_hd__dfxbp_1 s877 (.CLK(clknet_4_6_0_clk),
    .D(net479),
    .Q(net802),
    .Q_N(net801));
 sky130_fd_sc_hd__dfxtp_1 s878 (.CLK(clknet_4_6_0_clk),
    .D(net481),
    .Q(net803));
 sky130_fd_sc_hd__dfxtp_1 s879 (.CLK(clknet_4_6_0_clk),
    .D(net482),
    .Q(net804));
 sky130_fd_sc_hd__dfxtp_1 s880 (.CLK(clknet_4_13_0_clk),
    .D(net518),
    .Q(net805));
 sky130_fd_sc_hd__dlclkp_1 s881 (.CLK(clknet_4_15_0_clk),
    .GATE(net525),
    .GCLK(net806));
 sky130_fd_sc_hd__dlclkp_2 s882 (.CLK(clknet_4_15_0_clk),
    .GATE(net529),
    .GCLK(net807));
 sky130_fd_sc_hd__dlclkp_4 s883 (.CLK(clknet_4_14_0_clk),
    .GATE(net540),
    .GCLK(net808));
 sky130_fd_sc_hd__dlxbn_1 s884 (.D(net542),
    .GATE_N(clknet_4_14_0_clk),
    .Q(net901),
    .Q_N(net895));
 sky130_fd_sc_hd__dlxbn_1 s885 (.D(net543),
    .GATE_N(clknet_4_14_0_clk),
    .Q(net810),
    .Q_N(net809));
 sky130_fd_sc_hd__dlxbp_1 s886 (.D(net544),
    .GATE(clknet_4_15_0_clk),
    .Q(net812),
    .Q_N(net811));
 sky130_fd_sc_hd__dlxtn_1 s887 (.D(net545),
    .GATE_N(clknet_4_15_0_clk),
    .Q(net813));
 sky130_fd_sc_hd__dlxtn_1 s888 (.D(net546),
    .GATE_N(clknet_4_14_0_clk),
    .Q(net814));
 sky130_fd_sc_hd__dlxtn_2 s889 (.D(net565),
    .GATE_N(clknet_4_7_0_clk),
    .Q(net815));
 sky130_fd_sc_hd__dlxtp_1 s890 (.D(net592),
    .GATE(clknet_4_13_0_clk),
    .Q(net816));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s891 (.D(net594),
    .SLEEP_B(clknet_4_13_0_clk),
    .Q(net817));
 sky130_fd_sc_hd__dfxbp_1 s892 (.CLK(clknet_4_13_0_clk),
    .D(net617),
    .Q(net819),
    .Q_N(net818));
 sky130_fd_sc_hd__dfxbp_1 s893 (.CLK(clknet_4_12_0_clk),
    .D(net638),
    .Q(net821),
    .Q_N(net820));
 sky130_fd_sc_hd__dfxtp_1 s894 (.CLK(clknet_4_11_0_clk),
    .D(net640),
    .Q(net822));
 sky130_fd_sc_hd__dfxtp_1 s895 (.CLK(clknet_4_11_0_clk),
    .D(net641),
    .Q(net823));
 sky130_fd_sc_hd__dfxtp_1 s896 (.CLK(clknet_4_3_0_clk),
    .D(net663),
    .Q(net824));
 sky130_fd_sc_hd__dlclkp_1 s897 (.CLK(clknet_4_0_0_clk),
    .GATE(net682),
    .GCLK(net825));
 sky130_fd_sc_hd__dlclkp_2 s898 (.CLK(clknet_4_11_0_clk),
    .GATE(net685),
    .GCLK(net826));
 sky130_fd_sc_hd__dlclkp_4 s899 (.CLK(clknet_4_6_0_clk),
    .GATE(net687),
    .GCLK(net827));
 sky130_fd_sc_hd__dlxbn_1 s900 (.D(net689),
    .GATE_N(clknet_4_3_0_clk),
    .Q(net829),
    .Q_N(net828));
 sky130_fd_sc_hd__dlxbn_1 s901 (.D(net690),
    .GATE_N(clknet_4_7_0_clk),
    .Q(net831),
    .Q_N(net830));
 sky130_fd_sc_hd__dlxbp_1 s902 (.D(net694),
    .GATE(clknet_4_12_0_clk),
    .Q(net833),
    .Q_N(net832));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Right_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Right_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Right_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Right_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Right_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Right_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Right_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Right_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Right_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Right_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Right_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Right_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Right_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Right_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Right_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Right_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Right_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Right_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Right_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Right_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Right_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_161 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_162 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_163 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_164 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_165 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_166 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_167 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_168 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_169 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_170 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_171 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_172 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_173 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_174 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_175 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_176 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_177 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_178 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_179 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_180 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_181 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_182 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Left_183 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Left_184 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Left_185 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Left_186 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Left_187 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Left_188 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Left_189 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Left_190 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Left_191 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Left_192 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Left_193 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Left_194 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Left_195 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Left_196 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Left_197 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Left_198 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Left_199 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Left_200 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Left_201 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Left_202 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Left_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1347 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(in0),
    .X(net643));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(in1),
    .X(net675));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(in10),
    .X(net699));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(in11),
    .X(net834));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(in12),
    .X(net835));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(in13),
    .X(net836));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(in14),
    .X(net837));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(in15),
    .X(net838));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(in16),
    .X(net839));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(in17),
    .X(net840));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(in18),
    .X(net841));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(in19),
    .X(net842));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(in2),
    .X(net843));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(in20),
    .X(net844));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(in21),
    .X(net845));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(in22),
    .X(net846));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(in23),
    .X(net847));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(in24),
    .X(net848));
 sky130_fd_sc_hd__buf_1 input19 (.A(in25),
    .X(net849));
 sky130_fd_sc_hd__clkbuf_1 input20 (.A(in26),
    .X(net850));
 sky130_fd_sc_hd__clkbuf_1 input21 (.A(in27),
    .X(net851));
 sky130_fd_sc_hd__clkbuf_1 input22 (.A(in28),
    .X(net852));
 sky130_fd_sc_hd__clkbuf_1 input23 (.A(in29),
    .X(net853));
 sky130_fd_sc_hd__clkbuf_1 input24 (.A(in3),
    .X(net854));
 sky130_fd_sc_hd__clkbuf_1 input25 (.A(in30),
    .X(net855));
 sky130_fd_sc_hd__clkbuf_1 input26 (.A(in31),
    .X(net856));
 sky130_fd_sc_hd__clkbuf_1 input27 (.A(in32),
    .X(net857));
 sky130_fd_sc_hd__clkbuf_1 input28 (.A(in33),
    .X(net858));
 sky130_fd_sc_hd__clkbuf_1 input29 (.A(in34),
    .X(net859));
 sky130_fd_sc_hd__clkbuf_1 input30 (.A(in35),
    .X(net860));
 sky130_fd_sc_hd__clkbuf_1 input31 (.A(in36),
    .X(net861));
 sky130_fd_sc_hd__clkbuf_1 input32 (.A(in37),
    .X(net862));
 sky130_fd_sc_hd__clkbuf_1 input33 (.A(in38),
    .X(net863));
 sky130_fd_sc_hd__clkbuf_1 input34 (.A(in39),
    .X(net864));
 sky130_fd_sc_hd__clkbuf_1 input35 (.A(in4),
    .X(net865));
 sky130_fd_sc_hd__buf_1 input36 (.A(net953),
    .X(net866));
 sky130_fd_sc_hd__clkbuf_1 input37 (.A(in41),
    .X(net867));
 sky130_fd_sc_hd__clkbuf_1 input38 (.A(in42),
    .X(net868));
 sky130_fd_sc_hd__clkbuf_1 input39 (.A(in43),
    .X(net869));
 sky130_fd_sc_hd__clkbuf_1 input40 (.A(in44),
    .X(net870));
 sky130_fd_sc_hd__buf_1 input41 (.A(in45),
    .X(net871));
 sky130_fd_sc_hd__clkbuf_1 input42 (.A(in46),
    .X(net872));
 sky130_fd_sc_hd__clkbuf_1 input43 (.A(in47),
    .X(net873));
 sky130_fd_sc_hd__clkbuf_1 input44 (.A(in48),
    .X(net874));
 sky130_fd_sc_hd__buf_1 input45 (.A(in49),
    .X(net875));
 sky130_fd_sc_hd__clkbuf_1 input46 (.A(in5),
    .X(net876));
 sky130_fd_sc_hd__clkbuf_1 input47 (.A(in50),
    .X(net877));
 sky130_fd_sc_hd__clkbuf_1 input48 (.A(in51),
    .X(net878));
 sky130_fd_sc_hd__clkbuf_1 input49 (.A(in52),
    .X(net879));
 sky130_fd_sc_hd__clkbuf_1 input50 (.A(in53),
    .X(net880));
 sky130_fd_sc_hd__clkbuf_1 input51 (.A(in54),
    .X(net881));
 sky130_fd_sc_hd__clkbuf_1 input52 (.A(in55),
    .X(net882));
 sky130_fd_sc_hd__clkbuf_1 input53 (.A(in56),
    .X(net883));
 sky130_fd_sc_hd__clkbuf_1 input54 (.A(in57),
    .X(net884));
 sky130_fd_sc_hd__clkbuf_1 input55 (.A(in58),
    .X(net885));
 sky130_fd_sc_hd__clkbuf_1 input56 (.A(in59),
    .X(net886));
 sky130_fd_sc_hd__clkbuf_1 input57 (.A(in6),
    .X(net887));
 sky130_fd_sc_hd__clkbuf_1 input58 (.A(in60),
    .X(net888));
 sky130_fd_sc_hd__clkbuf_1 input59 (.A(in61),
    .X(net889));
 sky130_fd_sc_hd__clkbuf_1 input60 (.A(in7),
    .X(net890));
 sky130_fd_sc_hd__clkbuf_1 input61 (.A(in8),
    .X(net891));
 sky130_fd_sc_hd__clkbuf_1 input62 (.A(in9),
    .X(net892));
 sky130_fd_sc_hd__buf_2 output63 (.A(net893),
    .X(out0));
 sky130_fd_sc_hd__buf_2 output64 (.A(net894),
    .X(out10));
 sky130_fd_sc_hd__buf_2 output65 (.A(net895),
    .X(out14));
 sky130_fd_sc_hd__buf_2 output66 (.A(net896),
    .X(out16));
 sky130_fd_sc_hd__buf_2 output67 (.A(net897),
    .X(out17));
 sky130_fd_sc_hd__buf_2 output68 (.A(net898),
    .X(out19));
 sky130_fd_sc_hd__buf_2 output69 (.A(net899),
    .X(out22));
 sky130_fd_sc_hd__buf_2 output70 (.A(net900),
    .X(out28));
 sky130_fd_sc_hd__buf_2 output71 (.A(net901),
    .X(out3));
 sky130_fd_sc_hd__buf_2 output72 (.A(net902),
    .X(out31));
 sky130_fd_sc_hd__buf_2 output73 (.A(net903),
    .X(out32));
 sky130_fd_sc_hd__buf_2 output74 (.A(net904),
    .X(out39));
 sky130_fd_sc_hd__buf_2 output75 (.A(net905),
    .X(out4));
 sky130_fd_sc_hd__buf_2 output76 (.A(net906),
    .X(out40));
 sky130_fd_sc_hd__buf_2 output77 (.A(net907),
    .X(out41));
 sky130_fd_sc_hd__buf_2 output78 (.A(net908),
    .X(out42));
 sky130_fd_sc_hd__buf_2 output79 (.A(net909),
    .X(out43));
 sky130_fd_sc_hd__clkbuf_1 output80 (.A(clknet_1_1__leaf_net910),
    .X(out47));
 sky130_fd_sc_hd__buf_2 output81 (.A(net911),
    .X(out49));
 sky130_fd_sc_hd__buf_2 output82 (.A(net912),
    .X(out50));
 sky130_fd_sc_hd__clkbuf_1 output83 (.A(net913),
    .X(out54));
 sky130_fd_sc_hd__buf_2 output84 (.A(net914),
    .X(out7));
 sky130_fd_sc_hd__buf_2 fanout85 (.A(net230),
    .X(net915));
 sky130_fd_sc_hd__buf_2 fanout86 (.A(net230),
    .X(net916));
 sky130_fd_sc_hd__buf_2 fanout87 (.A(net506),
    .X(net917));
 sky130_fd_sc_hd__clkbuf_2 fanout88 (.A(net506),
    .X(net918));
 sky130_fd_sc_hd__clkbuf_2 fanout89 (.A(net29),
    .X(net919));
 sky130_fd_sc_hd__buf_8 fanout90 (.A(net148),
    .X(net920));
 sky130_fd_sc_hd__clkbuf_2 fanout91 (.A(net324),
    .X(net921));
 sky130_fd_sc_hd__buf_2 fanout92 (.A(net206),
    .X(net922));
 sky130_fd_sc_hd__clkbuf_2 fanout93 (.A(net189),
    .X(net923));
 sky130_fd_sc_hd__buf_1 fanout94 (.A(net189),
    .X(net924));
 sky130_fd_sc_hd__buf_6 fanout95 (.A(net144),
    .X(net925));
 sky130_fd_sc_hd__clkbuf_4 fanout96 (.A(net927),
    .X(net926));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout97 (.A(net928),
    .X(net927));
 sky130_fd_sc_hd__clkbuf_2 fanout98 (.A(net76),
    .X(net928));
 sky130_fd_sc_hd__buf_2 fanout99 (.A(net8),
    .X(net929));
 sky130_fd_sc_hd__clkbuf_2 fanout100 (.A(net51),
    .X(net930));
 sky130_fd_sc_hd__buf_2 fanout101 (.A(net94),
    .X(net931));
 sky130_fd_sc_hd__clkbuf_2 fanout102 (.A(net48),
    .X(net932));
 sky130_fd_sc_hd__buf_2 fanout103 (.A(net798),
    .X(net933));
 sky130_fd_sc_hd__buf_2 fanout104 (.A(net533),
    .X(net934));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net827 (.A(net827),
    .X(clknet_0_net827));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net827 (.A(clknet_0_net827),
    .X(clknet_1_0__leaf_net827));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net827 (.A(clknet_0_net827),
    .X(clknet_1_1__leaf_net827));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net597 (.A(net597),
    .X(clknet_0_net597));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net597 (.A(clknet_0_net597),
    .X(clknet_1_0__leaf_net597));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net597 (.A(clknet_0_net597),
    .X(clknet_1_1__leaf_net597));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net621 (.A(net621),
    .X(clknet_0_net621));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net621 (.A(clknet_0_net621),
    .X(clknet_1_0__leaf_net621));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net621 (.A(clknet_0_net621),
    .X(clknet_1_1__leaf_net621));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net644 (.A(net644),
    .X(clknet_0_net644));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net644 (.A(clknet_0_net644),
    .X(clknet_1_0__leaf_net644));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net644 (.A(clknet_0_net644),
    .X(clknet_1_1__leaf_net644));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net646 (.A(net646),
    .X(clknet_0_net646));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net646 (.A(clknet_0_net646),
    .X(clknet_1_0__leaf_net646));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net646 (.A(clknet_0_net646),
    .X(clknet_1_1__leaf_net646));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net826 (.A(net826),
    .X(clknet_0_net826));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net826 (.A(clknet_0_net826),
    .X(clknet_1_0__leaf_net826));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net826 (.A(clknet_0_net826),
    .X(clknet_1_1__leaf_net826));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net654 (.A(net654),
    .X(clknet_0_net654));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net654 (.A(clknet_0_net654),
    .X(clknet_1_0__leaf_net654));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net654 (.A(clknet_0_net654),
    .X(clknet_1_1__leaf_net654));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net653 (.A(net653),
    .X(clknet_0_net653));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net653 (.A(clknet_0_net653),
    .X(clknet_1_0__leaf_net653));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net653 (.A(clknet_0_net653),
    .X(clknet_1_1__leaf_net653));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net645 (.A(net645),
    .X(clknet_0_net645));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net645 (.A(clknet_0_net645),
    .X(clknet_1_0__leaf_net645));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net645 (.A(clknet_0_net645),
    .X(clknet_1_1__leaf_net645));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net655 (.A(net655),
    .X(clknet_0_net655));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net655 (.A(clknet_0_net655),
    .X(clknet_1_0__leaf_net655));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net655 (.A(clknet_0_net655),
    .X(clknet_1_1__leaf_net655));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net651 (.A(net651),
    .X(clknet_0_net651));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net651 (.A(clknet_0_net651),
    .X(clknet_1_0__leaf_net651));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net651 (.A(clknet_0_net651),
    .X(clknet_1_1__leaf_net651));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net625 (.A(net625),
    .X(clknet_0_net625));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net625 (.A(clknet_0_net625),
    .X(clknet_1_0__leaf_net625));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net625 (.A(clknet_0_net625),
    .X(clknet_1_1__leaf_net625));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net636 (.A(net636),
    .X(clknet_0_net636));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net636 (.A(clknet_0_net636),
    .X(clknet_1_0__leaf_net636));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net636 (.A(clknet_0_net636),
    .X(clknet_1_1__leaf_net636));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net623 (.A(net623),
    .X(clknet_0_net623));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net623 (.A(clknet_0_net623),
    .X(clknet_1_0__leaf_net623));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net623 (.A(clknet_0_net623),
    .X(clknet_1_1__leaf_net623));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net633 (.A(net633),
    .X(clknet_0_net633));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net633 (.A(clknet_0_net633),
    .X(clknet_1_0__leaf_net633));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net633 (.A(clknet_0_net633),
    .X(clknet_1_1__leaf_net633));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net629 (.A(net629),
    .X(clknet_0_net629));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net629 (.A(clknet_0_net629),
    .X(clknet_1_0__leaf_net629));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net629 (.A(clknet_0_net629),
    .X(clknet_1_1__leaf_net629));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net635 (.A(net635),
    .X(clknet_0_net635));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net635 (.A(clknet_0_net635),
    .X(clknet_1_0__leaf_net635));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net635 (.A(clknet_0_net635),
    .X(clknet_1_1__leaf_net635));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net634 (.A(net634),
    .X(clknet_0_net634));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net634 (.A(clknet_0_net634),
    .X(clknet_1_0__leaf_net634));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net634 (.A(clknet_0_net634),
    .X(clknet_1_1__leaf_net634));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net632 (.A(net632),
    .X(clknet_0_net632));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net632 (.A(clknet_0_net632),
    .X(clknet_1_0__leaf_net632));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net632 (.A(clknet_0_net632),
    .X(clknet_1_1__leaf_net632));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net631 (.A(net631),
    .X(clknet_0_net631));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net631 (.A(clknet_0_net631),
    .X(clknet_1_0__leaf_net631));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net631 (.A(clknet_0_net631),
    .X(clknet_1_1__leaf_net631));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net630 (.A(net630),
    .X(clknet_0_net630));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net630 (.A(clknet_0_net630),
    .X(clknet_1_0__leaf_net630));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net630 (.A(clknet_0_net630),
    .X(clknet_1_1__leaf_net630));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net626 (.A(net626),
    .X(clknet_0_net626));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net626 (.A(clknet_0_net626),
    .X(clknet_1_0__leaf_net626));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net626 (.A(clknet_0_net626),
    .X(clknet_1_1__leaf_net626));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net624 (.A(net624),
    .X(clknet_0_net624));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net624 (.A(clknet_0_net624),
    .X(clknet_1_0__leaf_net624));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net624 (.A(clknet_0_net624),
    .X(clknet_1_1__leaf_net624));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net622 (.A(net622),
    .X(clknet_0_net622));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net622 (.A(clknet_0_net622),
    .X(clknet_1_0__leaf_net622));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net622 (.A(clknet_0_net622),
    .X(clknet_1_1__leaf_net622));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net607 (.A(net607),
    .X(clknet_0_net607));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net607 (.A(clknet_0_net607),
    .X(clknet_1_0__leaf_net607));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net607 (.A(clknet_0_net607),
    .X(clknet_1_1__leaf_net607));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net609 (.A(net609),
    .X(clknet_0_net609));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net609 (.A(clknet_0_net609),
    .X(clknet_1_0__leaf_net609));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net609 (.A(clknet_0_net609),
    .X(clknet_1_1__leaf_net609));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net608 (.A(net608),
    .X(clknet_0_net608));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net608 (.A(clknet_0_net608),
    .X(clknet_1_0__leaf_net608));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net608 (.A(clknet_0_net608),
    .X(clknet_1_1__leaf_net608));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net600 (.A(net600),
    .X(clknet_0_net600));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net600 (.A(clknet_0_net600),
    .X(clknet_1_0__leaf_net600));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net600 (.A(clknet_0_net600),
    .X(clknet_1_1__leaf_net600));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net603 (.A(net603),
    .X(clknet_0_net603));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net603 (.A(clknet_0_net603),
    .X(clknet_1_0__leaf_net603));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net603 (.A(clknet_0_net603),
    .X(clknet_1_1__leaf_net603));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net604 (.A(net604),
    .X(clknet_0_net604));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net604 (.A(clknet_0_net604),
    .X(clknet_1_0__leaf_net604));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net604 (.A(clknet_0_net604),
    .X(clknet_1_1__leaf_net604));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net606 (.A(net606),
    .X(clknet_0_net606));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net606 (.A(clknet_0_net606),
    .X(clknet_1_0__leaf_net606));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net606 (.A(clknet_0_net606),
    .X(clknet_1_1__leaf_net606));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net468 (.A(net468),
    .X(clknet_0_net468));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net468 (.A(clknet_0_net468),
    .X(clknet_1_0__leaf_net468));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net468 (.A(clknet_0_net468),
    .X(clknet_1_1__leaf_net468));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net825 (.A(net825),
    .X(clknet_0_net825));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net825 (.A(clknet_0_net825),
    .X(clknet_1_0__leaf_net825));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net825 (.A(clknet_0_net825),
    .X(clknet_1_1__leaf_net825));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net238 (.A(net238),
    .X(clknet_0_net238));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net238 (.A(clknet_0_net238),
    .X(clknet_1_0__leaf_net238));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net238 (.A(clknet_0_net238),
    .X(clknet_1_1__leaf_net238));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net251 (.A(net251),
    .X(clknet_0_net251));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net251 (.A(clknet_0_net251),
    .X(clknet_1_0__leaf_net251));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net251 (.A(clknet_0_net251),
    .X(clknet_1_1__leaf_net251));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net239 (.A(net239),
    .X(clknet_0_net239));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net239 (.A(clknet_0_net239),
    .X(clknet_1_0__leaf_net239));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net239 (.A(clknet_0_net239),
    .X(clknet_1_1__leaf_net239));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net808 (.A(net808),
    .X(clknet_0_net808));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net808 (.A(clknet_0_net808),
    .X(clknet_1_0__leaf_net808));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net808 (.A(clknet_0_net808),
    .X(clknet_1_1__leaf_net808));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net541 (.A(net541),
    .X(clknet_0_net541));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net541 (.A(clknet_0_net541),
    .X(clknet_1_0__leaf_net541));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net541 (.A(clknet_0_net541),
    .X(clknet_1_1__leaf_net541));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net807 (.A(net807),
    .X(clknet_0_net807));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net807 (.A(clknet_0_net807),
    .X(clknet_1_0__leaf_net807));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net807 (.A(clknet_0_net807),
    .X(clknet_1_1__leaf_net807));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net806 (.A(net806),
    .X(clknet_0_net806));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net806 (.A(clknet_0_net806),
    .X(clknet_1_0__leaf_net806));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net806 (.A(clknet_0_net806),
    .X(clknet_1_1__leaf_net806));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net528 (.A(net528),
    .X(clknet_0_net528));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net528 (.A(clknet_0_net528),
    .X(clknet_1_0__leaf_net528));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net528 (.A(clknet_0_net528),
    .X(clknet_1_1__leaf_net528));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net788 (.A(net788),
    .X(clknet_0_net788));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net788 (.A(clknet_0_net788),
    .X(clknet_1_0__leaf_net788));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net788 (.A(clknet_0_net788),
    .X(clknet_1_1__leaf_net788));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net549 (.A(net549),
    .X(clknet_0_net549));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net549 (.A(clknet_0_net549),
    .X(clknet_1_0__leaf_net549));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net549 (.A(clknet_0_net549),
    .X(clknet_1_1__leaf_net549));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net567 (.A(net567),
    .X(clknet_0_net567));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net567 (.A(clknet_0_net567),
    .X(clknet_1_0__leaf_net567));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net567 (.A(clknet_0_net567),
    .X(clknet_1_1__leaf_net567));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net555 (.A(net555),
    .X(clknet_0_net555));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net555 (.A(clknet_0_net555),
    .X(clknet_1_0__leaf_net555));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net555 (.A(clknet_0_net555),
    .X(clknet_1_1__leaf_net555));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net563 (.A(net563),
    .X(clknet_0_net563));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net563 (.A(clknet_0_net563),
    .X(clknet_1_0__leaf_net563));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net563 (.A(clknet_0_net563),
    .X(clknet_1_1__leaf_net563));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net562 (.A(net562),
    .X(clknet_0_net562));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net562 (.A(clknet_0_net562),
    .X(clknet_1_0__leaf_net562));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net562 (.A(clknet_0_net562),
    .X(clknet_1_1__leaf_net562));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net566 (.A(net566),
    .X(clknet_0_net566));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net566 (.A(clknet_0_net566),
    .X(clknet_1_0__leaf_net566));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net566 (.A(clknet_0_net566),
    .X(clknet_1_1__leaf_net566));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net556 (.A(net556),
    .X(clknet_0_net556));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net556 (.A(clknet_0_net556),
    .X(clknet_1_0__leaf_net556));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net556 (.A(clknet_0_net556),
    .X(clknet_1_1__leaf_net556));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net560 (.A(net560),
    .X(clknet_0_net560));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net560 (.A(clknet_0_net560),
    .X(clknet_1_0__leaf_net560));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net560 (.A(clknet_0_net560),
    .X(clknet_1_1__leaf_net560));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net559 (.A(net559),
    .X(clknet_0_net559));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net559 (.A(clknet_0_net559),
    .X(clknet_1_0__leaf_net559));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net559 (.A(clknet_0_net559),
    .X(clknet_1_1__leaf_net559));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net557 (.A(net557),
    .X(clknet_0_net557));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net557 (.A(clknet_0_net557),
    .X(clknet_1_0__leaf_net557));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net557 (.A(clknet_0_net557),
    .X(clknet_1_1__leaf_net557));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net558 (.A(net558),
    .X(clknet_0_net558));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net558 (.A(clknet_0_net558),
    .X(clknet_1_0__leaf_net558));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net558 (.A(clknet_0_net558),
    .X(clknet_1_1__leaf_net558));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net561 (.A(net561),
    .X(clknet_0_net561));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net561 (.A(clknet_0_net561),
    .X(clknet_1_0__leaf_net561));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net561 (.A(clknet_0_net561),
    .X(clknet_1_1__leaf_net561));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net552 (.A(net552),
    .X(clknet_0_net552));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net552 (.A(clknet_0_net552),
    .X(clknet_1_0__leaf_net552));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net552 (.A(clknet_0_net552),
    .X(clknet_1_1__leaf_net552));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net554 (.A(net554),
    .X(clknet_0_net554));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net554 (.A(clknet_0_net554),
    .X(clknet_1_0__leaf_net554));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net554 (.A(clknet_0_net554),
    .X(clknet_1_1__leaf_net554));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net551 (.A(net551),
    .X(clknet_0_net551));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net551 (.A(clknet_0_net551),
    .X(clknet_1_0__leaf_net551));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net551 (.A(clknet_0_net551),
    .X(clknet_1_1__leaf_net551));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net550 (.A(net550),
    .X(clknet_0_net550));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net550 (.A(clknet_0_net550),
    .X(clknet_1_0__leaf_net550));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net550 (.A(clknet_0_net550),
    .X(clknet_1_1__leaf_net550));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net553 (.A(net553),
    .X(clknet_0_net553));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net553 (.A(clknet_0_net553),
    .X(clknet_1_0__leaf_net553));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net553 (.A(clknet_0_net553),
    .X(clknet_1_1__leaf_net553));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net439 (.A(net439),
    .X(clknet_0_net439));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net439 (.A(clknet_0_net439),
    .X(clknet_1_0__leaf_net439));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net439 (.A(clknet_0_net439),
    .X(clknet_1_1__leaf_net439));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net449 (.A(net449),
    .X(clknet_0_net449));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net449 (.A(clknet_0_net449),
    .X(clknet_1_0__leaf_net449));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net449 (.A(clknet_0_net449),
    .X(clknet_1_1__leaf_net449));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net450 (.A(net450),
    .X(clknet_0_net450));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net450 (.A(clknet_0_net450),
    .X(clknet_1_0__leaf_net450));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net450 (.A(clknet_0_net450),
    .X(clknet_1_1__leaf_net450));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net446 (.A(net446),
    .X(clknet_0_net446));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net446 (.A(clknet_0_net446),
    .X(clknet_1_0__leaf_net446));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net446 (.A(clknet_0_net446),
    .X(clknet_1_1__leaf_net446));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net444 (.A(net444),
    .X(clknet_0_net444));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net444 (.A(clknet_0_net444),
    .X(clknet_1_0__leaf_net444));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net444 (.A(clknet_0_net444),
    .X(clknet_1_1__leaf_net444));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net445 (.A(net445),
    .X(clknet_0_net445));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net445 (.A(clknet_0_net445),
    .X(clknet_1_0__leaf_net445));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net445 (.A(clknet_0_net445),
    .X(clknet_1_1__leaf_net445));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net447 (.A(net447),
    .X(clknet_0_net447));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net447 (.A(clknet_0_net447),
    .X(clknet_1_0__leaf_net447));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net447 (.A(clknet_0_net447),
    .X(clknet_1_1__leaf_net447));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net442 (.A(net442),
    .X(clknet_0_net442));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net442 (.A(clknet_0_net442),
    .X(clknet_1_0__leaf_net442));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net442 (.A(clknet_0_net442),
    .X(clknet_1_1__leaf_net442));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net443 (.A(net443),
    .X(clknet_0_net443));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net443 (.A(clknet_0_net443),
    .X(clknet_1_0__leaf_net443));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net443 (.A(clknet_0_net443),
    .X(clknet_1_1__leaf_net443));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net441 (.A(net441),
    .X(clknet_0_net441));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net441 (.A(clknet_0_net441),
    .X(clknet_1_0__leaf_net441));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net441 (.A(clknet_0_net441),
    .X(clknet_1_1__leaf_net441));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net440 (.A(net440),
    .X(clknet_0_net440));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net440 (.A(clknet_0_net440),
    .X(clknet_1_0__leaf_net440));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net440 (.A(clknet_0_net440),
    .X(clknet_1_1__leaf_net440));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net434 (.A(net434),
    .X(clknet_0_net434));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net434 (.A(clknet_0_net434),
    .X(clknet_1_0__leaf_net434));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net434 (.A(clknet_0_net434),
    .X(clknet_1_1__leaf_net434));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net436 (.A(net436),
    .X(clknet_0_net436));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net436 (.A(clknet_0_net436),
    .X(clknet_1_0__leaf_net436));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net436 (.A(clknet_0_net436),
    .X(clknet_1_1__leaf_net436));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net437 (.A(net437),
    .X(clknet_0_net437));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net437 (.A(clknet_0_net437),
    .X(clknet_1_0__leaf_net437));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net437 (.A(clknet_0_net437),
    .X(clknet_1_1__leaf_net437));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net438 (.A(net438),
    .X(clknet_0_net438));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net438 (.A(clknet_0_net438),
    .X(clknet_1_0__leaf_net438));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net438 (.A(clknet_0_net438),
    .X(clknet_1_1__leaf_net438));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net435 (.A(net435),
    .X(clknet_0_net435));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net435 (.A(clknet_0_net435),
    .X(clknet_1_0__leaf_net435));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net435 (.A(clknet_0_net435),
    .X(clknet_1_1__leaf_net435));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net346 (.A(net346),
    .X(clknet_0_net346));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net346 (.A(clknet_0_net346),
    .X(clknet_1_0__leaf_net346));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net346 (.A(clknet_0_net346),
    .X(clknet_1_1__leaf_net346));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net360 (.A(net360),
    .X(clknet_0_net360));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net360 (.A(clknet_0_net360),
    .X(clknet_1_0__leaf_net360));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net360 (.A(clknet_0_net360),
    .X(clknet_1_1__leaf_net360));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net363 (.A(net363),
    .X(clknet_0_net363));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net363 (.A(clknet_0_net363),
    .X(clknet_1_0__leaf_net363));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net363 (.A(clknet_0_net363),
    .X(clknet_1_1__leaf_net363));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net362 (.A(net362),
    .X(clknet_0_net362));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net362 (.A(clknet_0_net362),
    .X(clknet_1_0__leaf_net362));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net362 (.A(clknet_0_net362),
    .X(clknet_1_1__leaf_net362));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net361 (.A(net361),
    .X(clknet_0_net361));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net361 (.A(clknet_0_net361),
    .X(clknet_1_0__leaf_net361));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net361 (.A(clknet_0_net361),
    .X(clknet_1_1__leaf_net361));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net359 (.A(net359),
    .X(clknet_0_net359));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net359 (.A(clknet_0_net359),
    .X(clknet_1_0__leaf_net359));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net359 (.A(clknet_0_net359),
    .X(clknet_1_1__leaf_net359));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net572 (.A(net572),
    .X(clknet_0_net572));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net572 (.A(clknet_0_net572),
    .X(clknet_1_0__leaf_net572));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net572 (.A(clknet_0_net572),
    .X(clknet_1_1__leaf_net572));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net589 (.A(net589),
    .X(clknet_0_net589));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net589 (.A(clknet_0_net589),
    .X(clknet_1_0__leaf_net589));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net589 (.A(clknet_0_net589),
    .X(clknet_1_1__leaf_net589));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net591 (.A(net591),
    .X(clknet_0_net591));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net591 (.A(clknet_0_net591),
    .X(clknet_1_0__leaf_net591));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net591 (.A(clknet_0_net591),
    .X(clknet_1_1__leaf_net591));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net590 (.A(net590),
    .X(clknet_0_net590));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net590 (.A(clknet_0_net590),
    .X(clknet_1_0__leaf_net590));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net590 (.A(clknet_0_net590),
    .X(clknet_1_1__leaf_net590));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net576 (.A(net576),
    .X(clknet_0_net576));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net576 (.A(clknet_0_net576),
    .X(clknet_1_0__leaf_net576));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net576 (.A(clknet_0_net576),
    .X(clknet_1_1__leaf_net576));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net575 (.A(net575),
    .X(clknet_0_net575));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net575 (.A(clknet_0_net575),
    .X(clknet_1_0__leaf_net575));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net575 (.A(clknet_0_net575),
    .X(clknet_1_1__leaf_net575));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net574 (.A(net574),
    .X(clknet_0_net574));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net574 (.A(clknet_0_net574),
    .X(clknet_1_0__leaf_net574));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net574 (.A(clknet_0_net574),
    .X(clknet_1_1__leaf_net574));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net573 (.A(net573),
    .X(clknet_0_net573));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net573 (.A(clknet_0_net573),
    .X(clknet_1_0__leaf_net573));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net573 (.A(clknet_0_net573),
    .X(clknet_1_1__leaf_net573));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net460 (.A(net460),
    .X(clknet_0_net460));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net460 (.A(clknet_0_net460),
    .X(clknet_1_0__leaf_net460));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net460 (.A(clknet_0_net460),
    .X(clknet_1_1__leaf_net460));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net467 (.A(net467),
    .X(clknet_0_net467));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net467 (.A(clknet_0_net467),
    .X(clknet_1_0__leaf_net467));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net467 (.A(clknet_0_net467),
    .X(clknet_1_1__leaf_net467));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net463 (.A(net463),
    .X(clknet_0_net463));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net463 (.A(clknet_0_net463),
    .X(clknet_1_0__leaf_net463));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net463 (.A(clknet_0_net463),
    .X(clknet_1_1__leaf_net463));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net461 (.A(net461),
    .X(clknet_0_net461));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net461 (.A(clknet_0_net461),
    .X(clknet_1_0__leaf_net461));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net461 (.A(clknet_0_net461),
    .X(clknet_1_1__leaf_net461));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net462 (.A(net462),
    .X(clknet_0_net462));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net462 (.A(clknet_0_net462),
    .X(clknet_1_0__leaf_net462));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net462 (.A(clknet_0_net462),
    .X(clknet_1_1__leaf_net462));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net371 (.A(net371),
    .X(clknet_0_net371));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net371 (.A(clknet_0_net371),
    .X(clknet_1_0__leaf_net371));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net371 (.A(clknet_0_net371),
    .X(clknet_1_1__leaf_net371));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net380 (.A(net380),
    .X(clknet_0_net380));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net380 (.A(clknet_0_net380),
    .X(clknet_1_0__leaf_net380));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net380 (.A(clknet_0_net380),
    .X(clknet_1_1__leaf_net380));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net375 (.A(net375),
    .X(clknet_0_net375));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net375 (.A(clknet_0_net375),
    .X(clknet_1_0__leaf_net375));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net375 (.A(clknet_0_net375),
    .X(clknet_1_1__leaf_net375));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net373 (.A(net373),
    .X(clknet_0_net373));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net373 (.A(clknet_0_net373),
    .X(clknet_1_0__leaf_net373));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net373 (.A(clknet_0_net373),
    .X(clknet_1_1__leaf_net373));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net736 (.A(net736),
    .X(clknet_0_net736));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net736 (.A(clknet_0_net736),
    .X(clknet_1_0__leaf_net736));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net736 (.A(clknet_0_net736),
    .X(clknet_1_1__leaf_net736));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net668 (.A(net668),
    .X(clknet_0_net668));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net668 (.A(clknet_0_net668),
    .X(clknet_1_0__leaf_net668));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net668 (.A(clknet_0_net668),
    .X(clknet_1_1__leaf_net668));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net396 (.A(net396),
    .X(clknet_0_net396));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net396 (.A(clknet_0_net396),
    .X(clknet_1_0__leaf_net396));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net396 (.A(clknet_0_net396),
    .X(clknet_1_1__leaf_net396));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net403 (.A(net403),
    .X(clknet_0_net403));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net403 (.A(clknet_0_net403),
    .X(clknet_1_0__leaf_net403));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net403 (.A(clknet_0_net403),
    .X(clknet_1_1__leaf_net403));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net406 (.A(net406),
    .X(clknet_0_net406));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net406 (.A(clknet_0_net406),
    .X(clknet_1_0__leaf_net406));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net406 (.A(clknet_0_net406),
    .X(clknet_1_1__leaf_net406));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net411 (.A(net411),
    .X(clknet_0_net411));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net411 (.A(clknet_0_net411),
    .X(clknet_1_0__leaf_net411));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net411 (.A(clknet_0_net411),
    .X(clknet_1_1__leaf_net411));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net412 (.A(net412),
    .X(clknet_0_net412));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net412 (.A(clknet_0_net412),
    .X(clknet_1_0__leaf_net412));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net412 (.A(clknet_0_net412),
    .X(clknet_1_1__leaf_net412));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net410 (.A(net410),
    .X(clknet_0_net410));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net410 (.A(clknet_0_net410),
    .X(clknet_1_0__leaf_net410));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net410 (.A(clknet_0_net410),
    .X(clknet_1_1__leaf_net410));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net415 (.A(net415),
    .X(clknet_0_net415));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net415 (.A(clknet_0_net415),
    .X(clknet_1_0__leaf_net415));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net415 (.A(clknet_0_net415),
    .X(clknet_1_1__leaf_net415));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net408 (.A(net408),
    .X(clknet_0_net408));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net408 (.A(clknet_0_net408),
    .X(clknet_1_0__leaf_net408));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net408 (.A(clknet_0_net408),
    .X(clknet_1_1__leaf_net408));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net407 (.A(net407),
    .X(clknet_0_net407));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net407 (.A(clknet_0_net407),
    .X(clknet_1_0__leaf_net407));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net407 (.A(clknet_0_net407),
    .X(clknet_1_1__leaf_net407));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net401 (.A(net401),
    .X(clknet_0_net401));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net401 (.A(clknet_0_net401),
    .X(clknet_1_0__leaf_net401));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net401 (.A(clknet_0_net401),
    .X(clknet_1_1__leaf_net401));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net430 (.A(net430),
    .X(clknet_0_net430));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net430 (.A(clknet_0_net430),
    .X(clknet_1_0__leaf_net430));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net430 (.A(clknet_0_net430),
    .X(clknet_1_1__leaf_net430));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net404 (.A(net404),
    .X(clknet_0_net404));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net404 (.A(clknet_0_net404),
    .X(clknet_1_0__leaf_net404));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net404 (.A(clknet_0_net404),
    .X(clknet_1_1__leaf_net404));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net402 (.A(net402),
    .X(clknet_0_net402));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net402 (.A(clknet_0_net402),
    .X(clknet_1_0__leaf_net402));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net402 (.A(clknet_0_net402),
    .X(clknet_1_1__leaf_net402));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net400 (.A(net400),
    .X(clknet_0_net400));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net400 (.A(clknet_0_net400),
    .X(clknet_1_0__leaf_net400));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net400 (.A(clknet_0_net400),
    .X(clknet_1_1__leaf_net400));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net399 (.A(net399),
    .X(clknet_0_net399));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net399 (.A(clknet_0_net399),
    .X(clknet_1_0__leaf_net399));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net399 (.A(clknet_0_net399),
    .X(clknet_1_1__leaf_net399));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net398 (.A(net398),
    .X(clknet_0_net398));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net398 (.A(clknet_0_net398),
    .X(clknet_1_0__leaf_net398));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net398 (.A(clknet_0_net398),
    .X(clknet_1_1__leaf_net398));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net397 (.A(net397),
    .X(clknet_0_net397));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net397 (.A(clknet_0_net397),
    .X(clknet_1_0__leaf_net397));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net397 (.A(clknet_0_net397),
    .X(clknet_1_1__leaf_net397));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net394 (.A(net394),
    .X(clknet_0_net394));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net394 (.A(clknet_0_net394),
    .X(clknet_1_0__leaf_net394));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net394 (.A(clknet_0_net394),
    .X(clknet_1_1__leaf_net394));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net395 (.A(net395),
    .X(clknet_0_net395));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net395 (.A(clknet_0_net395),
    .X(clknet_1_0__leaf_net395));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net395 (.A(clknet_0_net395),
    .X(clknet_1_1__leaf_net395));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net299 (.A(net299),
    .X(clknet_0_net299));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net299 (.A(clknet_0_net299),
    .X(clknet_1_0__leaf_net299));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net299 (.A(clknet_0_net299),
    .X(clknet_1_1__leaf_net299));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net288 (.A(net288),
    .X(clknet_0_net288));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net288 (.A(clknet_0_net288),
    .X(clknet_1_0__leaf_net288));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net288 (.A(clknet_0_net288),
    .X(clknet_1_1__leaf_net288));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net297 (.A(net297),
    .X(clknet_0_net297));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net297 (.A(clknet_0_net297),
    .X(clknet_1_0__leaf_net297));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net297 (.A(clknet_0_net297),
    .X(clknet_1_1__leaf_net297));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net296 (.A(net296),
    .X(clknet_0_net296));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net296 (.A(clknet_0_net296),
    .X(clknet_1_0__leaf_net296));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net296 (.A(clknet_0_net296),
    .X(clknet_1_1__leaf_net296));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net294 (.A(net294),
    .X(clknet_0_net294));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net294 (.A(clknet_0_net294),
    .X(clknet_1_0__leaf_net294));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net294 (.A(clknet_0_net294),
    .X(clknet_1_1__leaf_net294));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net292 (.A(net292),
    .X(clknet_0_net292));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net292 (.A(clknet_0_net292),
    .X(clknet_1_0__leaf_net292));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net292 (.A(net939),
    .X(clknet_1_1__leaf_net292));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net295 (.A(net295),
    .X(clknet_0_net295));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net295 (.A(clknet_0_net295),
    .X(clknet_1_0__leaf_net295));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net295 (.A(clknet_0_net295),
    .X(clknet_1_1__leaf_net295));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net291 (.A(net291),
    .X(clknet_0_net291));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net291 (.A(clknet_0_net291),
    .X(clknet_1_0__leaf_net291));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net291 (.A(clknet_0_net291),
    .X(clknet_1_1__leaf_net291));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net289 (.A(net289),
    .X(clknet_0_net289));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net289 (.A(clknet_0_net289),
    .X(clknet_1_0__leaf_net289));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net289 (.A(clknet_0_net289),
    .X(clknet_1_1__leaf_net289));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net290 (.A(net290),
    .X(clknet_0_net290));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net290 (.A(clknet_0_net290),
    .X(clknet_1_0__leaf_net290));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net290 (.A(clknet_0_net290),
    .X(clknet_1_1__leaf_net290));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net910 (.A(net910),
    .X(clknet_0_net910));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net910 (.A(clknet_0_net910),
    .X(clknet_1_0__leaf_net910));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net910 (.A(clknet_0_net910),
    .X(clknet_1_1__leaf_net910));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net311 (.A(net311),
    .X(clknet_0_net311));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net311 (.A(clknet_0_net311),
    .X(clknet_1_0__leaf_net311));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net311 (.A(clknet_0_net311),
    .X(clknet_1_1__leaf_net311));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net305 (.A(net305),
    .X(clknet_0_net305));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net305 (.A(clknet_0_net305),
    .X(clknet_1_0__leaf_net305));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net305 (.A(clknet_0_net305),
    .X(clknet_1_1__leaf_net305));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net306 (.A(net306),
    .X(clknet_0_net306));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net306 (.A(clknet_0_net306),
    .X(clknet_1_0__leaf_net306));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net306 (.A(clknet_0_net306),
    .X(clknet_1_1__leaf_net306));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net312 (.A(net312),
    .X(clknet_0_net312));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net312 (.A(clknet_0_net312),
    .X(clknet_1_0__leaf_net312));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net312 (.A(clknet_0_net312),
    .X(clknet_1_1__leaf_net312));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net308 (.A(net308),
    .X(clknet_0_net308));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net308 (.A(clknet_0_net308),
    .X(clknet_1_0__leaf_net308));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net308 (.A(clknet_0_net308),
    .X(clknet_1_1__leaf_net308));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net314 (.A(net314),
    .X(clknet_0_net314));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net314 (.A(clknet_0_net314),
    .X(clknet_1_0__leaf_net314));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net314 (.A(clknet_0_net314),
    .X(clknet_1_1__leaf_net314));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net317 (.A(net317),
    .X(clknet_0_net317));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net317 (.A(clknet_0_net317),
    .X(clknet_1_0__leaf_net317));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net317 (.A(clknet_0_net317),
    .X(clknet_1_1__leaf_net317));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net303 (.A(net303),
    .X(clknet_0_net303));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net303 (.A(clknet_0_net303),
    .X(clknet_1_0__leaf_net303));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net303 (.A(clknet_0_net303),
    .X(clknet_1_1__leaf_net303));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net310 (.A(net310),
    .X(clknet_0_net310));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net310 (.A(clknet_0_net310),
    .X(clknet_1_0__leaf_net310));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net310 (.A(clknet_0_net310),
    .X(clknet_1_1__leaf_net310));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net307 (.A(net307),
    .X(clknet_0_net307));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net307 (.A(clknet_0_net307),
    .X(clknet_1_0__leaf_net307));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net307 (.A(clknet_0_net307),
    .X(clknet_1_1__leaf_net307));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net372 (.A(net372),
    .X(clknet_0_net372));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net372 (.A(clknet_0_net372),
    .X(clknet_1_0__leaf_net372));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net372 (.A(clknet_0_net372),
    .X(clknet_1_1__leaf_net372));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net386 (.A(net386),
    .X(clknet_0_net386));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net386 (.A(clknet_0_net386),
    .X(clknet_1_0__leaf_net386));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net386 (.A(clknet_0_net386),
    .X(clknet_1_1__leaf_net386));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net367 (.A(net367),
    .X(clknet_0_net367));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net367 (.A(clknet_0_net367),
    .X(clknet_1_0__leaf_net367));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net367 (.A(clknet_0_net367),
    .X(clknet_1_1__leaf_net367));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net381 (.A(net381),
    .X(clknet_0_net381));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net381 (.A(clknet_0_net381),
    .X(clknet_1_0__leaf_net381));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net381 (.A(clknet_0_net381),
    .X(clknet_1_1__leaf_net381));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net358 (.A(net358),
    .X(clknet_0_net358));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net358 (.A(clknet_0_net358),
    .X(clknet_1_0__leaf_net358));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net358 (.A(clknet_0_net358),
    .X(clknet_1_1__leaf_net358));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net357 (.A(net357),
    .X(clknet_0_net357));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net357 (.A(clknet_0_net357),
    .X(clknet_1_0__leaf_net357));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net357 (.A(clknet_0_net357),
    .X(clknet_1_1__leaf_net357));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net352 (.A(net352),
    .X(clknet_0_net352));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net352 (.A(clknet_0_net352),
    .X(clknet_1_0__leaf_net352));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net352 (.A(clknet_0_net352),
    .X(clknet_1_1__leaf_net352));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net351 (.A(net351),
    .X(clknet_0_net351));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net351 (.A(clknet_0_net351),
    .X(clknet_1_0__leaf_net351));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net351 (.A(clknet_0_net351),
    .X(clknet_1_1__leaf_net351));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net350 (.A(net350),
    .X(clknet_0_net350));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net350 (.A(clknet_0_net350),
    .X(clknet_1_0__leaf_net350));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net350 (.A(clknet_0_net350),
    .X(clknet_1_1__leaf_net350));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net354 (.A(net354),
    .X(clknet_0_net354));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net354 (.A(clknet_0_net354),
    .X(clknet_1_0__leaf_net354));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net354 (.A(clknet_0_net354),
    .X(clknet_1_1__leaf_net354));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net356 (.A(net356),
    .X(clknet_0_net356));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net356 (.A(clknet_0_net356),
    .X(clknet_1_0__leaf_net356));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net356 (.A(clknet_0_net356),
    .X(clknet_1_1__leaf_net356));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net353 (.A(net353),
    .X(clknet_0_net353));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net353 (.A(clknet_0_net353),
    .X(clknet_1_0__leaf_net353));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net353 (.A(clknet_0_net353),
    .X(clknet_1_1__leaf_net353));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net355 (.A(net355),
    .X(clknet_0_net355));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net355 (.A(clknet_0_net355),
    .X(clknet_1_0__leaf_net355));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net355 (.A(clknet_0_net355),
    .X(clknet_1_1__leaf_net355));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net349 (.A(net349),
    .X(clknet_0_net349));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net349 (.A(clknet_0_net349),
    .X(clknet_1_0__leaf_net349));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net349 (.A(clknet_0_net349),
    .X(clknet_1_1__leaf_net349));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net368 (.A(net368),
    .X(clknet_0_net368));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net368 (.A(clknet_0_net368),
    .X(clknet_1_0__leaf_net368));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net368 (.A(clknet_0_net368),
    .X(clknet_1_1__leaf_net368));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net376 (.A(net376),
    .X(clknet_0_net376));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net376 (.A(clknet_0_net376),
    .X(clknet_1_0__leaf_net376));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net376 (.A(clknet_0_net376),
    .X(clknet_1_1__leaf_net376));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net347 (.A(net347),
    .X(clknet_0_net347));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net347 (.A(clknet_0_net347),
    .X(clknet_1_0__leaf_net347));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net347 (.A(clknet_0_net347),
    .X(clknet_1_1__leaf_net347));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net787 (.A(net787),
    .X(clknet_0_net787));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net787 (.A(clknet_0_net787),
    .X(clknet_1_0__leaf_net787));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net787 (.A(clknet_0_net787),
    .X(clknet_1_1__leaf_net787));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net342 (.A(net342),
    .X(clknet_0_net342));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net342 (.A(clknet_0_net342),
    .X(clknet_1_0__leaf_net342));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net342 (.A(clknet_0_net342),
    .X(clknet_1_1__leaf_net342));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net786 (.A(net786),
    .X(clknet_0_net786));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net786 (.A(clknet_0_net786),
    .X(clknet_1_0__leaf_net786));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net786 (.A(clknet_0_net786),
    .X(clknet_1_1__leaf_net786));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net341 (.A(net341),
    .X(clknet_0_net341));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net341 (.A(clknet_0_net341),
    .X(clknet_1_0__leaf_net341));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net341 (.A(clknet_0_net341),
    .X(clknet_1_1__leaf_net341));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net769 (.A(net769),
    .X(clknet_0_net769));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net769 (.A(clknet_0_net769),
    .X(clknet_1_0__leaf_net769));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net769 (.A(clknet_0_net769),
    .X(clknet_1_1__leaf_net769));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net302 (.A(net302),
    .X(clknet_0_net302));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net302 (.A(clknet_0_net302),
    .X(clknet_1_0__leaf_net302));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net302 (.A(clknet_0_net302),
    .X(clknet_1_1__leaf_net302));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net737 (.A(net737),
    .X(clknet_0_net737));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net737 (.A(clknet_0_net737),
    .X(clknet_1_0__leaf_net737));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net737 (.A(clknet_0_net737),
    .X(clknet_1_1__leaf_net737));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net169 (.A(net169),
    .X(clknet_0_net169));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net169 (.A(clknet_0_net169),
    .X(clknet_1_0__leaf_net169));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net169 (.A(clknet_0_net169),
    .X(clknet_1_1__leaf_net169));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net176 (.A(net176),
    .X(clknet_0_net176));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net176 (.A(clknet_0_net176),
    .X(clknet_1_0__leaf_net176));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net176 (.A(clknet_0_net176),
    .X(clknet_1_1__leaf_net176));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net192 (.A(net192),
    .X(clknet_0_net192));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net192 (.A(clknet_0_net192),
    .X(clknet_1_0__leaf_net192));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net192 (.A(clknet_0_net192),
    .X(clknet_1_1__leaf_net192));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net166 (.A(net166),
    .X(clknet_0_net166));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net166 (.A(clknet_0_net166),
    .X(clknet_1_0__leaf_net166));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net166 (.A(clknet_0_net166),
    .X(clknet_1_1__leaf_net166));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net175 (.A(net175),
    .X(clknet_0_net175));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net175 (.A(clknet_0_net175),
    .X(clknet_1_0__leaf_net175));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net175 (.A(clknet_0_net175),
    .X(clknet_1_1__leaf_net175));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net180 (.A(net180),
    .X(clknet_0_net180));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net180 (.A(clknet_0_net180),
    .X(clknet_1_0__leaf_net180));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net180 (.A(clknet_0_net180),
    .X(clknet_1_1__leaf_net180));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net168 (.A(net168),
    .X(clknet_0_net168));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net168 (.A(clknet_0_net168),
    .X(clknet_1_0__leaf_net168));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net168 (.A(clknet_0_net168),
    .X(clknet_1_1__leaf_net168));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net768 (.A(net768),
    .X(clknet_0_net768));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net768 (.A(clknet_0_net768),
    .X(clknet_1_0__leaf_net768));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net768 (.A(clknet_0_net768),
    .X(clknet_1_1__leaf_net768));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net158 (.A(net158),
    .X(clknet_0_net158));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net158 (.A(clknet_0_net158),
    .X(clknet_1_0__leaf_net158));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net158 (.A(clknet_0_net158),
    .X(clknet_1_1__leaf_net158));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net157 (.A(net157),
    .X(clknet_0_net157));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net157 (.A(clknet_0_net157),
    .X(clknet_1_0__leaf_net157));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net157 (.A(clknet_0_net157),
    .X(clknet_1_1__leaf_net157));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net767 (.A(net767),
    .X(clknet_0_net767));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net767 (.A(clknet_0_net767),
    .X(clknet_1_0__leaf_net767));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net767 (.A(clknet_0_net767),
    .X(clknet_1_1__leaf_net767));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net256 (.A(net256),
    .X(clknet_0_net256));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net256 (.A(clknet_0_net256),
    .X(clknet_1_0__leaf_net256));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net256 (.A(clknet_0_net256),
    .X(clknet_1_1__leaf_net256));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net270 (.A(net270),
    .X(clknet_0_net270));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net270 (.A(clknet_0_net270),
    .X(clknet_1_0__leaf_net270));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net270 (.A(clknet_0_net270),
    .X(clknet_1_1__leaf_net270));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net257 (.A(net257),
    .X(clknet_0_net257));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net257 (.A(clknet_0_net257),
    .X(clknet_1_0__leaf_net257));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net257 (.A(clknet_0_net257),
    .X(clknet_1_1__leaf_net257));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net134 (.A(net134),
    .X(clknet_0_net134));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net134 (.A(clknet_0_net134),
    .X(clknet_1_0__leaf_net134));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net134 (.A(clknet_0_net134),
    .X(clknet_1_1__leaf_net134));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net133 (.A(net133),
    .X(clknet_0_net133));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net133 (.A(clknet_0_net133),
    .X(clknet_1_0__leaf_net133));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net133 (.A(clknet_0_net133),
    .X(clknet_1_1__leaf_net133));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net735 (.A(net735),
    .X(clknet_0_net735));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net735 (.A(clknet_0_net735),
    .X(clknet_1_0__leaf_net735));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net735 (.A(clknet_0_net735),
    .X(clknet_1_1__leaf_net735));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net118 (.A(net118),
    .X(clknet_0_net118));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net118 (.A(clknet_0_net118),
    .X(clknet_1_0__leaf_net118));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net118 (.A(clknet_0_net118),
    .X(clknet_1_1__leaf_net118));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net119 (.A(net119),
    .X(clknet_0_net119));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net119 (.A(clknet_0_net119),
    .X(clknet_1_0__leaf_net119));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net119 (.A(clknet_0_net119),
    .X(clknet_1_1__leaf_net119));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net117 (.A(net117),
    .X(clknet_0_net117));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net117 (.A(clknet_0_net117),
    .X(clknet_1_0__leaf_net117));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net117 (.A(clknet_0_net117),
    .X(clknet_1_1__leaf_net117));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net128 (.A(net128),
    .X(clknet_0_net128));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net128 (.A(clknet_0_net128),
    .X(clknet_1_0__leaf_net128));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net128 (.A(clknet_0_net128),
    .X(clknet_1_1__leaf_net128));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer1 (.A(net147),
    .X(net935));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer2 (.A(net147),
    .X(net936));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer3 (.A(net920),
    .X(net937));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer4 (.A(net937),
    .X(net938));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer5 (.A(clknet_0_net292),
    .X(net939));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer6 (.A(net942),
    .X(net940));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer7 (.A(net940),
    .X(net941));
 sky130_fd_sc_hd__clkbuf_1 clone8 (.A(net144),
    .X(net942));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(net383),
    .X(net943));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(net799),
    .X(net944));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(net126),
    .X(net945));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(net464),
    .X(net946));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(net122),
    .X(net947));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(net805),
    .X(net948));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(net240),
    .X(net949));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(net814),
    .X(net950));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(net744),
    .X(net951));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(net369),
    .X(net952));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(in40),
    .X(net953));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(net237),
    .X(net954));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(net524),
    .X(net955));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(net198),
    .X(net956));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(net757),
    .X(net957));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(net934),
    .X(net958));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(net764),
    .X(net959));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(net244),
    .X(net960));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(net765),
    .X(net961));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(net774),
    .X(net962));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(net763),
    .X(net963));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(net742),
    .X(net964));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(net820),
    .X(net965));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(net374),
    .X(net966));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(net809),
    .X(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_A (.DIODE(clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(in0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(in1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(in10));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(in11));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(in12));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(in13));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(in14));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(in15));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(in16));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(in17));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(in18));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(in19));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(in2));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(in20));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(in21));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(in22));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(in23));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(in24));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(in25));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(in26));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(in27));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_A (.DIODE(in28));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_A (.DIODE(in29));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_A (.DIODE(in3));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_A (.DIODE(in30));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_A (.DIODE(in31));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_A (.DIODE(in32));
 sky130_fd_sc_hd__diode_2 ANTENNA_input28_A (.DIODE(in33));
 sky130_fd_sc_hd__diode_2 ANTENNA_input29_A (.DIODE(in34));
 sky130_fd_sc_hd__diode_2 ANTENNA_input30_A (.DIODE(in35));
 sky130_fd_sc_hd__diode_2 ANTENNA_input31_A (.DIODE(in36));
 sky130_fd_sc_hd__diode_2 ANTENNA_input32_A (.DIODE(in37));
 sky130_fd_sc_hd__diode_2 ANTENNA_input33_A (.DIODE(in38));
 sky130_fd_sc_hd__diode_2 ANTENNA_input34_A (.DIODE(in39));
 sky130_fd_sc_hd__diode_2 ANTENNA_input35_A (.DIODE(in4));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold19_A (.DIODE(in40));
 sky130_fd_sc_hd__diode_2 ANTENNA_input37_A (.DIODE(in41));
 sky130_fd_sc_hd__diode_2 ANTENNA_input38_A (.DIODE(in42));
 sky130_fd_sc_hd__diode_2 ANTENNA_input39_A (.DIODE(in43));
 sky130_fd_sc_hd__diode_2 ANTENNA_input40_A (.DIODE(in44));
 sky130_fd_sc_hd__diode_2 ANTENNA_input41_A (.DIODE(in45));
 sky130_fd_sc_hd__diode_2 ANTENNA_input42_A (.DIODE(in46));
 sky130_fd_sc_hd__diode_2 ANTENNA_input43_A (.DIODE(in47));
 sky130_fd_sc_hd__diode_2 ANTENNA_input44_A (.DIODE(in48));
 sky130_fd_sc_hd__diode_2 ANTENNA_input45_A (.DIODE(in49));
 sky130_fd_sc_hd__diode_2 ANTENNA_input46_A (.DIODE(in5));
 sky130_fd_sc_hd__diode_2 ANTENNA_input47_A (.DIODE(in50));
 sky130_fd_sc_hd__diode_2 ANTENNA_input48_A (.DIODE(in51));
 sky130_fd_sc_hd__diode_2 ANTENNA_input49_A (.DIODE(in52));
 sky130_fd_sc_hd__diode_2 ANTENNA_input50_A (.DIODE(in53));
 sky130_fd_sc_hd__diode_2 ANTENNA_input51_A (.DIODE(in54));
 sky130_fd_sc_hd__diode_2 ANTENNA_input52_A (.DIODE(in55));
 sky130_fd_sc_hd__diode_2 ANTENNA_input53_A (.DIODE(in56));
 sky130_fd_sc_hd__diode_2 ANTENNA_input54_A (.DIODE(in57));
 sky130_fd_sc_hd__diode_2 ANTENNA_input55_A (.DIODE(in58));
 sky130_fd_sc_hd__diode_2 ANTENNA_input56_A (.DIODE(in59));
 sky130_fd_sc_hd__diode_2 ANTENNA_input57_A (.DIODE(in6));
 sky130_fd_sc_hd__diode_2 ANTENNA_input58_A (.DIODE(in60));
 sky130_fd_sc_hd__diode_2 ANTENNA_input59_A (.DIODE(in61));
 sky130_fd_sc_hd__diode_2 ANTENNA_input60_A (.DIODE(in7));
 sky130_fd_sc_hd__diode_2 ANTENNA_input61_A (.DIODE(in8));
 sky130_fd_sc_hd__diode_2 ANTENNA_input62_A (.DIODE(in9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_B (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_B (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_B (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c286_C (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_D (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_B (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_A (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_S1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_A2 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_A1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_X (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge769_C_N (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_SCE (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_S1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_X (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge793_C_N (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge789_S0 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge783_SCD (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge770_A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge767_D_N (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_S0 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_C1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c191_S1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_SET_B (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_X (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge784_B1 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge781_C_N (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_Q_N (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge778_D_N (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge772_D (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_A0 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA_c393_SCD (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA_c236_A2 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA_c235_A2 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA_c231_S1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_X (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge796_S0 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA_c238_A1 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA_c237_A2 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA_c235_A3 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA_c234_D1 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_C_N (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA_c232_B (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA_c231_A0 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA_c229_X (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout92_A (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA_c398_B (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_A (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA_c264_X (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge783_SCE (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA_c458_A3 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_B (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_A (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_A1 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA_c323_A0 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_X (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_B (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_B (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_A (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_A2 (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_c344_A2 (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_C_N (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_c340_S0 (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_X (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout91_A (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA_c413_B1 (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA_c664_B (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_A (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_X (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge786_A1 (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_B (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_B (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_A (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_B (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_X (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge794_A3 (.DIODE(net595));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge787_A3 (.DIODE(net595));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_A2 (.DIODE(net595));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_A2 (.DIODE(net595));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_X (.DIODE(net595));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge794_A0 (.DIODE(net599));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_B (.DIODE(net599));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_A3 (.DIODE(net599));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_SET_B (.DIODE(net599));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_RESET_B (.DIODE(net599));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_C (.DIODE(net599));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_C1 (.DIODE(net599));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_C (.DIODE(net599));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_SCD (.DIODE(net599));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_X (.DIODE(net599));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge779_X (.DIODE(net678));
 sky130_fd_sc_hd__diode_2 ANTENNA_c311_A (.DIODE(net678));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_A (.DIODE(net678));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge818_RESET_B (.DIODE(net686));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge786_X (.DIODE(net686));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge801_Q (.DIODE(net704));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_S1 (.DIODE(net704));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_D_N (.DIODE(net704));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_A (.DIODE(net704));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_A (.DIODE(net704));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_S1 (.DIODE(net729));
 sky130_fd_sc_hd__diode_2 ANTENNA_c611_SCE (.DIODE(net729));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_D1 (.DIODE(net729));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_C (.DIODE(net729));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_C (.DIODE(net729));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_B (.DIODE(net729));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_A (.DIODE(net729));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_D1 (.DIODE(net729));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout103_A (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_S1 (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_C (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA_s875_Q (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge789_A2 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge782_A3 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_c286_B (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_C (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_A1 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_A3 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_B1 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_C1 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_B (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_c159_B (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_c158_X (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_output69_A (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_s864_Q (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_C (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_B (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c395_D1 (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c392_D_N (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_output78_A (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_s862_Q (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_C (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_C (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c394_S1 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c392_C_N (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c370_S0 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c368_S1 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c365_S1 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer3_A (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout90_X (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_C (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_D1 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_A (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c215_S0 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_C (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c208_B (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge784_D1 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout92_X (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_c402_C (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_c278_S0 (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_c270_A (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge776_SCD (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_c269_B (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_c267_A (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_c266_B (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_c265_A (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_A1 (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_A (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout98_X (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_B1 (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c397_B (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c528_A (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout97_A (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_A (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c264_B (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout99_X (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_A (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c83_S0 (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c81_A2 (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c80_D1 (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c79_B (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c73_D_N (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c72_C (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c71_C (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c212_S1 (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c88_B (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout103_X (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_SCE (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge768_C_N (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c664_C (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c663_B (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c661_B (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c660_B (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_C (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_B (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_B (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c548_S1 (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_15_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_14_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_13_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_12_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_11_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_10_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_9_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_8_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_7_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_6_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_5_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_4_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_3_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_2_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_1_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_0_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_X (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_CLK_N (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c295_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c297_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge820_GATE (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge833_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge837_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s846_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s847_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s848_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s857_GATE_N (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s858_GATE (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s859_SLEEP_B (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_1_0_clk_X (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_CLK_N (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_CLK_N (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c190_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_CLK_N (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge798_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge826_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge841_GATE_N (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s849_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s850_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_2_0_clk_X (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_CLK_N (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge783_CLK_N (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge805_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge832_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge834_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge836_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s860_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s861_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s896_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s900_GATE_N (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_3_0_clk_X (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c563_CLK_N (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge809_GATE_N (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge810_GATE_N (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge814_GATE_N (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s865_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s866_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s867_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s868_GATE_N (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s875_SLEEP_B (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_4_0_clk_X (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c366_CLK_N (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge799_CLK_N (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge816_GATE_N (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge828_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge830_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge831_CLK_N (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s844_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s852_GATE_N (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s853_GATE_N (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_8_0_clk_X (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c253_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c256_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c393_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge802_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge803_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge811_GATE (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge839_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s851_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s854_GATE (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s855_GATE_N (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s856_GATE_N (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s864_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_10_0_clk_X (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c761_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge795_CLK_N (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge800_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge818_GATE_N (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge838_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge842_GATE_N (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s863_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s894_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s895_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s898_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_11_0_clk_X (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_CLK_N (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_CLK_N (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_CLK_N (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge780_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge801_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s869_GATE_N (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s893_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s902_GATE (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_12_0_clk_X (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_CLK_N (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c720_CLK_N (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge807_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge825_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s880_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s890_GATE (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s891_SLEEP_B (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s892_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_13_0_clk_X (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_A2 (.DIODE(clknet_1_1__leaf_net359));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_A1 (.DIODE(clknet_1_1__leaf_net359));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_A2 (.DIODE(clknet_1_1__leaf_net359));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_B1 (.DIODE(clknet_1_1__leaf_net359));
 sky130_fd_sc_hd__diode_2 ANTENNA_c554_D_N (.DIODE(clknet_1_1__leaf_net359));
 sky130_fd_sc_hd__diode_2 ANTENNA_c558_SET_B (.DIODE(clknet_1_1__leaf_net359));
 sky130_fd_sc_hd__diode_2 ANTENNA_c559_A1 (.DIODE(clknet_1_1__leaf_net359));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_B (.DIODE(clknet_1_1__leaf_net359));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net359_X (.DIODE(clknet_1_1__leaf_net359));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_D_N (.DIODE(clknet_1_0__leaf_net575));
 sky130_fd_sc_hd__diode_2 ANTENNA_c693_RESET_B (.DIODE(clknet_1_0__leaf_net575));
 sky130_fd_sc_hd__diode_2 ANTENNA_c695_SET_B (.DIODE(clknet_1_0__leaf_net575));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge774_SCD (.DIODE(clknet_1_0__leaf_net575));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge787_S0 (.DIODE(clknet_1_0__leaf_net575));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge791_RESET_B (.DIODE(clknet_1_0__leaf_net575));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net575_X (.DIODE(clknet_1_0__leaf_net575));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_DE (.DIODE(clknet_1_0__leaf_net373));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_D1 (.DIODE(clknet_1_0__leaf_net373));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_SCD (.DIODE(clknet_1_0__leaf_net373));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge766_A2 (.DIODE(clknet_1_0__leaf_net373));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge786_A2 (.DIODE(clknet_1_0__leaf_net373));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge792_A3 (.DIODE(clknet_1_0__leaf_net373));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net373_X (.DIODE(clknet_1_0__leaf_net373));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_B (.DIODE(clknet_1_1__leaf_net401));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_C1 (.DIODE(clknet_1_1__leaf_net401));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_B (.DIODE(clknet_1_1__leaf_net401));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_C_N (.DIODE(clknet_1_1__leaf_net401));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_D_N (.DIODE(clknet_1_1__leaf_net401));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_D_N (.DIODE(clknet_1_1__leaf_net401));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_S0 (.DIODE(clknet_1_1__leaf_net401));
 sky130_fd_sc_hd__diode_2 ANTENNA_c502_S0 (.DIODE(clknet_1_1__leaf_net401));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_A1 (.DIODE(clknet_1_1__leaf_net401));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net401_X (.DIODE(clknet_1_1__leaf_net401));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_A (.DIODE(clknet_1_1__leaf_net290));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_A (.DIODE(clknet_1_1__leaf_net290));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_C1 (.DIODE(clknet_1_1__leaf_net290));
 sky130_fd_sc_hd__diode_2 ANTENNA_c394_A2 (.DIODE(clknet_1_1__leaf_net290));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net290_X (.DIODE(clknet_1_1__leaf_net290));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_A2 (.DIODE(clknet_1_1__leaf_net270));
 sky130_fd_sc_hd__diode_2 ANTENNA_c344_D1 (.DIODE(clknet_1_1__leaf_net270));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_A3 (.DIODE(clknet_1_1__leaf_net270));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_D1 (.DIODE(clknet_1_1__leaf_net270));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge792_A2 (.DIODE(clknet_1_1__leaf_net270));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net270_X (.DIODE(clknet_1_1__leaf_net270));
 sky130_fd_sc_hd__clkbuf_1 clone1 (.A(net148),
    .X(net968));
 sky130_fd_sc_hd__and3_1 clone2 (.A(net970),
    .B(net280),
    .C(net282),
    .X(net969));
 sky130_fd_sc_hd__clkbuf_1 clone3 (.A(net148),
    .X(net970));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_301 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_282 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_554 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_8 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_25 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_280 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_580 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_8 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_20 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_355 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_395 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_568 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_450 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_527 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_58 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_359 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_8 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_188 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_8 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_511 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_168 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_31 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_254 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_8 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_188 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_582 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_78 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_8 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_624 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_547 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_572 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_572 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_20 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_310 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_20 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_17 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_245 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_385 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_230 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_582 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_312 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_578 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_170 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_546 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_497 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_441 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_617 ();
endmodule
