module netlist_1 (clk,
    in0,
    in1,
    in10,
    in11,
    in12,
    in13,
    in14,
    in15,
    in16,
    in17,
    in18,
    in19,
    in2,
    in20,
    in21,
    in22,
    in23,
    in24,
    in25,
    in26,
    in27,
    in28,
    in29,
    in3,
    in30,
    in31,
    in32,
    in33,
    in34,
    in35,
    in36,
    in37,
    in38,
    in39,
    in4,
    in40,
    in41,
    in42,
    in43,
    in44,
    in45,
    in46,
    in47,
    in48,
    in49,
    in5,
    in50,
    in51,
    in52,
    in53,
    in54,
    in55,
    in56,
    in57,
    in58,
    in59,
    in6,
    in60,
    in61,
    in62,
    in63,
    in64,
    in65,
    in66,
    in67,
    in68,
    in69,
    in7,
    in70,
    in71,
    in72,
    in73,
    in74,
    in75,
    in76,
    in77,
    in78,
    in79,
    in8,
    in80,
    in81,
    in82,
    in83,
    in84,
    in85,
    in86,
    in87,
    in88,
    in89,
    in9,
    in90,
    in91,
    in92,
    in93,
    in94,
    in95,
    in96,
    in97,
    in98,
    in99,
    out0,
    out1,
    out10,
    out11,
    out12,
    out13,
    out14,
    out15,
    out16,
    out17,
    out18,
    out19,
    out2,
    out20,
    out21,
    out22,
    out23,
    out24,
    out25,
    out26,
    out27,
    out28,
    out29,
    out3,
    out30,
    out31,
    out32,
    out33,
    out34,
    out35,
    out36,
    out37,
    out38,
    out39,
    out4,
    out40,
    out41,
    out42,
    out43,
    out44,
    out45,
    out46,
    out47,
    out48,
    out49,
    out5,
    out50,
    out51,
    out52,
    out53,
    out54,
    out55,
    out56,
    out57,
    out58,
    out59,
    out6,
    out60,
    out61,
    out62,
    out63,
    out64,
    out65,
    out66,
    out67,
    out68,
    out69,
    out7,
    out70,
    out71,
    out72,
    out73,
    out74,
    out75,
    out76,
    out77,
    out78,
    out79,
    out8,
    out80,
    out81,
    out82,
    out83,
    out84,
    out85,
    out86,
    out87,
    out88,
    out89,
    out9,
    out90,
    out91,
    out92,
    out93,
    out94,
    out95,
    out96,
    out97,
    out98,
    out99,
    rst);
 input clk;
 input in0;
 input in1;
 input in10;
 input in11;
 input in12;
 input in13;
 input in14;
 input in15;
 input in16;
 input in17;
 input in18;
 input in19;
 input in2;
 input in20;
 input in21;
 input in22;
 input in23;
 input in24;
 input in25;
 input in26;
 input in27;
 input in28;
 input in29;
 input in3;
 input in30;
 input in31;
 input in32;
 input in33;
 input in34;
 input in35;
 input in36;
 input in37;
 input in38;
 input in39;
 input in4;
 input in40;
 input in41;
 input in42;
 input in43;
 input in44;
 input in45;
 input in46;
 input in47;
 input in48;
 input in49;
 input in5;
 input in50;
 input in51;
 input in52;
 input in53;
 input in54;
 input in55;
 input in56;
 input in57;
 input in58;
 input in59;
 input in6;
 input in60;
 input in61;
 input in62;
 input in63;
 input in64;
 input in65;
 input in66;
 input in67;
 input in68;
 input in69;
 input in7;
 input in70;
 input in71;
 input in72;
 input in73;
 input in74;
 input in75;
 input in76;
 input in77;
 input in78;
 input in79;
 input in8;
 input in80;
 input in81;
 input in82;
 input in83;
 input in84;
 input in85;
 input in86;
 input in87;
 input in88;
 input in89;
 input in9;
 input in90;
 input in91;
 input in92;
 input in93;
 input in94;
 input in95;
 input in96;
 input in97;
 input in98;
 input in99;
 output out0;
 output out1;
 output out10;
 output out11;
 output out12;
 output out13;
 output out14;
 output out15;
 output out16;
 output out17;
 output out18;
 output out19;
 output out2;
 output out20;
 output out21;
 output out22;
 output out23;
 output out24;
 output out25;
 output out26;
 output out27;
 output out28;
 output out29;
 output out3;
 output out30;
 output out31;
 output out32;
 output out33;
 output out34;
 output out35;
 output out36;
 output out37;
 output out38;
 output out39;
 output out4;
 output out40;
 output out41;
 output out42;
 output out43;
 output out44;
 output out45;
 output out46;
 output out47;
 output out48;
 output out49;
 output out5;
 output out50;
 output out51;
 output out52;
 output out53;
 output out54;
 output out55;
 output out56;
 output out57;
 output out58;
 output out59;
 output out6;
 output out60;
 output out61;
 output out62;
 output out63;
 output out64;
 output out65;
 output out66;
 output out67;
 output out68;
 output out69;
 output out7;
 output out70;
 output out71;
 output out72;
 output out73;
 output out74;
 output out75;
 output out76;
 output out77;
 output out78;
 output out79;
 output out8;
 output out80;
 output out81;
 output out82;
 output out83;
 output out84;
 output out85;
 output out86;
 output out87;
 output out88;
 output out89;
 output out9;
 output out90;
 output out91;
 output out92;
 output out93;
 output out94;
 output out95;
 output out96;
 output out97;
 output out98;
 output out99;
 input rst;

 wire net0;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net63;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net64;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net65;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net66;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net67;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net68;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net69;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net7;
 wire net70;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net71;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net72;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net73;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net74;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net75;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net76;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net77;
 wire net770;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net484;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_0_net753;
 wire clknet_1_0__leaf_net753;
 wire clknet_1_1__leaf_net753;
 wire clknet_0_net517;
 wire clknet_1_0__leaf_net517;
 wire clknet_1_1__leaf_net517;
 wire clknet_0_net522;
 wire clknet_1_0__leaf_net522;
 wire clknet_1_1__leaf_net522;
 wire clknet_0_net412;
 wire clknet_1_0__leaf_net412;
 wire clknet_1_1__leaf_net412;
 wire clknet_0_net411;
 wire clknet_1_0__leaf_net411;
 wire clknet_1_1__leaf_net411;
 wire clknet_0_net407;
 wire clknet_1_0__leaf_net407;
 wire clknet_1_1__leaf_net407;
 wire clknet_0_net549;
 wire clknet_1_0__leaf_net549;
 wire clknet_1_1__leaf_net549;
 wire clknet_0_net752;
 wire clknet_1_0__leaf_net752;
 wire clknet_1_1__leaf_net752;
 wire clknet_0_net409;
 wire clknet_1_0__leaf_net409;
 wire clknet_1_1__leaf_net409;
 wire clknet_0_net403;
 wire clknet_1_0__leaf_net403;
 wire clknet_1_1__leaf_net403;
 wire clknet_0_net413;
 wire clknet_1_0__leaf_net413;
 wire clknet_1_1__leaf_net413;
 wire clknet_0_net751;
 wire clknet_1_0__leaf_net751;
 wire clknet_1_1__leaf_net751;
 wire clknet_0_net410;
 wire clknet_1_0__leaf_net410;
 wire clknet_1_1__leaf_net410;
 wire clknet_0_net392;
 wire clknet_1_0__leaf_net392;
 wire clknet_1_1__leaf_net392;
 wire clknet_0_net496;
 wire clknet_1_0__leaf_net496;
 wire clknet_1_1__leaf_net496;
 wire clknet_0_net939;
 wire clknet_1_0__leaf_net939;
 wire clknet_1_1__leaf_net939;
 wire clknet_0_net735;
 wire clknet_1_0__leaf_net735;
 wire clknet_1_1__leaf_net735;
 wire clknet_0_net310;
 wire clknet_1_0__leaf_net310;
 wire clknet_1_1__leaf_net310;
 wire clknet_0_net307;
 wire clknet_1_0__leaf_net307;
 wire clknet_1_1__leaf_net307;
 wire clknet_0_net905;
 wire clknet_1_0__leaf_net905;
 wire clknet_1_1__leaf_net905;
 wire clknet_0_net908;
 wire clknet_1_0__leaf_net908;
 wire clknet_1_1__leaf_net908;
 wire clknet_0_net296;
 wire clknet_1_0__leaf_net296;
 wire clknet_1_1__leaf_net296;
 wire clknet_0_net904;
 wire clknet_1_0__leaf_net904;
 wire clknet_1_1__leaf_net904;
 wire clknet_0_net394;
 wire clknet_1_0__leaf_net394;
 wire clknet_1_1__leaf_net394;
 wire clknet_0_net734;
 wire clknet_1_0__leaf_net734;
 wire clknet_1_1__leaf_net734;
 wire clknet_0_net733;
 wire clknet_1_0__leaf_net733;
 wire clknet_1_1__leaf_net733;
 wire clknet_0_net714;
 wire clknet_1_0__leaf_net714;
 wire clknet_1_1__leaf_net714;
 wire clknet_0_net460;
 wire clknet_1_0__leaf_net460;
 wire clknet_1_1__leaf_net460;
 wire clknet_0_net504;
 wire clknet_1_0__leaf_net504;
 wire clknet_1_1__leaf_net504;
 wire clknet_0_net462;
 wire clknet_1_0__leaf_net462;
 wire clknet_1_1__leaf_net462;
 wire clknet_0_net458;
 wire clknet_1_0__leaf_net458;
 wire clknet_1_1__leaf_net458;
 wire clknet_0_net641;
 wire clknet_1_0__leaf_net641;
 wire clknet_1_1__leaf_net641;
 wire clknet_0_net518;
 wire clknet_1_0__leaf_net518;
 wire clknet_1_1__leaf_net518;
 wire clknet_0_net509;
 wire clknet_1_0__leaf_net509;
 wire clknet_1_1__leaf_net509;
 wire clknet_0_net260;
 wire clknet_1_0__leaf_net260;
 wire clknet_1_1__leaf_net260;
 wire clknet_0_net893;
 wire clknet_1_0__leaf_net893;
 wire clknet_1_1__leaf_net893;
 wire clknet_0_net401;
 wire clknet_1_0__leaf_net401;
 wire clknet_1_1__leaf_net401;
 wire clknet_0_net713;
 wire clknet_1_0__leaf_net713;
 wire clknet_1_1__leaf_net713;
 wire clknet_0_net405;
 wire clknet_1_0__leaf_net405;
 wire clknet_1_1__leaf_net405;
 wire clknet_0_net336;
 wire clknet_1_0__leaf_net336;
 wire clknet_1_1__leaf_net336;
 wire clknet_0_net894;
 wire clknet_1_0__leaf_net894;
 wire clknet_1_1__leaf_net894;
 wire clknet_0_net277;
 wire clknet_1_0__leaf_net277;
 wire clknet_1_1__leaf_net277;
 wire clknet_0_net422;
 wire clknet_1_0__leaf_net422;
 wire clknet_1_1__leaf_net422;
 wire clknet_0_net373;
 wire clknet_1_0__leaf_net373;
 wire clknet_1_1__leaf_net373;
 wire clknet_0_net378;
 wire clknet_1_0__leaf_net378;
 wire clknet_1_1__leaf_net378;
 wire clknet_0_net898;
 wire clknet_1_0__leaf_net898;
 wire clknet_1_1__leaf_net898;
 wire clknet_0_net712;
 wire clknet_1_0__leaf_net712;
 wire clknet_1_1__leaf_net712;
 wire clknet_0_net512;
 wire clknet_1_0__leaf_net512;
 wire clknet_1_1__leaf_net512;
 wire clknet_0_net465;
 wire clknet_1_0__leaf_net465;
 wire clknet_1_1__leaf_net465;
 wire clknet_0_net346;
 wire clknet_1_0__leaf_net346;
 wire clknet_1_1__leaf_net346;
 wire clknet_0_net616;
 wire clknet_1_0__leaf_net616;
 wire clknet_1_1__leaf_net616;
 wire clknet_0_net354;
 wire clknet_1_0__leaf_net354;
 wire clknet_1_1__leaf_net354;
 wire clknet_0_net615;
 wire clknet_1_0__leaf_net615;
 wire clknet_1_1__leaf_net615;
 wire clknet_0_net390;
 wire clknet_1_0__leaf_net390;
 wire clknet_1_1__leaf_net390;
 wire clknet_0_net353;
 wire clknet_1_0__leaf_net353;
 wire clknet_1_1__leaf_net353;
 wire clknet_0_net273;
 wire clknet_1_0__leaf_net273;
 wire clknet_1_1__leaf_net273;
 wire clknet_0_net379;
 wire clknet_1_0__leaf_net379;
 wire clknet_1_1__leaf_net379;
 wire clknet_0_net276;
 wire clknet_1_0__leaf_net276;
 wire clknet_1_1__leaf_net276;
 wire clknet_0_net247;
 wire clknet_1_0__leaf_net247;
 wire clknet_1_1__leaf_net247;
 wire clknet_0_net695;
 wire clknet_1_0__leaf_net695;
 wire clknet_1_1__leaf_net695;
 wire clknet_0_net377;
 wire clknet_1_0__leaf_net377;
 wire clknet_1_1__leaf_net377;
 wire clknet_0_net399;
 wire clknet_1_0__leaf_net399;
 wire clknet_1_1__leaf_net399;
 wire clknet_0_net502;
 wire clknet_1_0__leaf_net502;
 wire clknet_1_1__leaf_net502;
 wire clknet_0_net532;
 wire clknet_1_0__leaf_net532;
 wire clknet_1_1__leaf_net532;
 wire clknet_0_net535;
 wire clknet_1_0__leaf_net535;
 wire clknet_1_1__leaf_net535;
 wire clknet_0_net167;
 wire clknet_1_0__leaf_net167;
 wire clknet_1_1__leaf_net167;
 wire clknet_0_net191;
 wire clknet_1_0__leaf_net191;
 wire clknet_1_1__leaf_net191;
 wire clknet_0_net887;
 wire clknet_1_0__leaf_net887;
 wire clknet_1_1__leaf_net887;
 wire clknet_0_net312;
 wire clknet_1_0__leaf_net312;
 wire clknet_1_1__leaf_net312;
 wire clknet_0_net168;
 wire clknet_1_0__leaf_net168;
 wire clknet_1_1__leaf_net168;
 wire clknet_0_net161;
 wire clknet_1_0__leaf_net161;
 wire clknet_1_1__leaf_net161;
 wire clknet_0_net263;
 wire clknet_1_0__leaf_net263;
 wire clknet_1_1__leaf_net263;
 wire clknet_0_net166;
 wire clknet_1_0__leaf_net166;
 wire clknet_1_1__leaf_net166;
 wire clknet_0_net283;
 wire clknet_1_0__leaf_net283;
 wire clknet_1_1__leaf_net283;
 wire clknet_0_net302;
 wire clknet_1_0__leaf_net302;
 wire clknet_1_1__leaf_net302;
 wire clknet_0_net178;
 wire clknet_1_0__leaf_net178;
 wire clknet_1_1__leaf_net178;
 wire clknet_0_net505;
 wire clknet_1_0__leaf_net505;
 wire clknet_1_1__leaf_net505;
 wire clknet_0_net922;
 wire clknet_1_0__leaf_net922;
 wire clknet_1_1__leaf_net922;
 wire clknet_0_net179;
 wire clknet_1_0__leaf_net179;
 wire clknet_1_1__leaf_net179;
 wire clknet_0_net613;
 wire clknet_1_0__leaf_net613;
 wire clknet_1_1__leaf_net613;
 wire clknet_0_net218;
 wire clknet_1_0__leaf_net218;
 wire clknet_1_1__leaf_net218;
 wire clknet_0_net219;
 wire clknet_1_0__leaf_net219;
 wire clknet_1_1__leaf_net219;
 wire clknet_0_net694;
 wire clknet_1_0__leaf_net694;
 wire clknet_1_1__leaf_net694;
 wire clknet_0_net935;
 wire clknet_1_0__leaf_net935;
 wire clknet_1_1__leaf_net935;
 wire clknet_0_net693;
 wire clknet_1_0__leaf_net693;
 wire clknet_1_1__leaf_net693;
 wire clknet_0_net895;
 wire clknet_1_0__leaf_net895;
 wire clknet_1_1__leaf_net895;
 wire clknet_0_net157;
 wire clknet_1_0__leaf_net157;
 wire clknet_1_1__leaf_net157;
 wire clknet_0_net293;
 wire clknet_1_0__leaf_net293;
 wire clknet_1_1__leaf_net293;
 wire clknet_0_net295;
 wire clknet_1_0__leaf_net295;
 wire clknet_1_1__leaf_net295;
 wire clknet_0_net900;
 wire clknet_1_0__leaf_net900;
 wire clknet_1_1__leaf_net900;
 wire clknet_0_net675;
 wire clknet_1_0__leaf_net675;
 wire clknet_1_1__leaf_net675;
 wire clknet_0_net284;
 wire clknet_1_0__leaf_net284;
 wire clknet_1_1__leaf_net284;
 wire clknet_0_net104;
 wire clknet_1_0__leaf_net104;
 wire clknet_1_1__leaf_net104;
 wire clknet_0_net890;
 wire clknet_1_0__leaf_net890;
 wire clknet_1_1__leaf_net890;
 wire clknet_0_net231;
 wire clknet_1_0__leaf_net231;
 wire clknet_1_1__leaf_net231;
 wire clknet_0_net333;
 wire clknet_1_0__leaf_net333;
 wire clknet_1_1__leaf_net333;
 wire clknet_0_net221;
 wire clknet_1_0__leaf_net221;
 wire clknet_1_1__leaf_net221;
 wire clknet_0_net674;
 wire clknet_1_0__leaf_net674;
 wire clknet_1_1__leaf_net674;
 wire clknet_0_net318;
 wire clknet_1_0__leaf_net318;
 wire clknet_1_1__leaf_net318;
 wire clknet_0_net199;
 wire clknet_1_0__leaf_net199;
 wire clknet_1_1__leaf_net199;
 wire clknet_0_net98;
 wire clknet_1_0__leaf_net98;
 wire clknet_1_1__leaf_net98;
 wire clknet_0_net100;
 wire clknet_1_0__leaf_net100;
 wire clknet_1_1__leaf_net100;
 wire clknet_0_net193;
 wire clknet_1_0__leaf_net193;
 wire clknet_1_1__leaf_net193;
 wire clknet_0_net916;
 wire clknet_1_0__leaf_net916;
 wire clknet_1_1__leaf_net916;
 wire clknet_0_net73;
 wire clknet_1_0__leaf_net73;
 wire clknet_1_1__leaf_net73;
 wire clknet_0_net530;
 wire clknet_1_0__leaf_net530;
 wire clknet_1_1__leaf_net530;
 wire clknet_0_net76;
 wire clknet_1_0__leaf_net76;
 wire clknet_1_1__leaf_net76;
 wire clknet_0_net182;
 wire clknet_1_0__leaf_net182;
 wire clknet_1_1__leaf_net182;
 wire clknet_0_net186;
 wire clknet_1_0__leaf_net186;
 wire clknet_1_1__leaf_net186;
 wire clknet_0_net78;
 wire clknet_1_0__leaf_net78;
 wire clknet_1_1__leaf_net78;
 wire clknet_0_net84;
 wire clknet_1_0__leaf_net84;
 wire clknet_1_1__leaf_net84;
 wire clknet_0_net938;
 wire clknet_1_0__leaf_net938;
 wire clknet_1_1__leaf_net938;
 wire clknet_0_net109;
 wire clknet_1_0__leaf_net109;
 wire clknet_1_1__leaf_net109;
 wire clknet_0_net651;
 wire clknet_1_0__leaf_net651;
 wire clknet_1_1__leaf_net651;
 wire clknet_0_net328;
 wire clknet_1_0__leaf_net328;
 wire clknet_1_1__leaf_net328;
 wire clknet_0_net113;
 wire clknet_1_0__leaf_net113;
 wire clknet_1_1__leaf_net113;
 wire clknet_0_net116;
 wire clknet_1_0__leaf_net116;
 wire clknet_1_1__leaf_net116;
 wire clknet_0_net923;
 wire clknet_1_0__leaf_net923;
 wire clknet_1_1__leaf_net923;
 wire clknet_0_net111;
 wire clknet_1_0__leaf_net111;
 wire clknet_1_1__leaf_net111;
 wire clknet_0_net83;
 wire clknet_1_0__leaf_net83;
 wire clknet_1_1__leaf_net83;
 wire clknet_0_net936;
 wire clknet_1_0__leaf_net936;
 wire clknet_1_1__leaf_net936;
 wire clknet_0_net79;
 wire clknet_1_0__leaf_net79;
 wire clknet_1_1__leaf_net79;
 wire clknet_0_net70;
 wire clknet_1_0__leaf_net70;
 wire clknet_1_1__leaf_net70;
 wire clknet_0_net74;
 wire clknet_1_0__leaf_net74;
 wire clknet_1_1__leaf_net74;
 wire clknet_0_net285;
 wire clknet_1_0__leaf_net285;
 wire clknet_1_1__leaf_net285;
 wire clknet_0_net72;
 wire clknet_1_0__leaf_net72;
 wire clknet_1_1__leaf_net72;
 wire clknet_0_net202;
 wire clknet_1_0__leaf_net202;
 wire clknet_1_1__leaf_net202;
 wire clknet_0_net208;
 wire clknet_1_0__leaf_net208;
 wire clknet_1_1__leaf_net208;
 wire clknet_0_net75;
 wire clknet_1_0__leaf_net75;
 wire clknet_1_1__leaf_net75;
 wire clknet_0_net77;
 wire clknet_1_0__leaf_net77;
 wire clknet_1_1__leaf_net77;
 wire clknet_0_net184;
 wire clknet_1_0__leaf_net184;
 wire clknet_1_1__leaf_net184;
 wire clknet_0_net288;
 wire clknet_1_0__leaf_net288;
 wire clknet_1_1__leaf_net288;
 wire clknet_0_net175;
 wire clknet_1_0__leaf_net175;
 wire clknet_1_1__leaf_net175;
 wire clknet_0_net673;
 wire clknet_1_0__leaf_net673;
 wire clknet_1_1__leaf_net673;
 wire clknet_0_net66;
 wire clknet_1_0__leaf_net66;
 wire clknet_1_1__leaf_net66;
 wire clknet_0_net174;
 wire clknet_1_0__leaf_net174;
 wire clknet_1_1__leaf_net174;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1108;

 sky130_fd_sc_hd__mux4_2 c100 (.A0(net861),
    .A1(net867),
    .A2(net833),
    .A3(net827),
    .S0(net1000),
    .S1(net863),
    .X(net0));
 sky130_fd_sc_hd__mux4_2 c101 (.A0(net843),
    .A1(net832),
    .A2(net864),
    .A3(net1082),
    .S0(net838),
    .S1(net1000),
    .X(net1));
 sky130_fd_sc_hd__mux4_2 c102 (.A0(net857),
    .A1(net833),
    .A2(net796),
    .A3(net864),
    .S0(net1000),
    .S1(net834),
    .X(net917));
 sky130_fd_sc_hd__mux4_2 c103 (.A0(net1000),
    .A1(net869),
    .A2(net828),
    .A3(net838),
    .S0(net853),
    .S1(net999),
    .X(net2));
 sky130_fd_sc_hd__mux4_2 c104 (.A0(net868),
    .A1(net862),
    .A2(net839),
    .A3(net1000),
    .S0(net999),
    .S1(net822),
    .X(net3));
 sky130_fd_sc_hd__mux4_1 c105 (.A0(net858),
    .A1(net831),
    .A2(net838),
    .A3(net832),
    .S0(net1021),
    .S1(net0),
    .X(net4));
 sky130_fd_sc_hd__mux4_2 c106 (.A0(net4),
    .A1(net866),
    .A2(net864),
    .A3(net1000),
    .S0(net999),
    .S1(net831),
    .X(net5));
 sky130_fd_sc_hd__mux4_2 c107 (.A0(net5),
    .A1(net1000),
    .A2(net1082),
    .A3(net866),
    .S0(net837),
    .S1(net857),
    .X(net6));
 sky130_fd_sc_hd__mux4_2 c108 (.A0(net3),
    .A1(net0),
    .A2(net4),
    .A3(net1000),
    .S0(net840),
    .S1(net5),
    .X(net7));
 sky130_fd_sc_hd__mux4_2 c109 (.A0(net863),
    .A1(net860),
    .A2(net7),
    .A3(net813),
    .S0(net1000),
    .S1(net5),
    .X(net918));
 sky130_fd_sc_hd__a2111o_1 c110 (.A1(net1000),
    .A2(net817),
    .B1(net837),
    .C1(net1060),
    .D1(net1002),
    .X(net943));
 sky130_fd_sc_hd__a2111o_1 c111 (.A1(net825),
    .A2(net1014),
    .B1(net917),
    .C1(net863),
    .D1(net1019),
    .X(net8));
 sky130_fd_sc_hd__a2111o_1 c112 (.A1(net837),
    .A2(net484),
    .B1(net1002),
    .C1(net1014),
    .D1(net1011),
    .X(net906));
 sky130_fd_sc_hd__a2111o_2 c113 (.A1(net834),
    .A2(net906),
    .B1(net843),
    .C1(net1019),
    .D1(net1002),
    .X(net9));
 sky130_fd_sc_hd__or4bb_1 c114 (.A(net785),
    .B(net828),
    .C_N(net834),
    .D_N(net6),
    .X(net932));
 sky130_fd_sc_hd__a2111o_1 c115 (.A1(net1009),
    .A2(net853),
    .B1(net790),
    .C1(net9),
    .D1(net1002),
    .X(net10));
 sky130_fd_sc_hd__a2111o_2 c116 (.A1(net4),
    .A2(net918),
    .B1(net863),
    .C1(net1029),
    .D1(net1014),
    .X(net11));
 sky130_fd_sc_hd__a2111o_1 c117 (.A1(net850),
    .A2(net11),
    .B1(net9),
    .C1(net834),
    .D1(net796),
    .X(net937));
 sky130_fd_sc_hd__a2111o_1 c118 (.A1(net10),
    .A2(net850),
    .B1(net866),
    .C1(net843),
    .D1(net1002),
    .X(net12));
 sky130_fd_sc_hd__a2111o_1 c119 (.A1(net1029),
    .A2(net11),
    .B1(net825),
    .C1(net865),
    .D1(net906),
    .X(net13));
 sky130_fd_sc_hd__a2111o_2 c120 (.A1(net794),
    .A2(net13),
    .B1(net862),
    .C1(net790),
    .D1(net937),
    .X(net910));
 sky130_fd_sc_hd__mux4_1 c121 (.A0(net853),
    .A1(net910),
    .A2(net794),
    .A3(net1019),
    .S0(net865),
    .S1(net807),
    .X(net929));
 sky130_fd_sc_hd__a2111o_1 c122 (.A1(net807),
    .A2(net825),
    .B1(net937),
    .C1(net943),
    .D1(net906),
    .X(net14));
 sky130_fd_sc_hd__a2111o_2 c123 (.A1(net9),
    .A2(net11),
    .B1(net943),
    .C1(net910),
    .D1(net929),
    .X(net946));
 sky130_fd_sc_hd__mux4_2 c124 (.A0(net14),
    .A1(net10),
    .A2(net929),
    .A3(net11),
    .S0(net9),
    .S1(net1009),
    .X(net880));
 sky130_fd_sc_hd__a2111o_1 c125 (.A1(net880),
    .A2(net11),
    .B1(net1060),
    .C1(net13),
    .D1(net14),
    .X(net15));
 sky130_fd_sc_hd__mux4_1 c126 (.A0(net15),
    .A1(net880),
    .A2(net937),
    .A3(net943),
    .S0(net11),
    .S1(net9),
    .X(net16));
 sky130_fd_sc_hd__mux4_2 c127 (.A0(net13),
    .A1(net880),
    .A2(net798),
    .A3(net946),
    .S0(net1009),
    .S1(net817),
    .X(net17));
 sky130_fd_sc_hd__mux4_1 c128 (.A0(net17),
    .A1(net932),
    .A2(net880),
    .A3(net865),
    .S0(net14),
    .S1(net16),
    .X(net944));
 sky130_fd_sc_hd__mux4_1 c129 (.A0(net863),
    .A1(net910),
    .A2(net17),
    .A3(net880),
    .S0(net1019),
    .S1(net1014),
    .X(net925));
 sky130_fd_sc_hd__mux4_1 c130 (.A0(net16),
    .A1(net880),
    .A2(net17),
    .A3(net865),
    .S0(net910),
    .S1(net925),
    .X(net926));
 sky130_fd_sc_hd__mux4_1 c131 (.A0(net12),
    .A1(net925),
    .A2(net926),
    .A3(net1014),
    .S0(net15),
    .S1(net17),
    .X(net947));
 sky130_fd_sc_hd__or4bb_4 c132 (.A(net1007),
    .B(net1084),
    .C_N(net1006),
    .D_N(net1011),
    .X(net18));
 sky130_fd_sc_hd__a2111o_2 c133 (.A1(net1026),
    .A2(net1081),
    .B1(net793),
    .C1(net1007),
    .D1(net998),
    .X(net19));
 sky130_fd_sc_hd__a2111o_2 c134 (.A1(net1027),
    .A2(net793),
    .B1(net1026),
    .C1(net1002),
    .D1(net1007),
    .X(net20));
 sky130_fd_sc_hd__mux4_2 c135 (.A0(net1007),
    .A1(net998),
    .A2(net1084),
    .A3(net1002),
    .S0(net1011),
    .S1(net1024),
    .X(net21));
 sky130_fd_sc_hd__a2111o_2 c136 (.A1(net1009),
    .A2(net837),
    .B1(net1079),
    .C1(net998),
    .D1(net997),
    .X(net22));
 sky130_fd_sc_hd__a2111o_4 c137 (.A1(net984),
    .A2(net1026),
    .B1(net998),
    .C1(net1080),
    .D1(net1011),
    .X(net23));
 sky130_fd_sc_hd__a2111o_4 c138 (.A1(net981),
    .A2(net1083),
    .B1(net1084),
    .C1(net1079),
    .D1(net1080),
    .X(net24));
 sky130_fd_sc_hd__mux4_2 c139 (.A0(net981),
    .A1(net1080),
    .A2(net982),
    .A3(net24),
    .S0(net997),
    .S1(net984),
    .X(net25));
 sky130_fd_sc_hd__mux4_2 c140 (.A0(net1084),
    .A1(net1082),
    .A2(net998),
    .A3(net771),
    .S0(net1007),
    .S1(net983),
    .X(net26));
 sky130_fd_sc_hd__mux4_2 c141 (.A0(net998),
    .A1(net26),
    .A2(net19),
    .A3(net1006),
    .S0(net24),
    .S1(net984),
    .X(net27));
 sky130_fd_sc_hd__mux4_2 c142 (.A0(net981),
    .A1(net1009),
    .A2(net1083),
    .A3(net1081),
    .S0(net984),
    .S1(net1026),
    .X(net934));
 sky130_fd_sc_hd__mux4_2 c143 (.A0(net1082),
    .A1(net1085),
    .A2(net1083),
    .A3(net1057),
    .S0(net27),
    .S1(net1079),
    .X(net28));
 sky130_fd_sc_hd__a2111o_2 c144 (.A1(net27),
    .A2(net26),
    .B1(net24),
    .C1(net997),
    .D1(net1079),
    .X(net29));
 sky130_fd_sc_hd__mux4_2 c145 (.A0(net25),
    .A1(net1011),
    .A2(net1057),
    .A3(net28),
    .S0(net1083),
    .S1(net1079),
    .X(net30));
 sky130_fd_sc_hd__mux4_2 c146 (.A0(net24),
    .A1(net484),
    .A2(net28),
    .A3(net26),
    .S0(net934),
    .S1(net1079),
    .X(net872));
 sky130_fd_sc_hd__mux4_2 c147 (.A0(net981),
    .A1(net1081),
    .A2(net28),
    .A3(net24),
    .S0(net26),
    .S1(net1079),
    .X(net31));
 sky130_fd_sc_hd__mux4_2 c148 (.A0(net975),
    .A1(net28),
    .A2(net1085),
    .A3(net1028),
    .S0(net978),
    .S1(net31),
    .X(net32));
 sky130_fd_sc_hd__a2111o_4 c149 (.A1(net31),
    .A2(net1001),
    .B1(net1081),
    .C1(net975),
    .D1(net1079),
    .X(net33));
 sky130_fd_sc_hd__mux4_2 c150 (.A0(net1026),
    .A1(net30),
    .A2(net973),
    .A3(net1029),
    .S0(net978),
    .S1(net986),
    .X(net34));
 sky130_fd_sc_hd__mux4_2 c151 (.A0(net978),
    .A1(net1037),
    .A2(net1084),
    .A3(net1079),
    .S0(net32),
    .S1(net971),
    .X(net885));
 sky130_fd_sc_hd__mux4_2 c152 (.A0(net934),
    .A1(net973),
    .A2(net974),
    .A3(net1057),
    .S0(net1054),
    .S1(net1007),
    .X(net35));
 sky130_fd_sc_hd__mux4_2 c153 (.A0(net969),
    .A1(net1037),
    .A2(net18),
    .A3(net1084),
    .S0(net35),
    .S1(net971),
    .X(net36));
 sky130_fd_sc_hd__a2111o_4 c154 (.A1(net36),
    .A2(net794),
    .B1(net805),
    .C1(net997),
    .D1(net787),
    .X(net37));
 sky130_fd_sc_hd__mux4_2 c155 (.A0(net963),
    .A1(net802),
    .A2(net1018),
    .A3(net1012),
    .S0(net795),
    .S1(net36),
    .X(net38));
 sky130_fd_sc_hd__a2111o_1 c156 (.A1(net805),
    .A2(net973),
    .B1(net793),
    .C1(net972),
    .D1(net1019),
    .X(net39));
 sky130_fd_sc_hd__a2111o_2 c157 (.A1(net38),
    .A2(net786),
    .B1(net36),
    .C1(net785),
    .D1(net790),
    .X(net40));
 sky130_fd_sc_hd__mux4_2 c158 (.A0(net40),
    .A1(net786),
    .A2(net1001),
    .A3(net794),
    .S0(net802),
    .S1(net1021),
    .X(net897));
 sky130_fd_sc_hd__a2111o_1 c159 (.A1(net800),
    .A2(net803),
    .B1(net1083),
    .C1(net958),
    .D1(net36),
    .X(net41));
 sky130_fd_sc_hd__a2111o_4 c160 (.A1(net968),
    .A2(net771),
    .B1(net800),
    .C1(net1021),
    .D1(net586),
    .X(net42));
 sky130_fd_sc_hd__sdfbbn_2 c161 (.CLK_N(clknet_4_4_0_clk),
    .D(net1081),
    .RESET_B(net978),
    .SCD(net1012),
    .SCE(net805),
    .SET_B(net958),
    .Q(net44),
    .Q_N(net43));
 sky130_fd_sc_hd__mux4_1 c162 (.A0(net1044),
    .A1(net38),
    .A2(net1018),
    .A3(net974),
    .S0(net968),
    .S1(net958),
    .X(net45));
 sky130_fd_sc_hd__mux4_2 c163 (.A0(net1060),
    .A1(net788),
    .A2(net807),
    .A3(net1054),
    .S0(net806),
    .S1(net963),
    .X(net46));
 sky130_fd_sc_hd__a2111o_1 c164 (.A1(net42),
    .A2(net40),
    .B1(net787),
    .C1(net1082),
    .D1(net586),
    .X(net47));
 sky130_fd_sc_hd__sdfbbn_2 c165 (.CLK_N(clknet_4_5_0_clk),
    .D(net802),
    .RESET_B(net955),
    .SCD(net795),
    .SCE(net958),
    .SET_B(net626),
    .Q(net49),
    .Q_N(net48));
 sky130_fd_sc_hd__mux4_1 c166 (.A0(net35),
    .A1(net803),
    .A2(net38),
    .A3(net955),
    .S0(net968),
    .X(net50));
 sky130_fd_sc_hd__mux4_1 c167 (.A0(net955),
    .A1(net790),
    .A2(net997),
    .A3(net958),
    .S0(net42),
    .S1(net626),
    .X(net51));
 sky130_fd_sc_hd__mux4_1 c168 (.A0(net974),
    .A1(net799),
    .A2(net39),
    .A3(net785),
    .S0(net955),
    .S1(net626),
    .X(net52));
 sky130_fd_sc_hd__mux4_2 c169 (.A0(net802),
    .A1(net42),
    .A2(net795),
    .A3(net963),
    .S0(net40),
    .S1(net586),
    .X(net53));
 sky130_fd_sc_hd__mux4_2 c170 (.A0(net1028),
    .A1(net40),
    .A2(net20),
    .A3(net793),
    .S0(net585),
    .S1(net623),
    .X(net54));
 sky130_fd_sc_hd__mux4_1 c171 (.A0(net786),
    .A1(net49),
    .A2(net1012),
    .A3(net955),
    .S0(net953),
    .S1(net586),
    .X(net55));
 sky130_fd_sc_hd__mux4_1 c172 (.A0(net803),
    .A1(net44),
    .A2(net46),
    .A3(net48),
    .S0(net953),
    .S1(net585),
    .X(net56));
 sky130_fd_sc_hd__mux4_1 c173 (.A0(net787),
    .A1(net46),
    .A2(net1010),
    .A3(net48),
    .S0(net955),
    .S1(net626),
    .X(net57));
 sky130_fd_sc_hd__mux4_1 c174 (.A0(net46),
    .A1(net793),
    .A2(net788),
    .A3(net955),
    .S0(net669),
    .S1(net671),
    .X(net58));
 sky130_fd_sc_hd__mux4_1 c175 (.A0(net953),
    .A1(net46),
    .A2(net585),
    .S0(net626),
    .S1(net672),
    .X(net59));
 sky130_fd_sc_hd__a2111o_4 c176 (.A1(net820),
    .A2(net818),
    .B1(net1029),
    .C1(net973),
    .D1(net828),
    .X(net60));
 sky130_fd_sc_hd__mux4_2 c177 (.A0(net823),
    .A1(net60),
    .A2(net797),
    .A3(net1035),
    .S0(net804),
    .S1(net812),
    .X(net61));
 sky130_fd_sc_hd__a2111o_2 c178 (.A1(net1035),
    .A2(net820),
    .B1(net831),
    .C1(net1009),
    .D1(net623),
    .X(net62));
 sky130_fd_sc_hd__mux4_1 c179 (.A0(net967),
    .A1(net820),
    .A2(net958),
    .A3(net60),
    .S0(net934),
    .S1(net956),
    .X(net63));
 sky130_fd_sc_hd__mux4_1 c180 (.A0(net811),
    .A1(net48),
    .A2(net62),
    .A3(net790),
    .S0(net955),
    .S1(net573),
    .X(net64));
 sky130_fd_sc_hd__mux4_1 c181 (.A0(net824),
    .A1(net62),
    .A2(net955),
    .A3(net1035),
    .S0(net954),
    .S1(net912),
    .X(net65));
 sky130_fd_sc_hd__mux4_1 c182 (.A0(net793),
    .A1(net788),
    .A2(net813),
    .A3(net816),
    .S0(net572),
    .S1(clknet_1_0__leaf_net673),
    .X(net66));
 sky130_fd_sc_hd__mux4_1 c183 (.A0(net1083),
    .A1(clknet_1_0__leaf_net66),
    .A2(net62),
    .A3(net958),
    .S0(net825),
    .S1(net912),
    .X(net67));
 sky130_fd_sc_hd__mux4_2 c184 (.A0(net816),
    .A1(net31),
    .A2(net1014),
    .A3(net48),
    .S0(net572),
    .S1(net623),
    .X(net68));
 sky130_fd_sc_hd__mux4_1 c185 (.A0(net794),
    .A1(net813),
    .A2(net967),
    .A3(net831),
    .S0(net956),
    .S1(net912),
    .X(net69));
 sky130_fd_sc_hd__mux4_2 c186 (.A0(clknet_1_0__leaf_net66),
    .A1(net816),
    .A2(net60),
    .A3(net788),
    .S0(net572),
    .S1(clknet_1_0__leaf_net674),
    .X(net70));
 sky130_fd_sc_hd__mux4_2 c187 (.A0(net798),
    .A1(net1015),
    .A2(net1014),
    .A3(net28),
    .S0(net816),
    .S1(net812),
    .X(net71));
 sky130_fd_sc_hd__mux4_2 c188 (.A0(net68),
    .A1(clknet_1_0__leaf_net70),
    .A2(net805),
    .A3(net823),
    .S0(net1080),
    .S1(net626),
    .X(net72));
 sky130_fd_sc_hd__mux4_1 c189 (.A0(clknet_1_0__leaf_net70),
    .A1(net824),
    .A2(net71),
    .A3(net808),
    .S0(clknet_1_0__leaf_net673),
    .S1(clknet_1_0__leaf_net674),
    .X(net73));
 sky130_fd_sc_hd__mux4_2 c190 (.A0(net71),
    .A1(clknet_1_1__leaf_net70),
    .A2(net974),
    .A3(net60),
    .S0(net820),
    .S1(net573),
    .X(net74));
 sky130_fd_sc_hd__mux4_2 c191 (.A0(net824),
    .A1(clknet_1_0__leaf_net72),
    .A2(net1021),
    .A3(net823),
    .S0(net68),
    .S1(clknet_1_0__leaf_net673),
    .X(net75));
 sky130_fd_sc_hd__mux4_1 c192 (.A0(net795),
    .A1(net816),
    .A2(clknet_1_0__leaf_net73),
    .A3(net670),
    .S0(net912),
    .S1(clknet_1_0__leaf_net673),
    .X(net76));
 sky130_fd_sc_hd__mux4_2 c193 (.A0(net60),
    .A1(net68),
    .A2(clknet_1_1__leaf_net75),
    .A3(net1015),
    .S0(net771),
    .S1(net623),
    .X(net77));
 sky130_fd_sc_hd__mux4_2 c194 (.A0(net46),
    .A1(clknet_1_0__leaf_net77),
    .A2(clknet_1_1__leaf_net75),
    .A3(clknet_1_0__leaf_net76),
    .S0(net573),
    .S1(clknet_1_0__leaf_net673),
    .X(net78));
 sky130_fd_sc_hd__mux4_2 c195 (.A0(clknet_1_0__leaf_net77),
    .A1(clknet_1_0__leaf_net74),
    .A2(clknet_1_0__leaf_net78),
    .A3(net1035),
    .S0(net980),
    .S1(net819),
    .X(net79));
 sky130_fd_sc_hd__mux4_1 c196 (.A0(clknet_1_0__leaf_net78),
    .A1(clknet_1_1__leaf_net70),
    .A2(net1009),
    .A3(clknet_1_1__leaf_net66),
    .S0(net829),
    .S1(net573),
    .X(net936));
 sky130_fd_sc_hd__mux4_1 c197 (.A0(net812),
    .A1(clknet_1_1__leaf_net936),
    .A2(clknet_1_0__leaf_net76),
    .A3(net967),
    .S0(net824),
    .S1(net626),
    .X(net80));
 sky130_fd_sc_hd__a2111o_4 c198 (.A1(net60),
    .A2(net817),
    .B1(net43),
    .C1(net809),
    .D1(net787),
    .X(net81));
 sky130_fd_sc_hd__mux4_1 c199 (.A0(net1009),
    .A1(net958),
    .A2(net81),
    .A3(net956),
    .S0(clknet_1_0__leaf_net936),
    .S1(net1015),
    .X(net82));
 sky130_fd_sc_hd__a2111o_1 c200 (.A1(net44),
    .A2(clknet_1_1__leaf_net78),
    .B1(net827),
    .C1(net798),
    .D1(net971),
    .X(net83));
 sky130_fd_sc_hd__a2111o_1 c201 (.A1(net819),
    .A2(net829),
    .B1(net846),
    .C1(net845),
    .D1(clknet_1_0__leaf_net78),
    .X(net84));
 sky130_fd_sc_hd__a2111o_2 c202 (.A1(net827),
    .A2(net838),
    .B1(net1060),
    .C1(net586),
    .D1(net626),
    .X(net85));
 sky130_fd_sc_hd__a2111o_2 c203 (.A1(net809),
    .A2(net841),
    .B1(net851),
    .C1(net1082),
    .D1(net671),
    .X(net86));
 sky130_fd_sc_hd__sdfbbp_1 c204 (.CLK(clknet_4_1_0_clk),
    .D(net849),
    .RESET_B(clknet_1_1__leaf_net83),
    .SCD(clknet_1_0__leaf_net84),
    .SCE(net978),
    .SET_B(net956),
    .Q(net88),
    .Q_N(net87));
 sky130_fd_sc_hd__mux4_1 c205 (.A0(clknet_1_0__leaf_net83),
    .A1(net840),
    .A2(clknet_1_0__leaf_net73),
    .A3(net1002),
    .S0(net85),
    .S1(clknet_1_0__leaf_net936),
    .X(net89));
 sky130_fd_sc_hd__a2111o_4 c206 (.A1(net81),
    .A2(net997),
    .B1(net854),
    .C1(net971),
    .D1(net977),
    .X(net90));
 sky130_fd_sc_hd__mux4_2 c207 (.A0(net788),
    .A1(net838),
    .A2(net484),
    .A3(net1016),
    .S0(net851),
    .S1(net81),
    .X(net91));
 sky130_fd_sc_hd__mux4_1 c208 (.A0(net484),
    .A1(net86),
    .A2(net85),
    .A3(clknet_1_0__leaf_net84),
    .S0(net827),
    .S1(net677),
    .X(net92));
 sky130_fd_sc_hd__mux4_1 c209 (.A0(net851),
    .A1(net88),
    .A2(clknet_1_1__leaf_net83),
    .A3(net62),
    .S0(net847),
    .S1(net1094),
    .X(net93));
 sky130_fd_sc_hd__a2111o_1 c210 (.A1(clknet_1_0__leaf_net84),
    .A2(net827),
    .B1(net91),
    .C1(net87),
    .D1(net85),
    .X(net94));
 sky130_fd_sc_hd__a2111o_2 c211 (.A1(net847),
    .A2(net977),
    .B1(net1029),
    .C1(net844),
    .D1(net681),
    .X(net896));
 sky130_fd_sc_hd__a2111o_2 c212 (.A1(net91),
    .A2(net997),
    .B1(net846),
    .C1(net626),
    .D1(net680),
    .X(net95));
 sky130_fd_sc_hd__mux4_1 c213 (.A0(net846),
    .A1(clknet_1_0__leaf_net84),
    .A2(net841),
    .A3(net88),
    .S0(net1009),
    .S1(net81),
    .X(net96));
 sky130_fd_sc_hd__a2111o_4 c214 (.A1(net829),
    .A2(net95),
    .B1(net980),
    .C1(net849),
    .D1(net570),
    .X(net97));
 sky130_fd_sc_hd__mux4_1 c215 (.A0(net997),
    .A1(net71),
    .A2(net1028),
    .A3(net807),
    .S0(net1014),
    .S1(clknet_1_0__leaf_net674),
    .X(net98));
 sky130_fd_sc_hd__mux4_1 c216 (.A0(clknet_1_0__leaf_net79),
    .A1(net97),
    .A2(net81),
    .A3(net43),
    .S0(clknet_1_0__leaf_net98),
    .S1(net623),
    .X(net99));
 sky130_fd_sc_hd__mux4_1 c217 (.A0(clknet_1_0__leaf_net98),
    .A1(net1006),
    .A2(net62),
    .A3(net90),
    .S0(net819),
    .S1(net97),
    .X(net100));
 sky130_fd_sc_hd__a2111o_1 c218 (.A1(net62),
    .A2(clknet_1_0__leaf_net100),
    .B1(net97),
    .C1(net570),
    .D1(net607),
    .X(net916));
 sky130_fd_sc_hd__a2111o_1 c219 (.A1(clknet_1_0__leaf_net72),
    .A2(clknet_1_1__leaf_net916),
    .B1(net87),
    .C1(net97),
    .D1(net679),
    .X(net101));
 sky130_fd_sc_hd__mux4_1 c220 (.A0(net839),
    .A1(net813),
    .A2(clknet_1_0__leaf_net79),
    .A3(net980),
    .S0(net832),
    .S1(net607),
    .X(net102));
 sky130_fd_sc_hd__mux4_1 c221 (.A0(net97),
    .A1(net839),
    .A2(net1015),
    .A3(net831),
    .S0(net671),
    .S1(net672),
    .X(net924));
 sky130_fd_sc_hd__mux4_1 c222 (.A0(net864),
    .A1(net958),
    .A2(net862),
    .A3(net956),
    .S0(net95),
    .S1(net980),
    .X(net103));
 sky130_fd_sc_hd__mux4_1 c223 (.A0(net807),
    .A1(net817),
    .A2(net1001),
    .A3(net999),
    .S0(net912),
    .S1(clknet_1_0__leaf_net675),
    .X(net104));
 sky130_fd_sc_hd__mux4_1 c224 (.A0(net831),
    .A1(clknet_1_0__leaf_net83),
    .A2(net0),
    .A3(net844),
    .S0(net832),
    .S1(net607),
    .X(net105));
 sky130_fd_sc_hd__mux4_1 c225 (.A0(net832),
    .A1(clknet_1_0__leaf_net75),
    .A2(net861),
    .A3(clknet_1_0__leaf_net84),
    .S0(net821),
    .S1(net607),
    .X(net106));
 sky130_fd_sc_hd__mux4_1 c226 (.A0(net6),
    .A1(net1021),
    .A2(net832),
    .A3(clknet_1_1__leaf_net936),
    .S0(net677),
    .S1(net682),
    .X(net107));
 sky130_fd_sc_hd__mux4_1 c227 (.A0(net813),
    .A1(clknet_1_0__leaf_net84),
    .A2(clknet_1_0__leaf_net75),
    .A3(net95),
    .S0(net835),
    .S1(net956),
    .X(net108));
 sky130_fd_sc_hd__a2111o_1 c228 (.A1(net6),
    .A2(net837),
    .B1(net629),
    .C1(clknet_1_0__leaf_net938),
    .D1(net680),
    .X(net923));
 sky130_fd_sc_hd__mux4_1 c229 (.A0(net1019),
    .A1(net1094),
    .A2(clknet_1_1__leaf_net923),
    .A3(net1001),
    .S0(net969),
    .S1(clknet_1_0__leaf_net938),
    .X(net109));
 sky130_fd_sc_hd__mux4_1 c230 (.A0(net95),
    .A1(net1021),
    .A2(net3),
    .A3(net785),
    .S0(net629),
    .S1(net679),
    .X(net110));
 sky130_fd_sc_hd__mux4_2 c231 (.A0(net963),
    .A1(net3),
    .A2(net999),
    .A3(net838),
    .S0(net942),
    .S1(net903),
    .X(net927));
 sky130_fd_sc_hd__mux4_1 c232 (.A0(net110),
    .A1(net801),
    .A2(net827),
    .A3(clknet_1_0__leaf_net923),
    .S0(net572),
    .S1(net607),
    .X(net111));
 sky130_fd_sc_hd__mux4_1 c233 (.A0(net844),
    .A1(net963),
    .A2(net999),
    .A3(net933),
    .S0(net572),
    .S1(net630),
    .X(net112));
 sky130_fd_sc_hd__mux4_1 c234 (.A0(net112),
    .A1(clknet_1_0__leaf_net109),
    .A2(net869),
    .A3(net861),
    .S0(net671),
    .S1(net682),
    .X(net113));
 sky130_fd_sc_hd__mux4_1 c235 (.A0(clknet_1_0__leaf_net113),
    .A1(net953),
    .A2(clknet_1_1__leaf_net109),
    .A3(net839),
    .S0(net680),
    .S1(net682),
    .X(net114));
 sky130_fd_sc_hd__mux4_1 c236 (.A0(net854),
    .A1(net1094),
    .A2(clknet_1_1__leaf_net109),
    .A3(net112),
    .S0(net95),
    .S1(net956),
    .X(net115));
 sky130_fd_sc_hd__mux4_1 c237 (.A0(net1016),
    .A1(net927),
    .A2(net862),
    .A3(clknet_1_1__leaf_net113),
    .S0(net110),
    .S1(net682),
    .X(net116));
 sky130_fd_sc_hd__mux4_1 c238 (.A0(clknet_1_0__leaf_net116),
    .A1(clknet_1_0__leaf_net104),
    .A2(net858),
    .A3(net71),
    .S0(net956),
    .S1(net607),
    .X(net117));
 sky130_fd_sc_hd__sdfbbn_2 c239 (.CLK_N(clknet_4_0_0_clk),
    .D(net801),
    .RESET_B(clknet_1_0__leaf_net116),
    .SCD(net860),
    .SCE(net630),
    .SET_B(clknet_1_0__leaf_net651),
    .Q(net119),
    .Q_N(net118));
 sky130_fd_sc_hd__mux4_1 c240 (.A0(clknet_1_0__leaf_net116),
    .A1(clknet_1_1__leaf_net109),
    .A2(net118),
    .A3(clknet_1_0__leaf_net70),
    .S0(clknet_1_0__leaf_net651),
    .S1(net677),
    .X(net120));
 sky130_fd_sc_hd__mux4_1 c241 (.A0(clknet_1_0__leaf_net109),
    .A1(net2),
    .A2(net118),
    .A3(clknet_1_0__leaf_net116),
    .S0(clknet_1_0__leaf_net651),
    .S1(net940),
    .X(net121));
 sky130_fd_sc_hd__mux4_1 c256 (.A0(net8),
    .A1(clknet_1_1__leaf_net936),
    .A2(net927),
    .A3(net11),
    .S0(net946),
    .S1(net572),
    .X(net122));
 sky130_fd_sc_hd__mux4_2 c257 (.A0(net1009),
    .A1(net946),
    .A2(net840),
    .A3(net969),
    .S0(net975),
    .S1(net630),
    .X(net914));
 sky130_fd_sc_hd__mux4_2 c258 (.A0(net845),
    .A1(net934),
    .A2(net975),
    .A3(net914),
    .S0(net825),
    .S1(net880),
    .X(net871));
 sky130_fd_sc_hd__mux4_1 c259 (.A0(net11),
    .A1(net484),
    .A2(net17),
    .A3(net927),
    .S0(net914),
    .S1(net871),
    .X(net941));
 sky130_fd_sc_hd__mux4_1 c260 (.A0(net1029),
    .A1(net934),
    .A2(net946),
    .A3(net871),
    .S0(net914),
    .S1(net907),
    .X(net892));
 sky130_fd_sc_hd__mux4_1 c261 (.A0(net796),
    .A1(net871),
    .A2(net947),
    .A3(net825),
    .S0(net927),
    .S1(net573),
    .X(net945));
 sky130_fd_sc_hd__mux4_1 c262 (.A0(net790),
    .A1(net12),
    .A2(net944),
    .A3(net892),
    .S0(net927),
    .S1(net822),
    .X(net881));
 sky130_fd_sc_hd__mux4_1 c263 (.A0(net6),
    .A1(net941),
    .A2(net8),
    .A3(net807),
    .S0(clknet_1_0__leaf_net916),
    .S1(net927),
    .X(net123));
 sky130_fd_sc_hd__a2111o_4 c264 (.A1(net793),
    .A2(net24),
    .B1(net1016),
    .C1(net19),
    .D1(net1002),
    .X(net124));
 sky130_fd_sc_hd__a2111o_1 c265 (.A1(net124),
    .A2(net26),
    .B1(net1084),
    .C1(net1001),
    .D1(net972),
    .X(net125));
 sky130_fd_sc_hd__mux4_2 c266 (.A0(net1029),
    .A1(net771),
    .A2(net1084),
    .A3(net20),
    .S0(net26),
    .S1(net965),
    .X(net126));
 sky130_fd_sc_hd__a2111o_4 c267 (.A1(net771),
    .A2(net1024),
    .B1(net1002),
    .C1(net965),
    .D1(net978),
    .X(net127));
 sky130_fd_sc_hd__a2111o_4 c268 (.A1(net1057),
    .A2(net1024),
    .B1(net124),
    .C1(net969),
    .D1(net964),
    .X(net128));
 sky130_fd_sc_hd__a2111o_4 c269 (.A1(net128),
    .A2(net1085),
    .B1(net36),
    .C1(net124),
    .D1(net25),
    .X(net129));
 sky130_fd_sc_hd__a2111o_1 c270 (.A1(net771),
    .A2(net129),
    .B1(net974),
    .C1(net965),
    .D1(net1029),
    .X(net130));
 sky130_fd_sc_hd__mux4_1 c271 (.A0(net837),
    .A1(net128),
    .A2(net960),
    .A3(net1050),
    .S0(net772),
    .S1(net1024),
    .X(net131));
 sky130_fd_sc_hd__sdfbbn_2 c272 (.CLK_N(clknet_4_13_0_clk),
    .D(net36),
    .RESET_B(net126),
    .SCD(net960),
    .SCE(net949),
    .SET_B(net980),
    .Q(net133),
    .Q_N(net132));
 sky130_fd_sc_hd__sdfbbp_1 c273 (.CLK(clknet_4_7_0_clk),
    .D(net1050),
    .RESET_B(net133),
    .SCD(net128),
    .SCE(net969),
    .SET_B(net949),
    .Q(net135),
    .Q_N(net134));
 sky130_fd_sc_hd__sdfbbn_2 c274 (.CLK_N(clknet_4_7_0_clk),
    .D(net129),
    .RESET_B(net1026),
    .SCD(net1050),
    .SCE(net960),
    .SET_B(net949),
    .Q(net137),
    .Q_N(net136));
 sky130_fd_sc_hd__mux4_2 c275 (.A0(net964),
    .A1(net20),
    .A2(net136),
    .A3(net969),
    .S0(net1085),
    .S1(net965),
    .X(net138));
 sky130_fd_sc_hd__mux4_1 c276 (.A0(net137),
    .A1(net960),
    .A2(net133),
    .A3(net949),
    .S0(net138),
    .S1(net128),
    .X(net139));
 sky130_fd_sc_hd__mux4_1 c277 (.A0(net1085),
    .A1(net20),
    .A2(net1081),
    .A3(net949),
    .S0(net124),
    .S1(net684),
    .X(net140));
 sky130_fd_sc_hd__mux4_1 c278 (.A0(net804),
    .A1(net138),
    .A2(net960),
    .A3(net949),
    .S0(net1063),
    .S1(net1074),
    .X(net141));
 sky130_fd_sc_hd__mux4_1 c279 (.A0(net949),
    .A1(net137),
    .A2(net965),
    .A3(net960),
    .S0(net576),
    .S1(net684),
    .X(net142));
 sky130_fd_sc_hd__mux4_2 c280 (.A0(net138),
    .A1(net32),
    .A2(net134),
    .A3(net132),
    .S0(net1081),
    .S1(net136),
    .X(net143));
 sky130_fd_sc_hd__mux4_2 c281 (.A0(net1085),
    .A1(net962),
    .A2(net837),
    .A3(net575),
    .S0(net684),
    .S1(net685),
    .X(net144));
 sky130_fd_sc_hd__mux4_1 c282 (.A0(net133),
    .A1(net962),
    .A2(net134),
    .A3(net144),
    .S0(net949),
    .S1(net575),
    .X(net145));
 sky130_fd_sc_hd__mux4_1 c283 (.A0(net144),
    .A1(net962),
    .A2(net950),
    .A3(net576),
    .S0(net685),
    .S1(net687),
    .X(net146));
 sky130_fd_sc_hd__mux4_1 c284 (.A0(net962),
    .A1(net949),
    .A2(net1029),
    .A3(net685),
    .S0(net687),
    .S1(net996),
    .X(net147));
 sky130_fd_sc_hd__a2111o_2 c285 (.A1(net144),
    .A2(net1012),
    .B1(net576),
    .C1(net620),
    .D1(net996),
    .X(net148));
 sky130_fd_sc_hd__mux4_1 c286 (.A0(net972),
    .A1(net897),
    .A2(net1018),
    .A3(net795),
    .S0(net126),
    .S1(net1012),
    .X(net149));
 sky130_fd_sc_hd__mux4_2 c287 (.A0(net42),
    .A1(net793),
    .A2(net798),
    .A3(net576),
    .S0(net668),
    .S1(net994),
    .X(net150));
 sky130_fd_sc_hd__mux4_1 c288 (.A0(net801),
    .A1(net953),
    .A2(net38),
    .A3(net950),
    .S0(net684),
    .S1(net994),
    .X(net151));
 sky130_fd_sc_hd__mux4_1 c289 (.A0(net144),
    .A1(net785),
    .A2(net956),
    .A3(net909),
    .S0(net684),
    .S1(net994),
    .X(net152));
 sky130_fd_sc_hd__mux4_1 c290 (.A0(net1027),
    .A1(net793),
    .A2(net1050),
    .A3(net1024),
    .S0(net955),
    .S1(net994),
    .X(net153));
 sky130_fd_sc_hd__mux4_2 c291 (.A0(net772),
    .A1(net799),
    .A2(net150),
    .A3(net975),
    .S0(net798),
    .S1(net993),
    .X(net154));
 sky130_fd_sc_hd__mux4_2 c292 (.A0(net38),
    .A1(net982),
    .A2(net960),
    .A3(net36),
    .S0(net994),
    .S1(net993),
    .X(net155));
 sky130_fd_sc_hd__mux4_1 c293 (.A0(net950),
    .A1(net771),
    .A2(net785),
    .A3(net909),
    .S0(net623),
    .S1(net994),
    .X(net156));
 sky130_fd_sc_hd__mux4_1 c294 (.A0(net150),
    .A1(net771),
    .A2(net1027),
    .A3(net982),
    .S0(net692),
    .S1(clknet_1_0__leaf_net693),
    .X(net157));
 sky130_fd_sc_hd__mux4_1 c295 (.A0(net977),
    .A1(net962),
    .A2(net144),
    .A3(net1022),
    .S0(clknet_1_0__leaf_net157),
    .S1(net686),
    .X(net900));
 sky130_fd_sc_hd__mux4_1 c296 (.A0(clknet_1_1__leaf_net900),
    .A1(net1021),
    .A2(net155),
    .A3(net994),
    .S0(net993),
    .S1(clknet_1_0__leaf_net693),
    .X(net158));
 sky130_fd_sc_hd__mux4_1 c297 (.A0(net155),
    .A1(net974),
    .A2(net154),
    .A3(net670),
    .S0(net994),
    .S1(clknet_1_0__leaf_net693),
    .X(net159));
 sky130_fd_sc_hd__mux4_1 c298 (.A0(net155),
    .A1(clknet_1_1__leaf_net900),
    .A2(net619),
    .A3(net686),
    .S0(clknet_1_0__leaf_net693),
    .S1(clknet_1_0__leaf_net694),
    .X(net160));
 sky130_fd_sc_hd__mux4_1 c299 (.A0(net575),
    .A1(net619),
    .A2(net687),
    .A3(clknet_1_0__leaf_net693),
    .S0(clknet_1_0__leaf_net694),
    .S1(clknet_1_0__leaf_net695),
    .X(net161));
 sky130_fd_sc_hd__mux4_1 c300 (.A0(clknet_1_1__leaf_net161),
    .A1(clknet_1_1__leaf_net900),
    .A2(net957),
    .A3(clknet_1_0__leaf_net693),
    .S0(clknet_1_0__leaf_net694),
    .S1(clknet_1_0__leaf_net695),
    .X(net162));
 sky130_fd_sc_hd__mux4_1 c301 (.A0(net28),
    .A1(net994),
    .A2(net993),
    .A3(clknet_1_0__leaf_net693),
    .S0(clknet_1_0__leaf_net694),
    .S1(net697),
    .X(net935));
 sky130_fd_sc_hd__mux4_1 c302 (.A0(net793),
    .A1(clknet_1_1__leaf_net900),
    .A2(clknet_1_0__leaf_net935),
    .A3(net150),
    .S0(clknet_1_0__leaf_net161),
    .S1(clknet_1_0__leaf_net694),
    .X(net163));
 sky130_fd_sc_hd__mux4_1 c303 (.A0(net1022),
    .A1(net985),
    .A2(clknet_1_1__leaf_net900),
    .A3(net626),
    .S0(net995),
    .S1(net698),
    .X(net164));
 sky130_fd_sc_hd__mux4_1 c304 (.A0(clknet_1_0__leaf_net161),
    .A1(net969),
    .A2(net953),
    .A3(net1019),
    .S0(net585),
    .S1(net698),
    .X(net165));
 sky130_fd_sc_hd__mux4_1 c305 (.A0(clknet_1_0__leaf_net935),
    .A1(clknet_1_0__leaf_net161),
    .A2(net1021),
    .A3(net785),
    .S0(clknet_1_0__leaf_net693),
    .S1(net697),
    .X(net166));
 sky130_fd_sc_hd__mux4_1 c306 (.A0(net138),
    .A1(clknet_1_1__leaf_net166),
    .A2(net692),
    .A3(clknet_1_0__leaf_net693),
    .S0(clknet_1_0__leaf_net695),
    .S1(net873),
    .X(net167));
 sky130_fd_sc_hd__mux4_1 c307 (.A0(clknet_1_1__leaf_net167),
    .A1(net787),
    .A2(net620),
    .A3(net626),
    .S0(net993),
    .S1(net873),
    .X(net168));
 sky130_fd_sc_hd__mux4_1 c308 (.A0(net785),
    .A1(net42),
    .A2(net830),
    .A3(net809),
    .S0(net155),
    .S1(net968),
    .X(net169));
 sky130_fd_sc_hd__mux4_1 c309 (.A0(net135),
    .A1(clknet_1_1__leaf_net75),
    .A2(net148),
    .A3(net1049),
    .S0(net129),
    .S1(net1019),
    .X(net170));
 sky130_fd_sc_hd__mux4_1 c310 (.A0(net997),
    .A1(net129),
    .A2(clknet_1_1__leaf_net76),
    .A3(clknet_1_1__leaf_net900),
    .S0(net1004),
    .S1(net42),
    .X(net171));
 sky130_fd_sc_hd__mux4_1 c311 (.A0(net954),
    .A1(net1063),
    .A2(net134),
    .A3(net994),
    .S0(net696),
    .S1(net701),
    .X(net172));
 sky130_fd_sc_hd__mux4_2 c312 (.A0(net825),
    .A1(net49),
    .A2(net985),
    .A3(net982),
    .S0(net42),
    .S1(net977),
    .X(net173));
 sky130_fd_sc_hd__mux4_1 c313 (.A0(clknet_1_1__leaf_net66),
    .A1(net173),
    .A2(net1021),
    .A3(net995),
    .S0(net701),
    .S1(net991),
    .X(net174));
 sky130_fd_sc_hd__mux4_2 c314 (.A0(clknet_1_1__leaf_net77),
    .A1(net44),
    .A2(net138),
    .A3(net796),
    .S0(net1015),
    .S1(net991),
    .X(net175));
 sky130_fd_sc_hd__mux4_1 c315 (.A0(net1060),
    .A1(net787),
    .A2(clknet_1_0__leaf_net175),
    .A3(clknet_1_0__leaf_net79),
    .S0(clknet_1_0__leaf_net900),
    .S1(net701),
    .X(net176));
 sky130_fd_sc_hd__mux4_1 c316 (.A0(clknet_1_0__leaf_net166),
    .A1(net952),
    .A2(net827),
    .A3(net830),
    .S0(net701),
    .S1(net703),
    .X(net177));
 sky130_fd_sc_hd__mux4_1 c317 (.A0(clknet_1_1__leaf_net166),
    .A1(net154),
    .A2(net964),
    .A3(net1021),
    .S0(net901),
    .S1(net703),
    .X(net178));
 sky130_fd_sc_hd__mux4_1 c318 (.A0(net967),
    .A1(net1006),
    .A2(clknet_1_0__leaf_net178),
    .A3(clknet_1_1__leaf_net613),
    .S0(net701),
    .S1(net703),
    .X(net179));
 sky130_fd_sc_hd__mux4_1 c319 (.A0(clknet_1_0__leaf_net174),
    .A1(clknet_1_1__leaf_net76),
    .A2(net952),
    .A3(clknet_1_1__leaf_net613),
    .S0(clknet_1_0__leaf_net694),
    .S1(net991),
    .X(net180));
 sky130_fd_sc_hd__mux4_1 c320 (.A0(clknet_1_0__leaf_net178),
    .A1(net897),
    .A2(net771),
    .A3(net982),
    .S0(net991),
    .S1(net703),
    .X(net181));
 sky130_fd_sc_hd__mux4_1 c321 (.A0(clknet_1_1__leaf_net76),
    .A1(clknet_1_1__leaf_net174),
    .A2(net798),
    .A3(net978),
    .S0(net567),
    .S1(net696),
    .X(net182));
 sky130_fd_sc_hd__mux4_1 c322 (.A0(net49),
    .A1(net795),
    .A2(net148),
    .A3(net909),
    .S0(net647),
    .S1(net991),
    .X(net183));
 sky130_fd_sc_hd__mux4_2 c323 (.A0(net971),
    .A1(clknet_1_1__leaf_net77),
    .A2(net173),
    .A3(net822),
    .S0(net991),
    .S1(net703),
    .X(net184));
 sky130_fd_sc_hd__mux4_1 c324 (.A0(net138),
    .A1(net958),
    .A2(clknet_1_0__leaf_net184),
    .A3(net1029),
    .S0(net701),
    .S1(net703),
    .X(net185));
 sky130_fd_sc_hd__mux4_2 c325 (.A0(clknet_1_0__leaf_net182),
    .A1(net71),
    .A2(clknet_1_0__leaf_net184),
    .A3(net1014),
    .S0(net670),
    .S1(net873),
    .X(net186));
 sky130_fd_sc_hd__mux4_1 c326 (.A0(clknet_1_0__leaf_net174),
    .A1(net982),
    .A2(clknet_1_1__leaf_net186),
    .A3(clknet_1_0__leaf_net182),
    .S0(net647),
    .S1(net883),
    .X(net187));
 sky130_fd_sc_hd__mux4_1 c327 (.A0(clknet_1_0__leaf_net186),
    .A1(net967),
    .A2(net568),
    .S0(net647),
    .S1(clknet_1_0__leaf_net673),
    .X(net188));
 sky130_fd_sc_hd__mux4_2 c328 (.A0(clknet_1_0__leaf_net178),
    .A1(clknet_1_0__leaf_net184),
    .A2(net623),
    .A3(net647),
    .S0(net873),
    .S1(net704),
    .X(net922));
 sky130_fd_sc_hd__mux4_1 c329 (.A0(clknet_1_0__leaf_net186),
    .A1(clknet_1_0__leaf_net167),
    .A2(clknet_1_1__leaf_net182),
    .A3(clknet_1_1__leaf_net922),
    .S0(net568),
    .S1(net704),
    .X(net189));
 sky130_fd_sc_hd__mux4_1 c330 (.A0(net855),
    .A1(clknet_1_1__leaf_net179),
    .A2(net86),
    .A3(net830),
    .S0(net1028),
    .S1(net991),
    .X(net190));
 sky130_fd_sc_hd__mux4_1 c331 (.A0(clknet_1_0__leaf_net167),
    .A1(net837),
    .A2(net806),
    .A3(clknet_1_0__leaf_net675),
    .S0(net701),
    .S1(net991),
    .X(net191));
 sky130_fd_sc_hd__mux4_2 c332 (.A0(net856),
    .A1(net830),
    .A2(net798),
    .A3(net805),
    .S0(net698),
    .S1(net704),
    .X(net192));
 sky130_fd_sc_hd__mux4_1 c333 (.A0(net771),
    .A1(clknet_1_0__leaf_net100),
    .A2(net997),
    .A3(net825),
    .S0(net697),
    .S1(net991),
    .X(net193));
 sky130_fd_sc_hd__mux4_1 c334 (.A0(net1080),
    .A1(clknet_1_0__leaf_net175),
    .A2(net801),
    .A3(clknet_1_0__leaf_net79),
    .S0(net138),
    .S1(clknet_1_0__leaf_net193),
    .X(net194));
 sky130_fd_sc_hd__mux4_1 c335 (.A0(net798),
    .A1(net1018),
    .A2(net948),
    .A3(net909),
    .S0(net644),
    .S1(net696),
    .X(net195));
 sky130_fd_sc_hd__mux4_1 c336 (.A0(net85),
    .A1(net1014),
    .A2(net896),
    .A3(net86),
    .S0(net954),
    .S1(clknet_1_0__leaf_net613),
    .X(net196));
 sky130_fd_sc_hd__mux4_1 c337 (.A0(net961),
    .A1(net801),
    .A2(net1019),
    .A3(net948),
    .S0(net796),
    .S1(net704),
    .X(net197));
 sky130_fd_sc_hd__mux4_2 c338 (.A0(net817),
    .A1(net797),
    .A2(net809),
    .A3(net856),
    .S0(net607),
    .S1(net700),
    .X(net198));
 sky130_fd_sc_hd__mux4_1 c339 (.A0(net138),
    .A1(net1018),
    .A2(net841),
    .A3(net909),
    .S0(clknet_1_0__leaf_net674),
    .S1(net706),
    .X(net199));
 sky130_fd_sc_hd__mux4_1 c340 (.A0(clknet_1_0__leaf_net193),
    .A1(net934),
    .A2(net804),
    .A3(net968),
    .S0(net948),
    .S1(net920),
    .X(net200));
 sky130_fd_sc_hd__mux4_1 c341 (.A0(net830),
    .A1(clknet_1_1__leaf_net916),
    .A2(net192),
    .A3(net1083),
    .S0(clknet_1_0__leaf_net179),
    .S1(net678),
    .X(net201));
 sky130_fd_sc_hd__mux4_1 c342 (.A0(net85),
    .A1(net81),
    .A2(clknet_1_1__leaf_net72),
    .A3(net198),
    .S0(net920),
    .S1(net678),
    .X(net202));
 sky130_fd_sc_hd__mux4_1 c343 (.A0(net837),
    .A1(net934),
    .A2(net1049),
    .A3(clknet_1_0__leaf_net202),
    .S0(clknet_1_1__leaf_net922),
    .S1(net86),
    .X(net203));
 sky130_fd_sc_hd__mux4_1 c344 (.A0(clknet_1_0__leaf_net179),
    .A1(net173),
    .A2(clknet_1_1__leaf_net72),
    .A3(clknet_1_0__leaf_net922),
    .S0(net920),
    .S1(net709),
    .X(net204));
 sky130_fd_sc_hd__mux4_1 c345 (.A0(net155),
    .A1(clknet_1_0__leaf_net98),
    .A2(net919),
    .A3(net701),
    .S0(net708),
    .S1(net989),
    .X(net205));
 sky130_fd_sc_hd__mux4_2 c346 (.A0(net830),
    .A1(net198),
    .A2(net644),
    .A3(net990),
    .S0(net709),
    .S1(net989),
    .X(net206));
 sky130_fd_sc_hd__mux4_2 c347 (.A0(net198),
    .A1(net86),
    .A2(net928),
    .A3(net671),
    .S0(net989),
    .S1(net710),
    .X(net207));
 sky130_fd_sc_hd__mux4_1 c348 (.A0(clknet_1_1__leaf_net202),
    .A1(net206),
    .A2(net198),
    .A3(net919),
    .S0(net708),
    .S1(net989),
    .X(net208));
 sky130_fd_sc_hd__mux4_1 c349 (.A0(net797),
    .A1(net855),
    .A2(net896),
    .A3(net709),
    .S0(net921),
    .S1(net710),
    .X(net209));
 sky130_fd_sc_hd__mux4_1 c350 (.A0(net954),
    .A1(net207),
    .A2(net912),
    .A3(net676),
    .S0(net707),
    .S1(net1077),
    .X(net210));
 sky130_fd_sc_hd__mux4_1 c351 (.A0(net838),
    .A1(clknet_1_0__leaf_net75),
    .A2(net87),
    .A3(clknet_1_1__leaf_net179),
    .S1(net710),
    .X(net211));
 sky130_fd_sc_hd__mux4_1 c352 (.A0(net948),
    .A1(net785),
    .A2(net860),
    .A3(net2),
    .S0(clknet_1_0__leaf_net613),
    .S1(net989),
    .X(net212));
 sky130_fd_sc_hd__mux4_1 c353 (.A0(clknet_1_0__leaf_net79),
    .A1(net97),
    .A2(net2),
    .A3(net838),
    .S0(net607),
    .S1(net678),
    .X(net213));
 sky130_fd_sc_hd__mux4_1 c354 (.A0(net118),
    .A1(net999),
    .A2(net840),
    .A3(net97),
    .S0(net607),
    .S1(net989),
    .X(net214));
 sky130_fd_sc_hd__mux4_1 c355 (.A0(net801),
    .A1(clknet_1_0__leaf_net900),
    .A2(net192),
    .A3(net931),
    .S0(net703),
    .S1(net708),
    .X(net215));
 sky130_fd_sc_hd__mux4_1 c356 (.A0(net838),
    .A1(net980),
    .A2(clknet_1_1__leaf_net84),
    .A3(net623),
    .S0(net683),
    .S1(net709),
    .X(net216));
 sky130_fd_sc_hd__mux4_1 c357 (.A0(net0),
    .A1(clknet_1_0__leaf_net936),
    .A2(net971),
    .A3(net804),
    .S0(net703),
    .S1(net989),
    .X(net217));
 sky130_fd_sc_hd__mux4_1 c358 (.A0(net7),
    .A1(net838),
    .A2(net2),
    .A3(net1030),
    .S0(clknet_1_0__leaf_net613),
    .S1(net711),
    .X(net218));
 sky130_fd_sc_hd__mux4_1 c359 (.A0(clknet_1_0__leaf_net218),
    .A1(net868),
    .A2(net484),
    .A3(net869),
    .S0(net909),
    .S1(net708),
    .X(net219));
 sky130_fd_sc_hd__mux4_1 c360 (.A0(net860),
    .A1(net828),
    .A2(clknet_1_0__leaf_net900),
    .A3(net909),
    .S0(net989),
    .S1(net711),
    .X(net220));
 sky130_fd_sc_hd__mux4_1 c361 (.A0(clknet_1_0__leaf_net104),
    .A1(net861),
    .A2(net924),
    .A3(net931),
    .S0(net704),
    .S1(net989),
    .X(net221));
 sky130_fd_sc_hd__mux4_1 c362 (.A0(net7),
    .A1(net817),
    .A2(net999),
    .A3(net806),
    .S0(net833),
    .S1(net934),
    .X(net222));
 sky130_fd_sc_hd__mux4_1 c363 (.A0(net2),
    .A1(clknet_1_1__leaf_net221),
    .A2(net828),
    .A3(net1059),
    .S0(net928),
    .S1(net683),
    .X(net223));
 sky130_fd_sc_hd__mux4_1 c364 (.A0(net97),
    .A1(clknet_1_0__leaf_net104),
    .A2(net917),
    .A3(net214),
    .S0(clknet_1_1__leaf_net693),
    .S1(net703),
    .X(net895));
 sky130_fd_sc_hd__mux4_1 c365 (.A0(net867),
    .A1(clknet_1_1__leaf_net104),
    .A2(clknet_1_1__leaf_net221),
    .A3(clknet_1_0__leaf_net895),
    .S0(net644),
    .S1(net662),
    .X(net224));
 sky130_fd_sc_hd__mux4_1 c366 (.A0(net222),
    .A1(clknet_1_0__leaf_net895),
    .A2(clknet_1_0__leaf_net936),
    .A3(net915),
    .S0(net709),
    .S1(net711),
    .X(net225));
 sky130_fd_sc_hd__mux4_1 c367 (.A0(net173),
    .A1(clknet_1_1__leaf_net218),
    .A2(clknet_1_1__leaf_net116),
    .A3(net833),
    .S0(clknet_1_0__leaf_net895),
    .S1(net711),
    .X(net226));
 sky130_fd_sc_hd__mux4_1 c368 (.A0(clknet_1_0__leaf_net221),
    .A1(clknet_1_1__leaf_net104),
    .A2(net825),
    .A3(net611),
    .S0(net662),
    .S1(net676),
    .X(net227));
 sky130_fd_sc_hd__a2111o_1 c369 (.A1(net917),
    .A2(clknet_1_0__leaf_net221),
    .B1(net837),
    .C1(net633),
    .D1(net662),
    .X(net228));
 sky130_fd_sc_hd__mux4_1 c370 (.A0(net214),
    .A1(net918),
    .A2(net1054),
    .A3(net2),
    .S0(clknet_1_0__leaf_net895),
    .S1(clknet_1_0__leaf_net83),
    .X(net229));
 sky130_fd_sc_hd__mux4_1 c371 (.A0(clknet_1_0__leaf_net75),
    .A1(clknet_1_0__leaf_net199),
    .A2(net2),
    .A3(clknet_1_0__leaf_net895),
    .S0(net611),
    .S1(net919),
    .X(net230));
 sky130_fd_sc_hd__mux4_1 c372 (.A0(clknet_1_1__leaf_net104),
    .A1(net0),
    .A2(net611),
    .A3(net648),
    .S0(net919),
    .S1(net915),
    .X(net231));
 sky130_fd_sc_hd__mux4_1 c373 (.A0(clknet_1_0__leaf_net219),
    .A1(clknet_1_0__leaf_net221),
    .A2(net97),
    .A3(net611),
    .S0(net633),
    .S1(net919),
    .X(net232));
 sky130_fd_sc_hd__a2111o_4 c396 (.A1(net32),
    .A2(net1028),
    .B1(net977),
    .C1(net985),
    .D1(net1003),
    .X(net233));
 sky130_fd_sc_hd__a2111o_2 c397 (.A1(net135),
    .A2(net129),
    .B1(net1024),
    .C1(net977),
    .D1(net686),
    .X(net234));
 sky130_fd_sc_hd__sdfbbn_2 c398 (.CLK_N(clknet_4_12_0_clk),
    .D(net233),
    .RESET_B(net950),
    .SCD(net780),
    .SCE(net1042),
    .SET_B(net686),
    .Q(net236),
    .Q_N(net235));
 sky130_fd_sc_hd__a2111o_2 c399 (.A1(net780),
    .A2(net959),
    .B1(net960),
    .C1(net1085),
    .D1(net686),
    .X(net237));
 sky130_fd_sc_hd__sdfbbp_1 c400 (.CLK(clknet_4_13_0_clk),
    .D(net236),
    .RESET_B(net26),
    .SCD(net1024),
    .SCE(net237),
    .SET_B(net1075),
    .Q(net239),
    .Q_N(net238));
 sky130_fd_sc_hd__a2111o_2 c401 (.A1(net982),
    .A2(net36),
    .B1(net1027),
    .C1(net1085),
    .D1(net132),
    .X(net240));
 sky130_fd_sc_hd__sdfbbn_1 c402 (.CLK_N(clknet_4_7_0_clk),
    .D(net1044),
    .RESET_B(net25),
    .SCD(net1003),
    .SCE(net950),
    .SET_B(net620),
    .Q(net242),
    .Q_N(net241));
 sky130_fd_sc_hd__a2111o_2 c403 (.A1(net242),
    .A2(net1063),
    .B1(net132),
    .C1(net960),
    .D1(net1003),
    .X(net243));
 sky130_fd_sc_hd__mux4_1 c404 (.A0(net35),
    .A1(net1083),
    .A2(net241),
    .A3(net243),
    .S0(net1084),
    .S1(net27),
    .X(net244));
 sky130_fd_sc_hd__sdfbbn_2 c405 (.CLK_N(clknet_4_13_0_clk),
    .D(net19),
    .RESET_B(net243),
    .SCD(net238),
    .SCE(net1010),
    .SET_B(net951),
    .Q(net246),
    .Q_N(net245));
 sky130_fd_sc_hd__a2111o_1 c406 (.A1(net1050),
    .A2(net959),
    .B1(net245),
    .C1(net240),
    .D1(clknet_1_0__leaf_net712),
    .X(net247));
 sky130_fd_sc_hd__a2111o_1 c407 (.A1(net1084),
    .A2(net242),
    .B1(net243),
    .C1(net949),
    .D1(clknet_1_0__leaf_net712),
    .X(net248));
 sky130_fd_sc_hd__mux4_1 c408 (.A0(net246),
    .A1(net243),
    .A2(net126),
    .A3(net124),
    .S0(net588),
    .S1(clknet_1_0__leaf_net712),
    .X(net249));
 sky130_fd_sc_hd__sdfbbp_1 c409 (.CLK(clknet_4_13_0_clk),
    .D(net246),
    .RESET_B(net959),
    .SCD(clknet_1_0__leaf_net247),
    .SCE(net588),
    .SET_B(net1069),
    .Q(net251),
    .Q_N(net250));
 sky130_fd_sc_hd__sdfbbn_1 c410 (.CLK_N(clknet_4_13_0_clk),
    .D(net36),
    .RESET_B(net241),
    .SCD(net243),
    .SCE(clknet_1_0__leaf_net712),
    .SET_B(clknet_1_1__leaf_net713),
    .Q(net253),
    .Q_N(net252));
 sky130_fd_sc_hd__sdfbbn_2 c411 (.CLK_N(clknet_4_13_0_clk),
    .D(net1076),
    .RESET_B(net951),
    .SCD(net245),
    .SCE(net1051),
    .SET_B(clknet_1_1__leaf_net713),
    .Q(net255),
    .Q_N(net254));
 sky130_fd_sc_hd__mux4_1 c412 (.A0(net1085),
    .A1(net242),
    .A2(net246),
    .A3(net133),
    .S0(net240),
    .S1(net243),
    .X(net256));
 sky130_fd_sc_hd__sdfbbp_1 c413 (.CLK(clknet_4_13_0_clk),
    .D(net255),
    .RESET_B(net243),
    .SCD(net960),
    .SCE(net589),
    .SET_B(clknet_1_0__leaf_net712),
    .Q(net258),
    .Q_N(net257));
 sky130_fd_sc_hd__mux4_1 c414 (.A0(net236),
    .A1(net239),
    .A2(net257),
    .A3(net252),
    .S0(clknet_1_1__leaf_net713),
    .S1(clknet_1_0__leaf_net714),
    .X(net893));
 sky130_fd_sc_hd__mux4_1 c415 (.A0(net251),
    .A1(net240),
    .A2(net948),
    .A3(net588),
    .S0(clknet_1_0__leaf_net712),
    .S1(clknet_1_0__leaf_net714),
    .X(net259));
 sky130_fd_sc_hd__mux4_1 c416 (.A0(net26),
    .A1(net253),
    .A2(net257),
    .A3(net959),
    .S0(net233),
    .S1(clknet_1_0__leaf_net714),
    .X(net260));
 sky130_fd_sc_hd__mux4_1 c417 (.A0(clknet_1_1__leaf_net260),
    .A1(clknet_1_1__leaf_net893),
    .A2(net245),
    .A3(net233),
    .S0(clknet_1_0__leaf_net714),
    .S1(net716),
    .X(net261));
 sky130_fd_sc_hd__mux4_1 c418 (.A0(net126),
    .A1(net258),
    .A2(net977),
    .A3(net957),
    .S0(clknet_1_1__leaf_net695),
    .S1(clknet_1_1__leaf_net713),
    .X(net262));
 sky130_fd_sc_hd__mux4_1 c419 (.A0(clknet_1_1__leaf_net161),
    .A1(net1003),
    .A2(net235),
    .A3(net964),
    .S0(net1022),
    .S1(net716),
    .X(net263));
 sky130_fd_sc_hd__mux4_1 c420 (.A0(clknet_1_1__leaf_net161),
    .A1(clknet_1_1__leaf_net166),
    .A2(net954),
    .A3(net1049),
    .S0(net985),
    .S1(net698),
    .X(net264));
 sky130_fd_sc_hd__mux4_1 c421 (.A0(clknet_1_1__leaf_net263),
    .A1(clknet_1_0__leaf_net168),
    .A2(net148),
    .A3(net589),
    .S0(net619),
    .S1(net717),
    .X(net265));
 sky130_fd_sc_hd__mux4_1 c422 (.A0(net1007),
    .A1(clknet_1_0__leaf_net260),
    .A2(net604),
    .A3(net688),
    .S0(clknet_1_0__leaf_net712),
    .S1(net719),
    .X(net266));
 sky130_fd_sc_hd__mux4_1 c423 (.A0(net1026),
    .A1(clknet_1_0__leaf_net168),
    .A2(net805),
    .A3(net148),
    .S0(net620),
    .S1(net720),
    .X(net267));
 sky130_fd_sc_hd__mux4_1 c424 (.A0(net49),
    .A1(net954),
    .A2(net1022),
    .A3(net686),
    .S0(net719),
    .S1(net988),
    .X(net268));
 sky130_fd_sc_hd__mux4_2 c425 (.A0(net26),
    .A1(net258),
    .A2(net970),
    .A3(net589),
    .S0(net604),
    .S1(net715),
    .X(net269));
 sky130_fd_sc_hd__mux4_1 c426 (.A0(net258),
    .A1(clknet_1_1__leaf_net166),
    .A2(net1018),
    .A3(net953),
    .S0(net48),
    .S1(net909),
    .X(net270));
 sky130_fd_sc_hd__mux4_2 c427 (.A0(net135),
    .A1(net36),
    .A2(net1007),
    .A3(net269),
    .S0(net715),
    .S1(net724),
    .X(net271));
 sky130_fd_sc_hd__mux4_1 c428 (.A0(clknet_1_1__leaf_net260),
    .A1(net269),
    .A2(net1019),
    .A3(net1049),
    .S0(net271),
    .S1(clknet_1_1__leaf_net713),
    .X(net272));
 sky130_fd_sc_hd__mux4_1 c429 (.A0(net129),
    .A1(net240),
    .A2(net269),
    .A3(clknet_1_0__leaf_net712),
    .S0(net723),
    .S1(net725),
    .X(net273));
 sky130_fd_sc_hd__mux4_1 c430 (.A0(net269),
    .A1(clknet_1_0__leaf_net247),
    .A2(clknet_1_1__leaf_net273),
    .A3(clknet_1_0__leaf_net157),
    .S0(net150),
    .S1(net725),
    .X(net274));
 sky130_fd_sc_hd__mux4_1 c431 (.A0(net240),
    .A1(net799),
    .A2(net1044),
    .A3(net954),
    .S0(net721),
    .S1(net727),
    .X(net275));
 sky130_fd_sc_hd__mux4_1 c432 (.A0(clknet_1_1__leaf_net273),
    .A1(net39),
    .A2(net671),
    .A3(clknet_1_1__leaf_net695),
    .S0(net719),
    .S1(net988),
    .X(net276));
 sky130_fd_sc_hd__mux4_1 c433 (.A0(clknet_1_1__leaf_net713),
    .A1(net721),
    .A2(net988),
    .A3(net724),
    .S0(net726),
    .S1(net728),
    .X(net277));
 sky130_fd_sc_hd__mux4_1 c434 (.A0(net40),
    .A1(net806),
    .A2(clknet_1_1__leaf_net263),
    .A3(clknet_1_0__leaf_net277),
    .S0(net974),
    .S1(net726),
    .X(net898));
 sky130_fd_sc_hd__mux4_1 c435 (.A0(clknet_1_1__leaf_net277),
    .A1(clknet_1_0__leaf_net276),
    .A2(net257),
    .A3(net589),
    .S0(net685),
    .S1(net728),
    .X(net278));
 sky130_fd_sc_hd__mux4_1 c436 (.A0(net124),
    .A1(net1063),
    .A2(clknet_1_1__leaf_net898),
    .A3(net717),
    .S0(net720),
    .S1(net729),
    .X(net279));
 sky130_fd_sc_hd__mux4_1 c437 (.A0(clknet_1_0__leaf_net273),
    .A1(net154),
    .A2(clknet_1_1__leaf_net898),
    .A3(net725),
    .S0(net727),
    .S1(net730),
    .X(net280));
 sky130_fd_sc_hd__mux4_1 c438 (.A0(net799),
    .A1(clknet_1_1__leaf_net277),
    .A2(clknet_1_0__leaf_net898),
    .A3(clknet_1_1__leaf_net273),
    .S0(clknet_1_0__leaf_net260),
    .S1(net729),
    .X(net281));
 sky130_fd_sc_hd__a2111o_1 c439 (.A1(net1063),
    .A2(clknet_1_0__leaf_net898),
    .B1(net591),
    .C1(net700),
    .D1(net730),
    .X(net282));
 sky130_fd_sc_hd__mux4_1 c440 (.A0(net68),
    .A1(net962),
    .A2(clknet_1_0__leaf_net166),
    .A3(net1018),
    .S0(net568),
    .S1(net601),
    .X(net283));
 sky130_fd_sc_hd__mux4_1 c441 (.A0(net239),
    .A1(net235),
    .A2(net601),
    .A3(clknet_1_0__leaf_net675),
    .S0(net719),
    .S1(net727),
    .X(net284));
 sky130_fd_sc_hd__mux4_1 c442 (.A0(clknet_1_0__leaf_net74),
    .A1(net968),
    .A2(net1024),
    .A3(net71),
    .S0(net601),
    .S1(net912),
    .X(net285));
 sky130_fd_sc_hd__mux4_1 c443 (.A0(net811),
    .A1(net47),
    .A2(net238),
    .A3(net967),
    .S0(net53),
    .S1(net591),
    .X(net286));
 sky130_fd_sc_hd__mux4_1 c444 (.A0(net1054),
    .A1(net1042),
    .A2(net591),
    .A3(net901),
    .S0(net692),
    .S1(net732),
    .X(net287));
 sky130_fd_sc_hd__mux4_1 c445 (.A0(clknet_1_1__leaf_net184),
    .A1(net287),
    .A2(net1015),
    .A3(net971),
    .S0(net912),
    .S1(net732),
    .X(net288));
 sky130_fd_sc_hd__mux4_1 c446 (.A0(clknet_1_1__leaf_net72),
    .A1(net235),
    .A2(clknet_1_1__leaf_net288),
    .A3(clknet_1_0__leaf_net263),
    .S0(net590),
    .S1(net696),
    .X(net289));
 sky130_fd_sc_hd__mux4_1 c447 (.A0(clknet_1_1__leaf_net288),
    .A1(net952),
    .A2(net49),
    .A3(net795),
    .S0(net647),
    .S1(net732),
    .X(net290));
 sky130_fd_sc_hd__mux4_1 c448 (.A0(clknet_1_1__leaf_net288),
    .A1(net567),
    .A2(net619),
    .A3(net665),
    .S0(net692),
    .S1(net725),
    .X(net291));
 sky130_fd_sc_hd__mux4_1 c449 (.A0(clknet_1_1__leaf_net70),
    .A1(clknet_1_0__leaf_net178),
    .A2(clknet_1_0__leaf_net893),
    .A3(net948),
    .S0(net1028),
    .S1(net720),
    .X(net292));
 sky130_fd_sc_hd__mux4_1 c450 (.A0(net974),
    .A1(net967),
    .A2(clknet_1_0__leaf_net157),
    .A3(net590),
    .S0(net726),
    .S1(net732),
    .X(net293));
 sky130_fd_sc_hd__mux4_1 c451 (.A0(clknet_1_0__leaf_net284),
    .A1(clknet_1_0__leaf_net73),
    .A2(clknet_1_0__leaf_net288),
    .A3(net805),
    .S0(net1003),
    .S1(net721),
    .X(net294));
 sky130_fd_sc_hd__mux4_1 c452 (.A0(net42),
    .A1(clknet_1_1__leaf_net174),
    .A2(net974),
    .A3(clknet_1_1__leaf_net674),
    .S0(clknet_1_0__leaf_net734),
    .S1(clknet_1_0__leaf_net735),
    .X(net904));
 sky130_fd_sc_hd__mux4_1 c453 (.A0(clknet_1_0__leaf_net293),
    .A1(net963),
    .A2(net982),
    .A3(net150),
    .S0(net619),
    .S1(net671),
    .X(net295));
 sky130_fd_sc_hd__mux4_1 c454 (.A0(net797),
    .A1(clknet_1_0__leaf_net283),
    .A2(clknet_1_0__leaf_net904),
    .A3(clknet_1_0__leaf_net713),
    .S0(clknet_1_0__leaf_net733),
    .S1(clknet_1_0__leaf_net735),
    .X(net296));
 sky130_fd_sc_hd__mux4_1 c455 (.A0(clknet_1_0__leaf_net157),
    .A1(clknet_1_0__leaf_net296),
    .A2(clknet_1_0__leaf_net904),
    .A3(clknet_1_0__leaf_net295),
    .S0(net901),
    .S1(net724),
    .X(net297));
 sky130_fd_sc_hd__mux4_1 c456 (.A0(clknet_1_1__leaf_net295),
    .A1(net982),
    .A2(clknet_1_0__leaf_net178),
    .A3(net647),
    .S0(net665),
    .S1(net732),
    .X(net298));
 sky130_fd_sc_hd__mux4_1 c457 (.A0(clknet_1_1__leaf_net296),
    .A1(clknet_1_1__leaf_net295),
    .A2(net811),
    .A3(net645),
    .S0(net911),
    .S1(clknet_1_0__leaf_net733),
    .X(net299));
 sky130_fd_sc_hd__mux4_1 c458 (.A0(clknet_1_1__leaf_net182),
    .A1(clknet_1_1__leaf_net284),
    .A2(clknet_1_1__leaf_net288),
    .A3(clknet_1_0__leaf_net296),
    .S0(net601),
    .S1(net665),
    .X(net300));
 sky130_fd_sc_hd__mux4_1 c459 (.A0(clknet_1_0__leaf_net295),
    .A1(clknet_1_0__leaf_net296),
    .A2(net953),
    .A3(net645),
    .S0(net901),
    .S1(clknet_1_1__leaf_net735),
    .X(net301));
 sky130_fd_sc_hd__mux4_1 c460 (.A0(clknet_1_1__leaf_net283),
    .A1(net974),
    .A2(net645),
    .A3(net732),
    .S0(net736),
    .S1(net889),
    .X(net302));
 sky130_fd_sc_hd__mux4_1 c461 (.A0(net796),
    .A1(clknet_1_1__leaf_net302),
    .A2(clknet_1_0__leaf_net898),
    .A3(net911),
    .S0(net723),
    .S1(net738),
    .X(net303));
 sky130_fd_sc_hd__mux4_1 c462 (.A0(clknet_1_1__leaf_net887),
    .A1(net1001),
    .A2(net646),
    .A3(net665),
    .S0(clknet_1_1__leaf_net674),
    .S1(net739),
    .X(net304));
 sky130_fd_sc_hd__mux4_1 c463 (.A0(clknet_1_0__leaf_net273),
    .A1(net90),
    .A2(net978),
    .A3(net911),
    .S0(net672),
    .S1(clknet_1_1__leaf_net735),
    .X(net908));
 sky130_fd_sc_hd__mux4_2 c464 (.A0(clknet_1_1__leaf_net175),
    .A1(net967),
    .A2(net975),
    .A3(net669),
    .S0(clknet_1_0__leaf_net713),
    .S1(clknet_1_0__leaf_net735),
    .X(net905));
 sky130_fd_sc_hd__mux4_1 c465 (.A0(clknet_1_0__leaf_net302),
    .A1(clknet_1_1__leaf_net78),
    .A2(clknet_1_1__leaf_net908),
    .A3(net604),
    .S0(net928),
    .S1(net992),
    .X(net305));
 sky130_fd_sc_hd__mux4_1 c466 (.A0(net841),
    .A1(net1043),
    .A2(net1080),
    .A3(net928),
    .S0(net995),
    .S1(net741),
    .X(net306));
 sky130_fd_sc_hd__mux4_1 c467 (.A0(net209),
    .A1(net961),
    .A2(net804),
    .A3(net238),
    .S0(net706),
    .S1(clknet_1_1__leaf_net735),
    .X(net307));
 sky130_fd_sc_hd__mux4_1 c468 (.A0(net306),
    .A1(net1080),
    .A2(clknet_1_0__leaf_net285),
    .A3(clknet_1_1__leaf_net887),
    .S0(net321),
    .S1(net1043),
    .X(net308));
 sky130_fd_sc_hd__mux4_1 c469 (.A0(net321),
    .A1(net1082),
    .A2(net81),
    .A3(net705),
    .S0(net723),
    .S1(net731),
    .X(net309));
 sky130_fd_sc_hd__mux4_2 c470 (.A0(clknet_1_0__leaf_net904),
    .A1(clknet_1_1__leaf_net78),
    .A2(net841),
    .A3(net1080),
    .S0(clknet_1_1__leaf_net735),
    .S1(net741),
    .X(net310));
 sky130_fd_sc_hd__mux4_1 c471 (.A0(net827),
    .A1(clknet_1_0__leaf_net288),
    .A2(net977),
    .A3(net822),
    .S0(net309),
    .S1(net570),
    .X(net311));
 sky130_fd_sc_hd__mux4_1 c472 (.A0(net309),
    .A1(clknet_1_0__leaf_net208),
    .A2(clknet_1_0__leaf_net938),
    .A3(clknet_1_1__leaf_net693),
    .S0(clknet_1_0__leaf_net713),
    .S1(net741),
    .X(net894));
 sky130_fd_sc_hd__mux4_1 c473 (.A0(clknet_1_1__leaf_net191),
    .A1(net1018),
    .A2(clknet_1_1__leaf_net100),
    .A3(net250),
    .S0(clknet_1_0__leaf_net208),
    .S1(net81),
    .X(net312));
 sky130_fd_sc_hd__mux4_1 c474 (.A0(clknet_1_0__leaf_net312),
    .A1(net980),
    .A2(clknet_1_0__leaf_net893),
    .A3(net828),
    .S0(net306),
    .S1(clknet_1_0__leaf_net307),
    .X(net313));
 sky130_fd_sc_hd__mux4_1 c475 (.A0(clknet_1_1__leaf_net193),
    .A1(clknet_1_1__leaf_net175),
    .A2(clknet_1_1__leaf_net887),
    .A3(net91),
    .S0(clknet_1_0__leaf_net893),
    .S1(net742),
    .X(net314));
 sky130_fd_sc_hd__mux4_1 c476 (.A0(net980),
    .A1(clknet_1_0__leaf_net887),
    .A2(net604),
    .A3(net609),
    .S0(clknet_1_1__leaf_net938),
    .S1(net742),
    .X(net315));
 sky130_fd_sc_hd__mux4_1 c477 (.A0(net1031),
    .A1(clknet_1_1__leaf_net84),
    .A2(net952),
    .A3(net604),
    .S0(net742),
    .S1(net743),
    .X(net316));
 sky130_fd_sc_hd__mux4_1 c478 (.A0(net978),
    .A1(clknet_1_1__leaf_net312),
    .A2(net1080),
    .A3(net609),
    .S0(net742),
    .S1(net743),
    .X(net317));
 sky130_fd_sc_hd__mux4_1 c479 (.A0(net209),
    .A1(clknet_1_0__leaf_net285),
    .A2(net646),
    .A3(clknet_1_1__leaf_net938),
    .S0(clknet_1_1__leaf_net674),
    .S1(net743),
    .X(net318));
 sky130_fd_sc_hd__mux4_1 c480 (.A0(clknet_1_1__leaf_net208),
    .A1(net1080),
    .A2(clknet_1_0__leaf_net98),
    .A3(clknet_1_0__leaf_net288),
    .S0(net1016),
    .S1(net705),
    .X(net319));
 sky130_fd_sc_hd__mux4_1 c481 (.A0(clknet_1_1__leaf_net193),
    .A1(clknet_1_0__leaf_net904),
    .A2(net836),
    .A3(net604),
    .S0(clknet_1_1__leaf_net674),
    .S1(net723),
    .X(net320));
 sky130_fd_sc_hd__mux4_1 c482 (.A0(net86),
    .A1(net896),
    .A2(net821),
    .A3(net676),
    .S0(net991),
    .S1(net913),
    .X(net321));
 sky130_fd_sc_hd__mux4_1 c483 (.A0(net91),
    .A1(net814),
    .A2(net250),
    .A3(clknet_1_0__leaf_net191),
    .S0(net821),
    .S1(net992),
    .X(net887));
 sky130_fd_sc_hd__mux4_1 c484 (.A0(clknet_1_0__leaf_net219),
    .A1(net251),
    .A2(net861),
    .A3(net833),
    .S0(net648),
    .S1(net743),
    .X(net322));
 sky130_fd_sc_hd__mux4_1 c485 (.A0(clknet_1_0__leaf_net905),
    .A1(net206),
    .A2(clknet_1_1__leaf_net79),
    .A3(net907),
    .S0(net626),
    .S1(net743),
    .X(net323));
 sky130_fd_sc_hd__mux4_1 c486 (.A0(net840),
    .A1(net239),
    .A2(clknet_1_1__leaf_net219),
    .A3(net646),
    .S0(net661),
    .S1(net743),
    .X(net899));
 sky130_fd_sc_hd__mux4_1 c487 (.A0(net322),
    .A1(net858),
    .A2(net948),
    .A3(clknet_1_0__leaf_net675),
    .S0(net724),
    .S1(net744),
    .X(net324));
 sky130_fd_sc_hd__mux4_1 c488 (.A0(net71),
    .A1(net1082),
    .A2(net484),
    .A3(net1015),
    .S0(net672),
    .S1(net990),
    .X(net325));
 sky130_fd_sc_hd__mux4_1 c489 (.A0(net833),
    .A1(clknet_1_0__leaf_net116),
    .A2(net821),
    .A3(net797),
    .S0(net954),
    .S1(net902),
    .X(net326));
 sky130_fd_sc_hd__mux4_1 c490 (.A0(net239),
    .A1(net150),
    .A2(net192),
    .A3(net858),
    .S0(net711),
    .S1(net988),
    .X(net327));
 sky130_fd_sc_hd__mux4_1 c491 (.A0(net868),
    .A1(net822),
    .A2(net1082),
    .A3(net626),
    .S0(net928),
    .S1(clknet_1_1__leaf_net651),
    .X(net328));
 sky130_fd_sc_hd__mux4_2 c492 (.A0(net5),
    .A1(net648),
    .A2(net940),
    .A3(net683),
    .S0(net990),
    .S1(net744),
    .X(net329));
 sky130_fd_sc_hd__mux4_1 c493 (.A0(net327),
    .A1(net71),
    .A2(net329),
    .A3(net948),
    .S0(net907),
    .S1(net901),
    .X(net330));
 sky130_fd_sc_hd__mux4_1 c494 (.A0(clknet_1_1__leaf_net104),
    .A1(net798),
    .A2(net999),
    .A3(net806),
    .S0(net1082),
    .S1(net990),
    .X(net890));
 sky130_fd_sc_hd__mux4_1 c495 (.A0(clknet_1_0__leaf_net263),
    .A1(net329),
    .A2(net971),
    .A3(net901),
    .S0(net940),
    .S1(net744),
    .X(net331));
 sky130_fd_sc_hd__mux4_1 c496 (.A0(clknet_1_0__leaf_net111),
    .A1(clknet_1_1__leaf_net84),
    .A2(clknet_1_1__leaf_net116),
    .A3(net329),
    .S0(clknet_1_1__leaf_net219),
    .S1(net671),
    .X(net332));
 sky130_fd_sc_hd__mux4_1 c497 (.A0(net5),
    .A1(net857),
    .A2(clknet_1_0__leaf_net231),
    .A3(net868),
    .S0(net1028),
    .S1(net720),
    .X(net333));
 sky130_fd_sc_hd__mux4_1 c498 (.A0(net206),
    .A1(net331),
    .A2(clknet_1_1__leaf_net111),
    .A3(net570),
    .S0(net683),
    .S1(net744),
    .X(net334));
 sky130_fd_sc_hd__mux4_1 c499 (.A0(net5),
    .A1(net329),
    .A2(net779),
    .A3(clknet_1_0__leaf_net616),
    .S0(net661),
    .S1(net903),
    .X(net335));
 sky130_fd_sc_hd__mux4_1 c500 (.A0(clknet_1_0__leaf_net328),
    .A1(clknet_1_0__leaf_net890),
    .A2(net329),
    .A3(clknet_1_0__leaf_net713),
    .S0(net724),
    .S1(net913),
    .X(net336));
 sky130_fd_sc_hd__mux4_1 c501 (.A0(clknet_1_0__leaf_net288),
    .A1(clknet_1_1__leaf_net328),
    .A2(clknet_1_0__leaf_net336),
    .A3(net646),
    .S0(net711),
    .S1(net988),
    .X(net337));
 sky130_fd_sc_hd__mux4_1 c502 (.A0(clknet_1_1__leaf_net336),
    .A1(net954),
    .A2(net1028),
    .A3(net90),
    .S0(clknet_1_0__leaf_net333),
    .S1(net805),
    .X(net338));
 sky130_fd_sc_hd__mux4_1 c503 (.A0(net325),
    .A1(clknet_1_1__leaf_net219),
    .A2(net858),
    .A3(net948),
    .S0(net635),
    .S1(net745),
    .X(net339));
 sky130_fd_sc_hd__mux4_1 c504 (.A0(net334),
    .A1(net1001),
    .A2(clknet_1_1__leaf_net890),
    .A3(clknet_1_0__leaf_net900),
    .S0(net901),
    .S1(net746),
    .X(net340));
 sky130_fd_sc_hd__mux4_1 c505 (.A0(net822),
    .A1(net948),
    .A2(net1),
    .A3(clknet_1_0__leaf_net616),
    .S0(net744),
    .S1(net746),
    .X(net341));
 sky130_fd_sc_hd__mux4_1 c528 (.A0(net961),
    .A1(clknet_1_1__leaf_net893),
    .A2(clknet_1_0__leaf_net247),
    .A3(net252),
    .S0(net959),
    .S1(net951),
    .X(net342));
 sky130_fd_sc_hd__sdfbbn_1 c529 (.CLK_N(clknet_4_13_0_clk),
    .D(net775),
    .RESET_B(net1071),
    .SCD(net951),
    .SCE(net35),
    .SET_B(net688),
    .Q(net344),
    .Q_N(net343));
 sky130_fd_sc_hd__a2111o_4 c530 (.A1(net128),
    .A2(net241),
    .B1(net970),
    .C1(net1013),
    .D1(net982),
    .X(net345));
 sky130_fd_sc_hd__a2111o_1 c531 (.A1(net22),
    .A2(net345),
    .B1(net1013),
    .C1(net688),
    .D1(clknet_1_0__leaf_net712),
    .X(net346));
 sky130_fd_sc_hd__sdfbbn_1 c532 (.CLK_N(clknet_4_15_0_clk),
    .D(net959),
    .RESET_B(net237),
    .SCD(net1007),
    .SCE(net986),
    .SET_B(net687),
    .Q(net348),
    .Q_N(net347));
 sky130_fd_sc_hd__sdfbbp_1 c533 (.CLK(clknet_4_13_0_clk),
    .D(net124),
    .RESET_B(net128),
    .SCD(net245),
    .SCE(net951),
    .SET_B(net1068),
    .Q(net350),
    .Q_N(net349));
 sky130_fd_sc_hd__sdfbbn_1 c534 (.CLK_N(clknet_4_13_0_clk),
    .D(net345),
    .RESET_B(net25),
    .SCD(clknet_1_0__leaf_net247),
    .SCE(net343),
    .SET_B(clknet_1_1__leaf_net712),
    .Q(net352),
    .Q_N(net351));
 sky130_fd_sc_hd__a2111o_1 c535 (.A1(clknet_1_1__leaf_net346),
    .A2(net347),
    .B1(net1007),
    .C1(net349),
    .D1(net747),
    .X(net353));
 sky130_fd_sc_hd__a2111o_1 c536 (.A1(net348),
    .A2(net970),
    .B1(clknet_1_1__leaf_net346),
    .C1(net143),
    .D1(net1010),
    .X(net354));
 sky130_fd_sc_hd__a2111o_1 c537 (.A1(net350),
    .A2(clknet_1_1__leaf_net354),
    .B1(net35),
    .C1(net22),
    .D1(net970),
    .X(net355));
 sky130_fd_sc_hd__sdfbbn_1 c538 (.CLK_N(clknet_4_15_0_clk),
    .D(net1072),
    .RESET_B(clknet_1_1__leaf_net353),
    .SCD(clknet_1_1__leaf_net354),
    .SCE(net1051),
    .SET_B(net687),
    .Q(net357),
    .Q_N(net356));
 sky130_fd_sc_hd__a2111o_1 c539 (.A1(net357),
    .A2(net253),
    .B1(net246),
    .C1(net237),
    .D1(clknet_1_1__leaf_net353),
    .X(net358));
 sky130_fd_sc_hd__sdfbbp_1 c540 (.CLK(clknet_4_15_0_clk),
    .D(net352),
    .RESET_B(net357),
    .SCD(clknet_1_1__leaf_net353),
    .SCE(net579),
    .SET_B(net1070),
    .Q(net360),
    .Q_N(net359));
 sky130_fd_sc_hd__sdfbbn_2 c541 (.CLK_N(clknet_4_15_0_clk),
    .D(net1076),
    .RESET_B(net1073),
    .SCD(net349),
    .SCE(clknet_1_1__leaf_net353),
    .SET_B(net579),
    .Q(net362),
    .Q_N(net361));
 sky130_fd_sc_hd__a2111o_1 c542 (.A1(net362),
    .A2(net1064),
    .B1(net360),
    .C1(net1045),
    .D1(net951),
    .X(net363));
 sky130_fd_sc_hd__a2111o_4 c543 (.A1(net360),
    .A2(net972),
    .B1(net361),
    .C1(net1003),
    .D1(net579),
    .X(net364));
 sky130_fd_sc_hd__mux4_1 c544 (.A0(net25),
    .A1(net364),
    .A2(net1041),
    .A3(net237),
    .S0(net361),
    .S1(net618),
    .X(net365));
 sky130_fd_sc_hd__mux4_2 c545 (.A0(net344),
    .A1(net362),
    .A2(net252),
    .A3(net364),
    .S0(net136),
    .S1(net891),
    .X(net366));
 sky130_fd_sc_hd__a2111o_1 c546 (.A1(net237),
    .A2(net126),
    .B1(clknet_1_1__leaf_net346),
    .C1(net364),
    .D1(net361),
    .X(net367));
 sky130_fd_sc_hd__mux4_1 c547 (.A0(net366),
    .A1(net361),
    .A2(net345),
    .A3(net241),
    .S0(net640),
    .S1(net891),
    .X(net368));
 sky130_fd_sc_hd__sdfbbn_1 c548 (.CLK_N(clknet_4_14_0_clk),
    .D(net368),
    .RESET_B(clknet_1_0__leaf_net354),
    .SCD(net364),
    .SCE(net361),
    .SET_B(net891),
    .Q(net370),
    .Q_N(net369));
 sky130_fd_sc_hd__mux4_1 c549 (.A0(net243),
    .A1(net364),
    .A2(net368),
    .A3(net1056),
    .S0(net361),
    .S1(net640),
    .X(net371));
 sky130_fd_sc_hd__sdfbbp_1 c550 (.CLK(clknet_4_12_0_clk),
    .D(clknet_1_1__leaf_net168),
    .RESET_B(net951),
    .SCD(net254),
    .SCE(clknet_1_1__leaf_net935),
    .SET_B(net1075),
    .Q(net874),
    .Q_N(net372));
 sky130_fd_sc_hd__a2111o_1 c551 (.A1(net1022),
    .A2(net233),
    .B1(clknet_1_1__leaf_net277),
    .C1(clknet_1_1__leaf_net157),
    .D1(net271),
    .X(net373));
 sky130_fd_sc_hd__a2111o_1 c552 (.A1(net25),
    .A2(net978),
    .B1(net27),
    .C1(net685),
    .D1(net692),
    .X(net374));
 sky130_fd_sc_hd__a2111o_2 c553 (.A1(net368),
    .A2(net966),
    .B1(net961),
    .C1(net579),
    .D1(net722),
    .X(net375));
 sky130_fd_sc_hd__mux4_1 c554 (.A0(net352),
    .A1(net375),
    .A2(net271),
    .A3(net957),
    .S0(net484),
    .S1(net688),
    .X(net376));
 sky130_fd_sc_hd__mux4_1 c555 (.A0(net374),
    .A1(net1022),
    .A2(clknet_1_1__leaf_net695),
    .A3(net699),
    .S0(net717),
    .S1(net721),
    .X(net377));
 sky130_fd_sc_hd__mux4_1 c556 (.A0(net364),
    .A1(clknet_1_1__leaf_net168),
    .A2(clknet_1_0__leaf_net373),
    .A3(net1018),
    .S0(net808),
    .S1(net692),
    .X(net378));
 sky130_fd_sc_hd__a2111o_1 c557 (.A1(net799),
    .A2(net271),
    .B1(net1024),
    .C1(clknet_1_1__leaf_net273),
    .D1(clknet_1_0__leaf_net377),
    .X(net379));
 sky130_fd_sc_hd__mux4_1 c558 (.A0(clknet_1_1__leaf_net378),
    .A1(net1066),
    .A2(net1041),
    .A3(clknet_1_1__leaf_net157),
    .S0(net953),
    .S1(net749),
    .X(net380));
 sky130_fd_sc_hd__a2111o_1 c559 (.A1(net369),
    .A2(net43),
    .B1(net351),
    .C1(net604),
    .D1(net749),
    .X(net381));
 sky130_fd_sc_hd__sdfbbn_2 c560 (.CLK_N(clknet_4_9_0_clk),
    .D(net966),
    .RESET_B(clknet_1_1__leaf_net277),
    .SCD(net957),
    .SCE(net579),
    .SET_B(net748),
    .Q(net383),
    .Q_N(net382));
 sky130_fd_sc_hd__a2111o_1 c561 (.A1(net381),
    .A2(clknet_1_0__leaf_net276),
    .B1(net236),
    .C1(net668),
    .D1(net697),
    .X(net384));
 sky130_fd_sc_hd__sdfbbn_1 c562 (.CLK_N(clknet_4_12_0_clk),
    .D(clknet_1_0__leaf_net379),
    .RESET_B(net374),
    .SCD(net966),
    .SCE(net569),
    .SET_B(net672),
    .Q(net888),
    .Q_N(net385));
 sky130_fd_sc_hd__a2111o_1 c563 (.A1(clknet_1_0__leaf_net354),
    .A2(net888),
    .B1(net381),
    .C1(net1020),
    .D1(net382),
    .X(net386));
 sky130_fd_sc_hd__mux4_1 c564 (.A0(net385),
    .A1(net964),
    .A2(net382),
    .A3(net604),
    .S0(net730),
    .S1(net749),
    .X(net387));
 sky130_fd_sc_hd__mux4_1 c565 (.A0(net387),
    .A1(clknet_1_1__leaf_net377),
    .A2(net43),
    .A3(net951),
    .S0(net796),
    .S1(net640),
    .X(net388));
 sky130_fd_sc_hd__mux4_1 c566 (.A0(clknet_1_0__leaf_net378),
    .A1(net124),
    .A2(clknet_1_1__leaf_net379),
    .A3(net1094),
    .S0(net381),
    .S1(net749),
    .X(net389));
 sky130_fd_sc_hd__a2111o_1 c567 (.A1(net233),
    .A2(net1027),
    .B1(clknet_1_0__leaf_net377),
    .C1(net569),
    .D1(clknet_1_1__leaf_net615),
    .X(net390));
 sky130_fd_sc_hd__mux4_1 c568 (.A0(net271),
    .A1(clknet_1_0__leaf_net379),
    .A2(net385),
    .A3(net254),
    .S0(clknet_1_1__leaf_net615),
    .S1(net749),
    .X(net391));
 sky130_fd_sc_hd__a2111o_1 c569 (.A1(net383),
    .A2(clknet_1_1__leaf_net615),
    .B1(net996),
    .C1(net995),
    .D1(clknet_1_1__leaf_net751),
    .X(net392));
 sky130_fd_sc_hd__a2111o_1 c570 (.A1(clknet_1_0__leaf_net392),
    .A2(net387),
    .B1(net383),
    .C1(net235),
    .D1(clknet_1_0__leaf_net377),
    .X(net393));
 sky130_fd_sc_hd__mux4_1 c571 (.A0(net393),
    .A1(clknet_1_1__leaf_net390),
    .A2(net374),
    .A3(net1006),
    .S0(net385),
    .S1(clknet_1_0__leaf_net615),
    .X(net939));
 sky130_fd_sc_hd__mux4_1 c572 (.A0(clknet_1_1__leaf_net74),
    .A1(net828),
    .A2(clknet_1_0__leaf_net904),
    .A3(net569),
    .S0(net668),
    .S1(clknet_1_0__leaf_net734),
    .X(net394));
 sky130_fd_sc_hd__mux4_1 c573 (.A0(net375),
    .A1(net962),
    .A2(net800),
    .A3(net569),
    .S0(clknet_1_1__leaf_net734),
    .S1(net889),
    .X(net395));
 sky130_fd_sc_hd__mux4_1 c574 (.A0(net818),
    .A1(clknet_1_0__leaf_net247),
    .A2(clknet_1_0__leaf_net373),
    .A3(net811),
    .S0(net828),
    .S1(net1018),
    .X(net396));
 sky130_fd_sc_hd__mux4_1 c575 (.A0(net236),
    .A1(net795),
    .A2(net1016),
    .A3(net375),
    .S0(net382),
    .S1(net569),
    .X(net397));
 sky130_fd_sc_hd__mux4_1 c576 (.A0(clknet_1_0__leaf_net378),
    .A1(net366),
    .A2(net814),
    .A3(net800),
    .S0(net1024),
    .S1(net579),
    .X(net398));
 sky130_fd_sc_hd__mux4_1 c577 (.A0(net370),
    .A1(net44),
    .A2(clknet_1_1__leaf_net377),
    .A3(net818),
    .S0(clknet_1_1__leaf_net74),
    .S1(clknet_1_1__leaf_net694),
    .X(net399));
 sky130_fd_sc_hd__mux4_2 c578 (.A0(net254),
    .A1(net797),
    .A2(net721),
    .A3(net736),
    .S0(net740),
    .S1(net748),
    .X(net400));
 sky130_fd_sc_hd__mux4_1 c579 (.A0(net800),
    .A1(net400),
    .A2(clknet_1_1__leaf_net893),
    .A3(net573),
    .S0(net605),
    .S1(net992),
    .X(net401));
 sky130_fd_sc_hd__mux4_2 c580 (.A0(net888),
    .A1(net154),
    .A2(net23),
    .A3(net484),
    .S0(net966),
    .S1(net601),
    .X(net402));
 sky130_fd_sc_hd__mux4_1 c581 (.A0(net255),
    .A1(net1042),
    .A2(clknet_1_1__leaf_net673),
    .A3(net721),
    .S0(clknet_1_0__leaf_net751),
    .S1(clknet_1_1__leaf_net752),
    .X(net403));
 sky130_fd_sc_hd__mux4_1 c582 (.A0(clknet_1_0__leaf_net403),
    .A1(net953),
    .A2(clknet_1_1__leaf_net74),
    .A3(net1025),
    .S0(net804),
    .S1(net645),
    .X(net404));
 sky130_fd_sc_hd__mux4_1 c583 (.A0(net1042),
    .A1(net245),
    .A2(clknet_1_0__leaf_net615),
    .A3(net647),
    .S0(net658),
    .S1(clknet_1_0__leaf_net713),
    .X(net405));
 sky130_fd_sc_hd__mux4_1 c584 (.A0(net154),
    .A1(clknet_1_1__leaf_net403),
    .A2(net1001),
    .A3(clknet_1_1__leaf_net296),
    .S0(net1039),
    .S1(clknet_1_1__leaf_net752),
    .X(net406));
 sky130_fd_sc_hd__mux4_1 c585 (.A0(net818),
    .A1(net1013),
    .A2(net647),
    .A3(clknet_1_1__leaf_net733),
    .S0(clknet_1_1__leaf_net734),
    .S1(clknet_1_0__leaf_net753),
    .X(net407));
 sky130_fd_sc_hd__mux4_1 c586 (.A0(net811),
    .A1(clknet_1_1__leaf_net296),
    .A2(net400),
    .A3(net382),
    .S0(net814),
    .S1(net698),
    .X(net408));
 sky130_fd_sc_hd__mux4_1 c587 (.A0(net1027),
    .A1(clknet_1_1__leaf_net401),
    .A2(net780),
    .A3(net254),
    .S0(net995),
    .S1(clknet_1_0__leaf_net752),
    .X(net409));
 sky130_fd_sc_hd__mux4_1 c588 (.A0(clknet_1_1__leaf_net293),
    .A1(net795),
    .A2(net569),
    .A3(net668),
    .S0(clknet_1_0__leaf_net751),
    .S1(net756),
    .X(net410));
 sky130_fd_sc_hd__mux4_1 c589 (.A0(net366),
    .A1(net874),
    .A2(net800),
    .A3(clknet_1_1__leaf_net751),
    .S0(clknet_1_1__leaf_net752),
    .S1(clknet_1_1__leaf_net753),
    .X(net411));
 sky130_fd_sc_hd__mux4_1 c590 (.A0(net287),
    .A1(net400),
    .A2(net967),
    .A3(net658),
    .S0(clknet_1_0__leaf_net752),
    .S1(clknet_1_0__leaf_net753),
    .X(net412));
 sky130_fd_sc_hd__mux4_1 c591 (.A0(clknet_1_0__leaf_net403),
    .A1(clknet_1_1__leaf_net904),
    .A2(net780),
    .A3(clknet_1_0__leaf_net405),
    .S0(net645),
    .S1(net755),
    .X(net413));
 sky130_fd_sc_hd__mux4_1 c592 (.A0(clknet_1_1__leaf_net184),
    .A1(clknet_1_1__leaf_net409),
    .A2(net818),
    .A3(clknet_1_1__leaf_net413),
    .S0(clknet_1_1__leaf_net296),
    .S1(clknet_1_1__leaf_net411),
    .X(net414));
 sky130_fd_sc_hd__mux4_1 c593 (.A0(clknet_1_1__leaf_net394),
    .A1(clknet_1_1__leaf_net413),
    .A2(net573),
    .A3(net605),
    .S0(clknet_1_1__leaf_net695),
    .S1(net755),
    .X(net415));
 sky130_fd_sc_hd__mux4_1 c594 (.A0(net1016),
    .A1(clknet_1_0__leaf_net939),
    .A2(net570),
    .A3(clknet_1_0__leaf_net615),
    .S0(net623),
    .S1(net707),
    .X(net416));
 sky130_fd_sc_hd__mux4_1 c595 (.A0(clknet_1_0__leaf_net390),
    .A1(net841),
    .A2(net570),
    .A3(net681),
    .S0(clknet_1_1__leaf_net694),
    .S1(net723),
    .X(net417));
 sky130_fd_sc_hd__mux4_1 c596 (.A0(net836),
    .A1(net967),
    .A2(net402),
    .A3(clknet_1_0__leaf_net904),
    .S0(net995),
    .S1(net913),
    .X(net418));
 sky130_fd_sc_hd__mux4_1 c597 (.A0(clknet_1_0__leaf_net166),
    .A1(clknet_1_0__leaf_net273),
    .A2(net968),
    .A3(net969),
    .S0(net623),
    .S1(net738),
    .X(net419));
 sky130_fd_sc_hd__mux4_1 c598 (.A0(clknet_1_0__leaf_net296),
    .A1(clknet_1_0__leaf_net904),
    .A2(net805),
    .A3(net1049),
    .S0(net996),
    .S1(net707),
    .X(net420));
 sky130_fd_sc_hd__mux4_1 c599 (.A0(net207),
    .A1(clknet_1_0__leaf_net887),
    .A2(net961),
    .A3(net836),
    .S0(net610),
    .S1(net737),
    .X(net421));
 sky130_fd_sc_hd__mux4_1 c600 (.A0(net795),
    .A1(net255),
    .A2(clknet_1_0__leaf_net277),
    .A3(net650),
    .S0(net883),
    .S1(net996),
    .X(net422));
 sky130_fd_sc_hd__mux4_1 c601 (.A0(clknet_1_0__leaf_net390),
    .A1(net402),
    .A2(net968),
    .A3(clknet_1_0__leaf_net410),
    .S0(net692),
    .S1(clknet_1_1__leaf_net693),
    .X(net423));
 sky130_fd_sc_hd__mux4_1 c602 (.A0(net81),
    .A1(clknet_1_0__leaf_net318),
    .A2(clknet_1_0__leaf_net422),
    .A3(clknet_1_1__leaf_net79),
    .S0(clknet_1_1__leaf_net694),
    .S1(net741),
    .X(net424));
 sky130_fd_sc_hd__mux4_1 c603 (.A0(clknet_1_1__leaf_net79),
    .A1(net1058),
    .A2(clknet_1_0__leaf_net401),
    .A3(net622),
    .S0(net707),
    .S1(net723),
    .X(net425));
 sky130_fd_sc_hd__mux4_1 c604 (.A0(net207),
    .A1(net1016),
    .A2(net1047),
    .A3(net245),
    .S0(net992),
    .S1(net759),
    .X(net426));
 sky130_fd_sc_hd__mux4_1 c605 (.A0(net852),
    .A1(clknet_1_1__leaf_net422),
    .A2(clknet_1_0__leaf_net713),
    .A3(net889),
    .S0(net750),
    .S1(net759),
    .X(net427));
 sky130_fd_sc_hd__mux4_1 c606 (.A0(net841),
    .A1(net809),
    .A2(clknet_1_0__leaf_net422),
    .A3(net402),
    .S0(net876),
    .S1(net759),
    .X(net428));
 sky130_fd_sc_hd__mux4_1 c607 (.A0(clknet_1_0__leaf_net277),
    .A1(clknet_1_1__leaf_net98),
    .A2(net372),
    .A3(net61),
    .S0(net633),
    .S1(net759),
    .X(net429));
 sky130_fd_sc_hd__mux4_1 c608 (.A0(clknet_1_1__leaf_net401),
    .A1(net852),
    .A2(clknet_1_0__leaf_net405),
    .A3(net633),
    .S0(net697),
    .S1(net992),
    .X(net430));
 sky130_fd_sc_hd__mux4_1 c609 (.A0(clknet_1_1__leaf_net157),
    .A1(net1003),
    .A2(clknet_1_0__leaf_net412),
    .A3(net796),
    .S0(net776),
    .S1(net891),
    .X(net431));
 sky130_fd_sc_hd__mux4_1 c610 (.A0(net426),
    .A1(clknet_1_1__leaf_net199),
    .A2(net979),
    .A3(net383),
    .S0(clknet_1_0__leaf_net422),
    .S1(net759),
    .X(net882));
 sky130_fd_sc_hd__mux4_1 c611 (.A0(net1081),
    .A1(net992),
    .A2(net706),
    .A3(net710),
    .S0(net723),
    .S1(net759),
    .X(net432));
 sky130_fd_sc_hd__mux4_1 c612 (.A0(net432),
    .A1(net973),
    .A2(net779),
    .A3(net484),
    .S0(net841),
    .S1(net610),
    .X(net433));
 sky130_fd_sc_hd__mux4_1 c613 (.A0(net431),
    .A1(net428),
    .A2(clknet_1_1__leaf_net318),
    .A3(net432),
    .S0(net646),
    .X(net434));
 sky130_fd_sc_hd__mux4_2 c614 (.A0(net792),
    .A1(net433),
    .A2(net90),
    .A3(net650),
    .S0(net738),
    .S1(net757),
    .X(net435));
 sky130_fd_sc_hd__mux4_1 c615 (.A0(net418),
    .A1(net416),
    .A2(net435),
    .A3(net705),
    .S0(net736),
    .S1(net754),
    .X(net436));
 sky130_fd_sc_hd__mux4_1 c616 (.A0(net54),
    .A1(net999),
    .A2(net1058),
    .A3(net650),
    .S0(net990),
    .S1(net758),
    .X(net437));
 sky130_fd_sc_hd__mux4_1 c617 (.A0(clknet_1_1__leaf_net318),
    .A1(net1028),
    .A2(net90),
    .A3(net605),
    .S0(clknet_1_0__leaf_net713),
    .S1(net988),
    .X(net870));
 sky130_fd_sc_hd__mux4_1 c618 (.A0(clknet_1_1__leaf_net79),
    .A1(net980),
    .A2(net119),
    .A3(net1001),
    .S0(net672),
    .S1(net891),
    .X(net438));
 sky130_fd_sc_hd__mux4_1 c619 (.A0(clknet_1_0__leaf_net231),
    .A1(net969),
    .A2(clknet_1_0__leaf_net939),
    .A3(net672),
    .S0(net683),
    .S1(net988),
    .X(net886));
 sky130_fd_sc_hd__mux4_1 c620 (.A0(clknet_1_0__leaf_net394),
    .A1(net1022),
    .A2(net192),
    .A3(net623),
    .S0(net649),
    .S1(net990),
    .X(net439));
 sky130_fd_sc_hd__mux4_1 c621 (.A0(net430),
    .A1(net805),
    .A2(net643),
    .A3(net650),
    .S0(net988),
    .S1(net737),
    .X(net440));
 sky130_fd_sc_hd__mux4_1 c622 (.A0(net255),
    .A1(clknet_1_1__leaf_net231),
    .A2(clknet_1_1__leaf_net894),
    .A3(net808),
    .S0(net643),
    .S1(net883),
    .X(net441));
 sky130_fd_sc_hd__mux4_1 c623 (.A0(net90),
    .A1(clknet_1_0__leaf_net413),
    .A2(net806),
    .A3(net779),
    .S0(net672),
    .S1(net757),
    .X(net442));
 sky130_fd_sc_hd__mux4_1 c624 (.A0(net335),
    .A1(net968),
    .A2(net1016),
    .A3(clknet_1_0__leaf_net413),
    .S0(net631),
    .S1(net988),
    .X(net443));
 sky130_fd_sc_hd__mux4_1 c625 (.A0(net440),
    .A1(clknet_1_1__leaf_net895),
    .A2(net635),
    .A3(net931),
    .S0(net746),
    .S1(net750),
    .X(net444));
 sky130_fd_sc_hd__mux4_1 c626 (.A0(net954),
    .A1(clknet_1_0__leaf_net401),
    .A2(clknet_1_0__leaf_net318),
    .A3(net980),
    .S0(net192),
    .S1(clknet_1_0__leaf_net394),
    .X(net445));
 sky130_fd_sc_hd__mux4_1 c627 (.A0(net383),
    .A1(net821),
    .A2(net119),
    .A3(net3),
    .S0(net618),
    .S1(net745),
    .X(net446));
 sky130_fd_sc_hd__mux4_1 c628 (.A0(net821),
    .A1(net54),
    .A2(net806),
    .A3(clknet_1_0__leaf_net346),
    .S0(net618),
    .S1(net760),
    .X(net447));
 sky130_fd_sc_hd__mux4_1 c629 (.A0(net1028),
    .A1(clknet_1_0__leaf_net409),
    .A2(clknet_1_1__leaf_net333),
    .A3(clknet_1_1__leaf_net651),
    .S0(net988),
    .S1(net741),
    .X(net884));
 sky130_fd_sc_hd__mux4_1 c630 (.A0(net419),
    .A1(net329),
    .A2(net968),
    .A3(net119),
    .S0(clknet_1_0__leaf_net893),
    .S1(net990),
    .X(net448));
 sky130_fd_sc_hd__mux4_1 c631 (.A0(net969),
    .A1(clknet_1_0__leaf_net333),
    .A2(net649),
    .A3(net650),
    .S0(clknet_1_1__leaf_net651),
    .S1(net658),
    .X(net449));
 sky130_fd_sc_hd__mux4_1 c632 (.A0(net417),
    .A1(net435),
    .A2(net962),
    .A3(clknet_1_0__leaf_net939),
    .S0(net814),
    .S1(net570),
    .X(net450));
 sky130_fd_sc_hd__mux4_1 c633 (.A0(clknet_1_1__leaf_net307),
    .A1(net427),
    .A2(net797),
    .A3(net246),
    .S0(net861),
    .S1(clknet_1_1__leaf_net895),
    .X(net451));
 sky130_fd_sc_hd__mux4_1 c634 (.A0(clknet_1_0__leaf_net346),
    .A1(net821),
    .A2(clknet_1_0__leaf_net307),
    .A3(clknet_1_0__leaf_net409),
    .S0(clknet_1_1__leaf_net616),
    .S1(net643),
    .X(net452));
 sky130_fd_sc_hd__mux4_1 c635 (.A0(net1020),
    .A1(net635),
    .A2(net655),
    .A3(net658),
    .S0(net737),
    .S1(net760),
    .X(net453));
 sky130_fd_sc_hd__mux4_1 c636 (.A0(net808),
    .A1(net450),
    .A2(net453),
    .A3(clknet_1_1__leaf_net895),
    .S0(net655),
    .S1(net760),
    .X(net454));
 sky130_fd_sc_hd__mux4_1 c637 (.A0(net449),
    .A1(net1058),
    .A2(net971),
    .A3(net649),
    .S0(net683),
    .S1(net758),
    .X(net455));
 sky130_fd_sc_hd__a2111o_2 c660 (.A1(net1037),
    .A2(net350),
    .B1(net979),
    .C1(net1004),
    .D1(net688),
    .X(net456));
 sky130_fd_sc_hd__a2111o_2 c661 (.A1(net345),
    .A2(net359),
    .B1(net343),
    .C1(net1010),
    .D1(net356),
    .X(net457));
 sky130_fd_sc_hd__a2111o_1 c662 (.A1(net457),
    .A2(net986),
    .B1(net349),
    .C1(net359),
    .D1(clknet_1_1__leaf_net714),
    .X(net458));
 sky130_fd_sc_hd__a2111o_1 c663 (.A1(net456),
    .A2(clknet_1_1__leaf_net458),
    .B1(net1041),
    .C1(net688),
    .D1(clknet_1_1__leaf_net714),
    .X(net459));
 sky130_fd_sc_hd__mux4_1 c664 (.A0(net344),
    .A1(net1027),
    .A2(net126),
    .A3(net347),
    .S0(net132),
    .S1(clknet_1_1__leaf_net714),
    .X(net460));
 sky130_fd_sc_hd__a2111o_1 c665 (.A1(net456),
    .A2(net143),
    .B1(net976),
    .C1(net1042),
    .D1(net359),
    .X(net461));
 sky130_fd_sc_hd__a2111o_1 c666 (.A1(net461),
    .A2(net457),
    .B1(net1083),
    .C1(clknet_1_1__leaf_net460),
    .D1(net361),
    .X(net462));
 sky130_fd_sc_hd__mux4_1 c667 (.A0(net1027),
    .A1(net1033),
    .A2(clknet_1_1__leaf_net462),
    .A3(net233),
    .S0(net660),
    .S1(clknet_1_1__leaf_net712),
    .X(net463));
 sky130_fd_sc_hd__mux4_2 c668 (.A0(net1025),
    .A1(net457),
    .A2(net1008),
    .A3(net1004),
    .S0(net361),
    .S1(net688),
    .X(net464));
 sky130_fd_sc_hd__a2111o_1 c669 (.A1(net457),
    .A2(net456),
    .B1(net1037),
    .C1(net972),
    .D1(clknet_1_1__leaf_net712),
    .X(net465));
 sky130_fd_sc_hd__a2111o_1 c670 (.A1(net133),
    .A2(clknet_1_1__leaf_net353),
    .B1(net464),
    .C1(clknet_1_0__leaf_net462),
    .D1(net35),
    .X(net466));
 sky130_fd_sc_hd__a2111o_1 c671 (.A1(clknet_1_0__leaf_net462),
    .A2(net457),
    .B1(net356),
    .C1(net1008),
    .D1(net1004),
    .X(net467));
 sky130_fd_sc_hd__a2111o_1 c672 (.A1(net456),
    .A2(clknet_1_1__leaf_net462),
    .B1(net464),
    .C1(net660),
    .D1(clknet_1_1__leaf_net714),
    .X(net468));
 sky130_fd_sc_hd__mux4_1 c673 (.A0(net137),
    .A1(net1008),
    .A2(clknet_1_1__leaf_net462),
    .A3(net654),
    .S0(net688),
    .S1(clknet_1_1__leaf_net714),
    .X(net469));
 sky130_fd_sc_hd__mux4_1 c674 (.A0(net357),
    .A1(clknet_1_1__leaf_net247),
    .A2(net1008),
    .A3(net578),
    .S0(net654),
    .S1(net663),
    .X(net470));
 sky130_fd_sc_hd__a2111o_1 c675 (.A1(net464),
    .A2(net1027),
    .B1(clknet_1_0__leaf_net462),
    .C1(net664),
    .D1(net1108),
    .X(net471));
 sky130_fd_sc_hd__mux4_2 c676 (.A0(net364),
    .A1(net132),
    .A2(net136),
    .A3(net578),
    .S0(net664),
    .S1(net762),
    .X(net472));
 sky130_fd_sc_hd__mux4_1 c677 (.A0(net359),
    .A1(net951),
    .A2(net1026),
    .A3(net578),
    .S0(net664),
    .S1(net762),
    .X(net473));
 sky130_fd_sc_hd__mux4_2 c678 (.A0(net456),
    .A1(net959),
    .A2(net457),
    .A3(net660),
    .S0(net762),
    .S1(net763),
    .X(net474));
 sky130_fd_sc_hd__mux4_1 c679 (.A0(net461),
    .A1(net474),
    .A2(net143),
    .A3(net137),
    .S0(net654),
    .S1(net761),
    .X(net475));
 sky130_fd_sc_hd__mux4_1 c680 (.A0(net474),
    .A1(net143),
    .A2(net596),
    .A3(net689),
    .S0(net761),
    .S1(net763),
    .X(net476));
 sky130_fd_sc_hd__mux4_1 c681 (.A0(net233),
    .A1(clknet_1_1__leaf_net354),
    .A2(net457),
    .A3(net578),
    .S0(net596),
    .S1(clknet_1_1__leaf_net712),
    .X(net477));
 sky130_fd_sc_hd__mux4_1 c682 (.A0(net1026),
    .A1(net387),
    .A2(net957),
    .A3(net1020),
    .S0(net233),
    .S1(net472),
    .X(net478));
 sky130_fd_sc_hd__mux4_2 c683 (.A0(net25),
    .A1(net456),
    .A2(net1026),
    .A3(net1016),
    .S0(net472),
    .S1(net972),
    .X(net479));
 sky130_fd_sc_hd__mux4_1 c684 (.A0(net479),
    .A1(net959),
    .A2(net126),
    .A3(net369),
    .S0(net731),
    .S1(net761),
    .X(net480));
 sky130_fd_sc_hd__mux4_1 c685 (.A0(net480),
    .A1(net972),
    .A2(net360),
    .A3(net977),
    .S0(net782),
    .S1(net779),
    .X(net481));
 sky130_fd_sc_hd__mux4_1 c686 (.A0(net1025),
    .A1(clknet_1_0__leaf_net465),
    .A2(net364),
    .A3(net1027),
    .S0(net730),
    .S1(net765),
    .X(net482));
 sky130_fd_sc_hd__mux4_1 c687 (.A0(clknet_1_1__leaf_net465),
    .A1(net233),
    .A2(net480),
    .A3(net456),
    .S0(clknet_1_1__leaf_net458),
    .S1(net1020),
    .X(net483));
 sky130_fd_sc_hd__mux4_2 c688 (.A0(net963),
    .A1(clknet_1_0__leaf_net353),
    .A2(net1020),
    .S0(net993),
    .S1(net765),
    .X(net641));
 sky130_fd_sc_hd__mux4_1 c689 (.A0(net25),
    .A1(net957),
    .A2(net687),
    .A3(net993),
    .S0(net731),
    .S1(net764),
    .X(net485));
 sky130_fd_sc_hd__mux4_1 c690 (.A0(net126),
    .A1(net808),
    .A2(net35),
    .A3(net781),
    .S0(net993),
    .S1(net768),
    .X(net486));
 sky130_fd_sc_hd__mux4_1 c691 (.A0(clknet_1_1__leaf_net276),
    .A1(net375),
    .A2(net486),
    .A3(net959),
    .S0(net664),
    .S1(net768),
    .X(net487));
 sky130_fd_sc_hd__mux4_2 c692 (.A0(net986),
    .A1(net479),
    .A2(net472),
    .A3(net804),
    .S0(net963),
    .S1(net768),
    .X(net488));
 sky130_fd_sc_hd__mux4_1 c693 (.A0(clknet_1_0__leaf_net354),
    .A1(net486),
    .A2(net474),
    .A3(clknet_1_1__leaf_net693),
    .S0(net767),
    .S1(net1067),
    .X(net489));
 sky130_fd_sc_hd__mux4_1 c694 (.A0(net1008),
    .A1(net480),
    .A2(net1078),
    .A3(net25),
    .S0(net993),
    .S1(net1067),
    .X(net490));
 sky130_fd_sc_hd__mux4_1 c695 (.A0(net486),
    .A1(net360),
    .A2(clknet_1_1__leaf_net247),
    .A3(net488),
    .S0(net993),
    .S1(net1067),
    .X(net491));
 sky130_fd_sc_hd__mux4_1 c696 (.A0(net1065),
    .A1(net480),
    .A2(net1020),
    .A3(net571),
    .S0(net659),
    .S1(net768),
    .X(net492));
 sky130_fd_sc_hd__mux4_2 c697 (.A0(net976),
    .A1(net1081),
    .A2(net642),
    .A3(net659),
    .S0(net691),
    .S1(net768),
    .X(net493));
 sky130_fd_sc_hd__mux4_1 c698 (.A0(net486),
    .A1(net493),
    .A2(net595),
    .A3(net617),
    .S0(net766),
    .S1(net768),
    .X(net494));
 sky130_fd_sc_hd__mux4_2 c699 (.A0(net1016),
    .A1(net493),
    .A2(net571),
    .A3(net595),
    .S0(net642),
    .S1(net659),
    .X(net495));
 sky130_fd_sc_hd__mux4_1 c700 (.A0(net959),
    .A1(net493),
    .A2(net479),
    .A3(clknet_1_0__leaf_net392),
    .S0(net617),
    .S1(net642),
    .X(net496));
 sky130_fd_sc_hd__mux4_1 c701 (.A0(clknet_1_1__leaf_net496),
    .A1(net495),
    .A2(net493),
    .A3(net234),
    .S0(net1041),
    .S1(net766),
    .X(net497));
 sky130_fd_sc_hd__mux4_1 c702 (.A0(net479),
    .A1(net1008),
    .A2(net493),
    .A3(net963),
    .S0(net571),
    .S1(net718),
    .X(net498));
 sky130_fd_sc_hd__mux4_1 c703 (.A0(clknet_1_1__leaf_net392),
    .A1(net488),
    .A2(clknet_1_0__leaf_net496),
    .A3(net571),
    .S0(net699),
    .S1(net769),
    .X(net499));
 sky130_fd_sc_hd__mux4_1 c704 (.A0(net494),
    .A1(net874),
    .A2(net35),
    .A3(net963),
    .S0(net700),
    .S1(net718),
    .X(net500));
 sky130_fd_sc_hd__mux4_1 c705 (.A0(net21),
    .A1(net68),
    .A2(net1081),
    .A3(net996),
    .S0(net736),
    .S1(net770),
    .X(net501));
 sky130_fd_sc_hd__mux4_2 c706 (.A0(net33),
    .A1(net362),
    .A2(net1025),
    .A3(clknet_1_0__leaf_net399),
    .S0(net663),
    .S1(net737),
    .X(net502));
 sky130_fd_sc_hd__mux4_1 c707 (.A0(net784),
    .A1(net402),
    .A2(clknet_1_0__leaf_net502),
    .A3(clknet_1_1__leaf_net904),
    .S0(net362),
    .S1(net658),
    .X(net503));
 sky130_fd_sc_hd__mux4_1 c708 (.A0(clknet_1_0__leaf_net460),
    .A1(net1052),
    .A2(clknet_1_1__leaf_net178),
    .A3(net1062),
    .S0(net761),
    .S1(net767),
    .X(net504));
 sky130_fd_sc_hd__mux4_1 c709 (.A0(clknet_1_1__leaf_net178),
    .A1(net809),
    .A2(net781),
    .A3(net666),
    .S0(net699),
    .S1(net739),
    .X(net505));
 sky130_fd_sc_hd__mux4_1 c710 (.A0(net498),
    .A1(net1015),
    .A2(net375),
    .A3(net666),
    .S0(clknet_1_1__leaf_net675),
    .S1(net769),
    .X(net506));
 sky130_fd_sc_hd__mux4_1 c711 (.A0(clknet_1_1__leaf_net504),
    .A1(net1020),
    .A2(net1003),
    .A3(net617),
    .S0(clknet_1_1__leaf_net673),
    .S1(net756),
    .X(net507));
 sky130_fd_sc_hd__mux4_1 c712 (.A0(net1025),
    .A1(net494),
    .A2(clknet_1_1__leaf_net502),
    .A3(net370),
    .S0(clknet_1_1__leaf_net712),
    .S1(clknet_1_1__leaf_net734),
    .X(net508));
 sky130_fd_sc_hd__mux4_1 c713 (.A0(net808),
    .A1(net501),
    .A2(net350),
    .A3(net37),
    .S0(clknet_1_0__leaf_net641),
    .S1(net721),
    .X(net509));
 sky130_fd_sc_hd__mux4_1 c714 (.A0(clknet_1_1__leaf_net373),
    .A1(clknet_1_1__leaf_net505),
    .A2(net498),
    .A3(clknet_1_0__leaf_net502),
    .S0(clknet_1_1__leaf_net178),
    .S1(clknet_1_1__leaf_net673),
    .X(net510));
 sky130_fd_sc_hd__mux4_1 c715 (.A0(net1041),
    .A1(net68),
    .A2(clknet_1_1__leaf_net410),
    .A3(net602),
    .S0(clknet_1_1__leaf_net733),
    .S1(net750),
    .X(net511));
 sky130_fd_sc_hd__mux4_1 c716 (.A0(clknet_1_1__leaf_net502),
    .A1(net498),
    .A2(net493),
    .A3(clknet_1_1__leaf_net712),
    .S0(net761),
    .S1(net763),
    .X(net512));
 sky130_fd_sc_hd__mux4_1 c717 (.A0(net503),
    .A1(net508),
    .A2(net494),
    .A3(net350),
    .S0(net361),
    .S1(net602),
    .X(net513));
 sky130_fd_sc_hd__mux4_1 c718 (.A0(clknet_1_1__leaf_net399),
    .A1(net1053),
    .A2(net957),
    .A3(net808),
    .S0(clknet_1_1__leaf_net512),
    .S1(clknet_1_1__leaf_net712),
    .X(net514));
 sky130_fd_sc_hd__mux4_1 c719 (.A0(net350),
    .A1(net35),
    .A2(clknet_1_1__leaf_net512),
    .A3(net1025),
    .S0(net653),
    .S1(clknet_1_1__leaf_net733),
    .X(net515));
 sky130_fd_sc_hd__mux4_1 c720 (.A0(net515),
    .A1(net37),
    .A2(clknet_1_1__leaf_net178),
    .A3(net493),
    .S0(clknet_1_1__leaf_net512),
    .S1(net769),
    .X(net516));
 sky130_fd_sc_hd__mux4_2 c721 (.A0(clknet_1_1__leaf_net377),
    .A1(clknet_1_1__leaf_net502),
    .A2(net349),
    .A3(net663),
    .S0(clknet_1_1__leaf_net753),
    .S1(net769),
    .X(net517));
 sky130_fd_sc_hd__mux4_2 c722 (.A0(clknet_1_1__leaf_net178),
    .A1(clknet_1_1__leaf_net641),
    .A2(net645),
    .A3(net666),
    .S0(net750),
    .S1(net769),
    .X(net518));
 sky130_fd_sc_hd__mux4_1 c723 (.A0(net370),
    .A1(clknet_1_1__leaf_net247),
    .A2(clknet_1_1__leaf_net512),
    .A3(clknet_1_1__leaf_net502),
    .S1(net718),
    .X(net519));
 sky130_fd_sc_hd__mux4_1 c724 (.A0(clknet_1_0__leaf_net512),
    .A1(net602),
    .A2(net638),
    .A3(net915),
    .S0(net761),
    .S1(net763),
    .X(net520));
 sky130_fd_sc_hd__mux4_1 c725 (.A0(net520),
    .A1(clknet_1_1__leaf_net517),
    .A2(net35),
    .A3(clknet_1_0__leaf_net460),
    .S0(net776),
    .S1(net731),
    .X(net521));
 sky130_fd_sc_hd__mux4_2 c726 (.A0(net776),
    .A1(clknet_1_0__leaf_net517),
    .A2(net787),
    .A3(clknet_1_0__leaf_net411),
    .S0(clknet_1_0__leaf_net939),
    .S1(net624),
    .X(net522));
 sky130_fd_sc_hd__mux4_1 c727 (.A0(clknet_1_1__leaf_net100),
    .A1(net809),
    .A2(net362),
    .A3(clknet_1_1__leaf_net522),
    .S0(net624),
    .S1(net740),
    .X(net523));
 sky130_fd_sc_hd__mux4_1 c728 (.A0(clknet_1_1__leaf_net405),
    .A1(clknet_1_0__leaf_net512),
    .A2(net488),
    .A3(clknet_1_1__leaf_net422),
    .S0(net730),
    .S1(net739),
    .X(net930));
 sky130_fd_sc_hd__mux4_2 c729 (.A0(clknet_1_0__leaf_net458),
    .A1(clknet_1_1__leaf_net310),
    .A2(net842),
    .A3(net915),
    .S0(net664),
    .S1(net770),
    .X(net524));
 sky130_fd_sc_hd__mux4_1 c730 (.A0(clknet_1_1__leaf_net422),
    .A1(clknet_1_0__leaf_net458),
    .A2(net952),
    .A3(clknet_1_1__leaf_net904),
    .S0(net639),
    .S1(net763),
    .X(net525));
 sky130_fd_sc_hd__mux4_2 c731 (.A0(net88),
    .A1(clknet_1_1__leaf_net518),
    .A2(net804),
    .A3(net902),
    .S0(net622),
    .S1(net731),
    .X(net526));
 sky130_fd_sc_hd__mux4_1 c732 (.A0(net501),
    .A1(net30),
    .A2(net1033),
    .A3(net667),
    .S0(net730),
    .S1(net763),
    .X(net527));
 sky130_fd_sc_hd__mux4_1 c733 (.A0(clknet_1_1__leaf_net73),
    .A1(net1033),
    .A2(net842),
    .A3(clknet_1_1__leaf_net247),
    .S0(net37),
    .S1(net873),
    .X(net528));
 sky130_fd_sc_hd__mux4_1 c734 (.A0(net796),
    .A1(clknet_1_0__leaf_net518),
    .A2(net400),
    .A3(net622),
    .S0(net996),
    .S1(net731),
    .X(net529));
 sky130_fd_sc_hd__mux4_1 c735 (.A0(clknet_1_1__leaf_net285),
    .A1(net246),
    .A2(clknet_1_1__leaf_net73),
    .A3(net663),
    .S0(net681),
    .S1(net996),
    .X(net530));
 sky130_fd_sc_hd__mux4_1 c736 (.A0(net472),
    .A1(clknet_1_1__leaf_net522),
    .A2(net962),
    .A3(net877),
    .S0(net669),
    .S1(clknet_1_1__leaf_net675),
    .X(net531));
 sky130_fd_sc_hd__mux4_1 c737 (.A0(clknet_1_0__leaf_net502),
    .A1(net472),
    .A2(net1001),
    .A3(net602),
    .S0(net730),
    .S1(net741),
    .X(net532));
 sky130_fd_sc_hd__mux4_1 c738 (.A0(net495),
    .A1(net362),
    .A2(clknet_1_1__leaf_net73),
    .A3(net877),
    .S0(net656),
    .S1(net667),
    .X(net533));
 sky130_fd_sc_hd__mux4_1 c739 (.A0(net493),
    .A1(clknet_1_0__leaf_net517),
    .A2(net500),
    .A3(clknet_1_1__leaf_net247),
    .S0(net976),
    .S1(net770),
    .X(net534));
 sky130_fd_sc_hd__mux4_1 c740 (.A0(clknet_1_0__leaf_net532),
    .A1(net977),
    .A2(net488),
    .A3(net362),
    .S0(clknet_1_1__leaf_net530),
    .S1(net667),
    .X(net535));
 sky130_fd_sc_hd__mux4_1 c741 (.A0(clknet_1_1__leaf_net73),
    .A1(net33),
    .A2(net902),
    .A3(net605),
    .S0(net915),
    .S1(net996),
    .X(net536));
 sky130_fd_sc_hd__mux4_1 c742 (.A0(net488),
    .A1(net402),
    .A2(clknet_1_0__leaf_net512),
    .A3(clknet_1_0__leaf_net522),
    .S0(net657),
    .S1(net995),
    .X(net537));
 sky130_fd_sc_hd__mux4_1 c743 (.A0(net400),
    .A1(clknet_1_0__leaf_net522),
    .A2(net639),
    .A3(net669),
    .S0(net995),
    .S1(net913),
    .X(net538));
 sky130_fd_sc_hd__mux4_1 c744 (.A0(clknet_1_1__leaf_net412),
    .A1(clknet_1_1__leaf_net522),
    .A2(net493),
    .A3(net664),
    .S0(clknet_1_1__leaf_net675),
    .S1(net700),
    .X(net539));
 sky130_fd_sc_hd__mux4_1 c745 (.A0(clknet_1_0__leaf_net505),
    .A1(net533),
    .A2(clknet_1_1__leaf_net509),
    .A3(clknet_1_1__leaf_net530),
    .S0(net784),
    .S1(net657),
    .X(net540));
 sky130_fd_sc_hd__mux4_1 c746 (.A0(clknet_1_0__leaf_net410),
    .A1(net429),
    .A2(net536),
    .A3(clknet_1_1__leaf_net532),
    .S0(net979),
    .S1(net656),
    .X(net541));
 sky130_fd_sc_hd__mux4_1 c747 (.A0(clknet_1_0__leaf_net530),
    .A1(net622),
    .A2(net638),
    .A3(net656),
    .S0(net657),
    .S1(net731),
    .X(net542));
 sky130_fd_sc_hd__mux4_1 c748 (.A0(net362),
    .A1(net867),
    .A2(net653),
    .A3(net658),
    .S0(net683),
    .S1(net996),
    .X(net543));
 sky130_fd_sc_hd__mux4_1 c749 (.A0(net842),
    .A1(net1048),
    .A2(net861),
    .A3(net773),
    .S0(net1015),
    .S1(net3),
    .X(net544));
 sky130_fd_sc_hd__mux4_1 c750 (.A0(clknet_1_1__leaf_net333),
    .A1(clknet_1_1__leaf_net535),
    .A2(net1005),
    .A3(clknet_1_0__leaf_net504),
    .S0(clknet_1_1__leaf_net407),
    .S1(net741),
    .X(net545));
 sky130_fd_sc_hd__mux4_1 c751 (.A0(net1),
    .A1(net543),
    .A2(net842),
    .A3(net435),
    .S0(net632),
    .S1(net750),
    .X(net546));
 sky130_fd_sc_hd__mux4_1 c752 (.A0(net474),
    .A1(net979),
    .A2(net859),
    .A3(net435),
    .S0(net605),
    .S1(net740),
    .X(net547));
 sky130_fd_sc_hd__mux4_1 c753 (.A0(net192),
    .A1(net957),
    .A2(net542),
    .A3(net848),
    .S0(clknet_1_1__leaf_net693),
    .S1(net760),
    .X(net548));
 sky130_fd_sc_hd__mux4_1 c754 (.A0(net867),
    .A1(clknet_1_0__leaf_net407),
    .A2(net976),
    .A3(net804),
    .S0(net877),
    .S1(net646),
    .X(net549));
 sky130_fd_sc_hd__mux4_1 c755 (.A0(clknet_1_0__leaf_net411),
    .A1(net857),
    .A2(net527),
    .A3(net435),
    .S0(clknet_1_1__leaf_net616),
    .S1(net681),
    .X(net550));
 sky130_fd_sc_hd__mux4_1 c756 (.A0(clknet_1_0__leaf_net522),
    .A1(net546),
    .A2(net804),
    .A3(clknet_1_0__leaf_net549),
    .S0(net653),
    .S1(net770),
    .X(net551));
 sky130_fd_sc_hd__mux4_1 c757 (.A0(clknet_1_0__leaf_net549),
    .A1(net119),
    .A2(net1062),
    .A3(net632),
    .S0(net639),
    .S1(net656),
    .X(net552));
 sky130_fd_sc_hd__mux4_1 c758 (.A0(clknet_1_0__leaf_net310),
    .A1(net441),
    .A2(net552),
    .A3(net1015),
    .S0(net1040),
    .S1(clknet_1_1__leaf_net675),
    .X(net553));
 sky130_fd_sc_hd__mux4_1 c759 (.A0(net810),
    .A1(clknet_1_0__leaf_net509),
    .A2(net979),
    .A3(clknet_1_1__leaf_net549),
    .S0(net878),
    .S1(net875),
    .X(net554));
 sky130_fd_sc_hd__a2111o_1 c760 (.A1(net773),
    .A2(clknet_1_1__leaf_net549),
    .B1(net362),
    .C1(net931),
    .D1(net878),
    .X(net555));
 sky130_fd_sc_hd__mux4_1 c761 (.A0(clknet_1_1__leaf_net247),
    .A1(net952),
    .A2(clknet_1_1__leaf_net83),
    .A3(net1003),
    .S0(net624),
    .S1(clknet_1_1__leaf_net675),
    .X(net556));
 sky130_fd_sc_hd__mux4_1 c762 (.A0(net3),
    .A1(net435),
    .A2(clknet_1_1__leaf_net675),
    .A3(net681),
    .S0(clknet_1_1__leaf_net693),
    .S1(net740),
    .X(net557));
 sky130_fd_sc_hd__mux4_1 c763 (.A0(net554),
    .A1(net962),
    .A2(net787),
    .A3(net550),
    .S0(net1),
    .S1(clknet_1_1__leaf_net693),
    .X(net558));
 sky130_fd_sc_hd__mux4_1 c764 (.A0(net544),
    .A1(net435),
    .A2(net558),
    .A3(clknet_1_0__leaf_net535),
    .S0(net635),
    .S1(net754),
    .X(net559));
 sky130_fd_sc_hd__mux4_1 c765 (.A0(net33),
    .A1(net859),
    .A2(net446),
    .A3(net957),
    .S0(net495),
    .S1(net657),
    .X(net560));
 sky130_fd_sc_hd__mux4_1 c766 (.A0(net246),
    .A1(net455),
    .A2(clknet_1_0__leaf_net530),
    .A3(net1003),
    .S0(net737),
    .S1(net760),
    .X(net561));
 sky130_fd_sc_hd__a2111o_1 c767 (.A1(net495),
    .A2(net557),
    .B1(net362),
    .C1(net631),
    .D1(net663),
    .X(net562));
 sky130_fd_sc_hd__mux4_1 c768 (.A0(net555),
    .A1(net848),
    .A2(clknet_1_0__leaf_net504),
    .A3(net562),
    .S0(net1032),
    .S1(net1020),
    .X(net563));
 sky130_fd_sc_hd__mux4_1 c769 (.A0(net971),
    .A1(clknet_1_0__leaf_net199),
    .A2(net561),
    .A3(net435),
    .S0(net878),
    .S1(net663));
 sky130_fd_sc_hd__and2_0 merge790 (.A(net324),
    .B(net330),
    .X(net564));
 sky130_fd_sc_hd__and2_0 merge791 (.A(net290),
    .B(net291),
    .X(net565));
 sky130_fd_sc_hd__and2_0 merge792 (.A(net423),
    .B(net424),
    .X(net566));
 sky130_fd_sc_hd__dfrbp_1 merge793 (.CLK(clknet_4_6_0_clk),
    .D(net187),
    .RESET_B(net171),
    .Q(net568),
    .Q_N(net567));
 sky130_fd_sc_hd__dfrbp_1 merge794 (.CLK(clknet_4_0_0_clk),
    .D(net102),
    .RESET_B(net106),
    .Q(net933),
    .Q_N(net942));
 sky130_fd_sc_hd__dfrtn_1 merge795 (.CLK_N(clknet_4_8_0_clk),
    .D(net304),
    .RESET_B(net308),
    .Q(net902));
 sky130_fd_sc_hd__dfrtp_4 merge796 (.CLK(clknet_4_14_0_clk),
    .D(net380),
    .RESET_B(net384),
    .Q(net569));
 sky130_fd_sc_hd__dfrtp_4 merge797 (.CLK(clknet_4_1_0_clk),
    .D(net101),
    .RESET_B(net94),
    .Q(net570));
 sky130_fd_sc_hd__dfrtp_1 merge798 (.CLK(clknet_4_14_0_clk),
    .D(net487),
    .RESET_B(net491),
    .Q(net571));
 sky130_fd_sc_hd__dfsbp_2 merge799 (.CLK(clknet_4_1_0_clk),
    .D(net67),
    .SET_B(net63),
    .Q(net573),
    .Q_N(net572));
 sky130_fd_sc_hd__and2_0 merge800 (.A(net437),
    .B(net438),
    .X(net574));
 sky130_fd_sc_hd__dfsbp_2 merge801 (.CLK(clknet_4_7_0_clk),
    .D(net140),
    .SET_B(net141),
    .Q(net576),
    .Q_N(net575));
 sky130_fd_sc_hd__and2_0 merge802 (.A(net196),
    .B(net197),
    .X(net577));
 sky130_fd_sc_hd__dfstp_2 merge803 (.CLK(clknet_4_5_0_clk),
    .D(net165),
    .SET_B(net151),
    .Q(net909));
 sky130_fd_sc_hd__dfstp_1 merge804 (.CLK(clknet_4_15_0_clk),
    .D(net466),
    .SET_B(net471),
    .Q(net578));
 sky130_fd_sc_hd__dfstp_2 merge805 (.CLK(clknet_4_15_0_clk),
    .D(net355),
    .SET_B(net358),
    .Q(net579));
 sky130_fd_sc_hd__and2_0 merge806 (.A(net232),
    .B(net216),
    .X(net580));
 sky130_fd_sc_hd__and2_0 merge807 (.A(net506),
    .B(net514),
    .X(net581));
 sky130_fd_sc_hd__and2_0 merge808 (.A(net545),
    .B(net547),
    .X(net582));
 sky130_fd_sc_hd__and2_0 merge809 (.A(net415),
    .B(net396),
    .X(net583));
 sky130_fd_sc_hd__and2_4 merge810 (.A(net523),
    .B(net524),
    .X(net584));
 sky130_fd_sc_hd__dlrbn_2 merge811 (.D(net41),
    .GATE_N(clknet_4_5_0_clk),
    .RESET_B(net52),
    .Q(net586),
    .Q_N(net585));
 sky130_fd_sc_hd__and2_0 merge812 (.A(net122),
    .B(net123),
    .X(net587));
 sky130_fd_sc_hd__dlrbn_1 merge813 (.D(net261),
    .GATE_N(clknet_4_13_0_clk),
    .RESET_B(net248),
    .Q(net589),
    .Q_N(net588));
 sky130_fd_sc_hd__dlrbp_1 merge814 (.D(net278),
    .GATE(clknet_4_12_0_clk),
    .RESET_B(net281),
    .Q(net591),
    .Q_N(net590));
 sky130_fd_sc_hd__and2_0 merge815 (.A(net516),
    .B(net541),
    .X(net592));
 sky130_fd_sc_hd__and2_0 merge816 (.A(net534),
    .B(net525),
    .X(net593));
 sky130_fd_sc_hd__and2_0 merge817 (.A(net445),
    .B(net563),
    .X(net594));
 sky130_fd_sc_hd__dlrbp_1 merge818 (.D(net475),
    .GATE(clknet_4_15_0_clk),
    .RESET_B(net492),
    .Q(net596),
    .Q_N(net595));
 sky130_fd_sc_hd__and2_0 merge819 (.A(net332),
    .B(net340),
    .X(net597));
 sky130_fd_sc_hd__and2_0 merge820 (.A(net528),
    .B(net560),
    .X(net598));
 sky130_fd_sc_hd__and2_0 merge821 (.A(net300),
    .B(net298),
    .X(net599));
 sky130_fd_sc_hd__and2_0 merge822 (.A(net107),
    .B(net108),
    .X(net600));
 sky130_fd_sc_hd__dlrtn_1 merge823 (.GATE_N(clknet_4_4_0_clk),
    .RESET_B(net181),
    .Q(net188));
 sky130_fd_sc_hd__dlrtn_1 merge824 (.D(net477),
    .GATE_N(clknet_4_11_0_clk),
    .RESET_B(net581),
    .Q(net602));
 sky130_fd_sc_hd__and2_0 merge825 (.A(net114),
    .B(net115),
    .X(net603));
 sky130_fd_sc_hd__dlrtn_2 merge826 (.D(net265),
    .GATE_N(clknet_4_12_0_clk),
    .RESET_B(net282),
    .Q(net604));
 sky130_fd_sc_hd__dlrtp_2 merge827 (.D(net414),
    .GATE(clknet_4_11_0_clk),
    .RESET_B(net395),
    .Q(net605));
 sky130_fd_sc_hd__and2_0 merge828 (.A(net442),
    .B(net337),
    .X(net606));
 sky130_fd_sc_hd__dlrtp_4 merge829 (.D(net99),
    .GATE(clknet_4_1_0_clk),
    .RESET_B(net96),
    .Q(net607));
 sky130_fd_sc_hd__dlrtp_2 merge830 (.D(net587),
    .GATE(clknet_4_0_0_clk),
    .RESET_B(net229),
    .Q(net907));
 sky130_fd_sc_hd__and2_0 merge831 (.A(net439),
    .B(net559),
    .X(net608));
 sky130_fd_sc_hd__edfxbp_1 merge832 (.CLK(clknet_4_2_0_clk),
    .D(net316),
    .DE(net314),
    .Q(net610),
    .Q_N(net609));
 sky130_fd_sc_hd__edfxtp_1 merge833 (.CLK(clknet_4_0_0_clk),
    .D(net228),
    .DE(net226),
    .Q(net611));
 sky130_fd_sc_hd__and2_0 merge834 (.A(net339),
    .B(net447),
    .X(net612));
 sky130_fd_sc_hd__sdlclkp_1 merge835 (.CLK(clknet_4_3_0_clk),
    .GATE(net201),
    .SCE(net177),
    .GCLK(net613));
 sky130_fd_sc_hd__and2_0 merge836 (.A(net448),
    .B(net452),
    .X(net614));
 sky130_fd_sc_hd__sdlclkp_2 merge837 (.CLK(clknet_4_14_0_clk),
    .GATE(net388),
    .SCE(net386),
    .GCLK(net615));
 sky130_fd_sc_hd__sdlclkp_4 merge838 (.CLK(clknet_4_8_0_clk),
    .GATE(net612),
    .SCE(net597),
    .GCLK(net616));
 sky130_fd_sc_hd__dfrbp_2 merge839 (.CLK(clknet_4_14_0_clk),
    .D(net363),
    .RESET_B(net490),
    .Q(net618),
    .Q_N(net617));
 sky130_fd_sc_hd__dfrbp_2 merge840 (.CLK(clknet_4_7_0_clk),
    .D(net147),
    .RESET_B(net158),
    .Q(net620),
    .Q_N(net619));
 sky130_fd_sc_hd__and2_0 merge841 (.A(net531),
    .B(net556),
    .X(net621));
 sky130_fd_sc_hd__dfrtn_1 merge842 (.CLK_N(clknet_4_8_0_clk),
    .D(net436),
    .RESET_B(net566),
    .Q(net622));
 sky130_fd_sc_hd__dfrtp_1 merge843 (.CLK(clknet_4_5_0_clk),
    .D(net51),
    .Q(net59));
 sky130_fd_sc_hd__dfrtp_1 merge844 (.CLK(clknet_4_11_0_clk),
    .RESET_B(net513),
    .Q(net519));
 sky130_fd_sc_hd__and2_0 merge845 (.A(net454),
    .B(net614),
    .X(net625));
 sky130_fd_sc_hd__dfrtp_1 merge846 (.CLK(clknet_4_5_0_clk),
    .D(net45),
    .Q(net50));
 sky130_fd_sc_hd__and2_0 merge847 (.A(net225),
    .B(net120),
    .X(net627));
 sky130_fd_sc_hd__and2_0 merge848 (.A(net220),
    .B(net564),
    .X(net628));
 sky130_fd_sc_hd__dfsbp_1 merge849 (.CLK(clknet_4_0_0_clk),
    .D(net117),
    .SET_B(net103),
    .Q(net630),
    .Q_N(net629));
 sky130_fd_sc_hd__dfsbp_1 merge850 (.CLK(clknet_4_10_0_clk),
    .D(net444),
    .SET_B(net608),
    .Q(net632),
    .Q_N(net631));
 sky130_fd_sc_hd__dfstp_2 merge851 (.CLK(clknet_4_2_0_clk),
    .D(net420),
    .SET_B(net224),
    .Q(net633));
 sky130_fd_sc_hd__and2_0 merge852 (.A(net537),
    .B(net539),
    .X(net634));
 sky130_fd_sc_hd__dfstp_1 merge853 (.CLK(clknet_4_8_0_clk),
    .D(net574),
    .SET_B(net606),
    .Q(net635));
 sky130_fd_sc_hd__and2_0 merge854 (.A(net634),
    .B(net553),
    .X(net636));
 sky130_fd_sc_hd__and2_0 merge855 (.A(net551),
    .B(net548),
    .X(net637));
 sky130_fd_sc_hd__dfstp_1 merge856 (.CLK(clknet_4_10_0_clk),
    .D(net507),
    .SET_B(net582),
    .Q(net877));
 sky130_fd_sc_hd__dlrbn_1 merge857 (.D(net592),
    .GATE_N(clknet_4_10_0_clk),
    .RESET_B(net637),
    .Q(net638),
    .Q_N(net879));
 sky130_fd_sc_hd__dlrbn_1 merge858 (.D(net367),
    .GATE_N(clknet_4_11_0_clk),
    .RESET_B(net521),
    .Q(net640),
    .Q_N(net639));
 sky130_fd_sc_hd__dlrbp_1 merge859 (.GATE(clknet_4_14_0_clk),
    .RESET_B(net483),
    .Q(net642),
    .Q_N(net641));
 sky130_fd_sc_hd__dlrbp_1 merge860 (.D(net190),
    .GATE(clknet_4_2_0_clk),
    .RESET_B(net341),
    .Q(net644),
    .Q_N(net643));
 sky130_fd_sc_hd__dlrtn_1 merge861 (.GATE_N(clknet_4_3_0_clk),
    .RESET_B(net210),
    .Q(net211));
 sky130_fd_sc_hd__dlrtn_2 merge862 (.D(net580),
    .GATE_N(clknet_4_2_0_clk),
    .RESET_B(net194),
    .Q(net928));
 sky130_fd_sc_hd__dlrtn_2 merge863 (.D(net297),
    .GATE_N(clknet_4_9_0_clk),
    .RESET_B(net583),
    .Q(net645));
 sky130_fd_sc_hd__dlrtp_2 merge864 (.D(net320),
    .GATE(clknet_4_8_0_clk),
    .RESET_B(net317),
    .Q(net646));
 sky130_fd_sc_hd__dlrtp_2 merge865 (.D(net185),
    .GATE(clknet_4_4_0_clk),
    .RESET_B(net180),
    .Q(net647));
 sky130_fd_sc_hd__dlrtp_1 merge866 (.D(net636),
    .GATE(clknet_4_10_0_clk),
    .RESET_B(net594),
    .Q(net878));
 sky130_fd_sc_hd__edfxbp_1 merge867 (.CLK(clknet_4_2_0_clk),
    .D(net213),
    .DE(net230),
    .Q(net649),
    .Q_N(net648));
 sky130_fd_sc_hd__edfxtp_1 merge868 (.CLK(clknet_4_2_0_clk),
    .D(net227),
    .DE(net200),
    .Q(net919));
 sky130_fd_sc_hd__sdlclkp_1 merge869 (.CLK(clknet_4_15_0_clk),
    .GATE(net371),
    .GCLK(net434));
 sky130_fd_sc_hd__sdlclkp_2 merge870 (.CLK(clknet_4_1_0_clk),
    .GATE(net311),
    .SCE(net600),
    .GCLK(net938));
 sky130_fd_sc_hd__sdlclkp_4 merge871 (.CLK(clknet_4_0_0_clk),
    .GATE(net326),
    .SCE(net603),
    .GCLK(net651));
 sky130_fd_sc_hd__and2_0 merge872 (.A(net621),
    .B(net598),
    .X(net652));
 sky130_fd_sc_hd__dfrbp_2 merge873 (.CLK(clknet_4_15_0_clk),
    .D(net467),
    .RESET_B(net511),
    .Q(net654),
    .Q_N(net653));
 sky130_fd_sc_hd__dfrbp_1 merge874 (.CLK(clknet_4_10_0_clk),
    .D(net451),
    .RESET_B(net593),
    .Q(net655),
    .Q_N(net875));
 sky130_fd_sc_hd__dfrtn_1 merge875 (.CLK_N(clknet_4_10_0_clk),
    .D(net584),
    .RESET_B(net540),
    .Q(net656));
 sky130_fd_sc_hd__dfrtp_2 merge876 (.CLK(clknet_4_10_0_clk),
    .D(net538),
    .RESET_B(net529),
    .Q(net657));
 sky130_fd_sc_hd__dfrtp_4 merge877 (.CLK(clknet_4_8_0_clk),
    .D(net397),
    .RESET_B(net625),
    .Q(net658));
 sky130_fd_sc_hd__dfrtp_4 merge878 (.CLK(clknet_4_10_0_clk),
    .D(net510),
    .RESET_B(net223),
    .Q(net915));
 sky130_fd_sc_hd__dfsbp_1 merge879 (.CLK(clknet_4_14_0_clk),
    .D(net459),
    .SET_B(net489),
    .Q(net660),
    .Q_N(net659));
 sky130_fd_sc_hd__dfsbp_1 merge880 (.CLK(clknet_4_2_0_clk),
    .D(net215),
    .SET_B(net212),
    .Q(net662),
    .Q_N(net661));
 sky130_fd_sc_hd__dfstp_2 merge881 (.CLK(clknet_4_15_0_clk),
    .D(net468),
    .SET_B(net652),
    .Q(net663));
 sky130_fd_sc_hd__dfstp_4 merge882 (.CLK(clknet_4_2_0_clk),
    .D(net169),
    .SET_B(net628),
    .Q(net901));
 sky130_fd_sc_hd__dfstp_2 merge883 (.CLK(clknet_4_15_0_clk),
    .D(net476),
    .SET_B(net469),
    .Q(net664));
 sky130_fd_sc_hd__dlrbn_2 merge884 (.D(net577),
    .GATE_N(clknet_4_0_0_clk),
    .RESET_B(net627),
    .Q(net920),
    .Q_N(net940));
 sky130_fd_sc_hd__dlrbn_2 merge885 (.D(net599),
    .GATE_N(clknet_4_6_0_clk),
    .RESET_B(net565),
    .Q(net911),
    .Q_N(net665));
 sky130_fd_sc_hd__dlrbp_1 merge886 (.D(net526),
    .GATE(clknet_4_11_0_clk),
    .RESET_B(net481),
    .Q(net667),
    .Q_N(net666));
 sky130_fd_sc_hd__dfxbp_2 s887 (.CLK(clknet_4_5_0_clk),
    .D(net55),
    .Q(net669),
    .Q_N(net668));
 sky130_fd_sc_hd__dfxbp_2 s888 (.CLK(clknet_4_4_0_clk),
    .D(net56),
    .Q(net883),
    .Q_N(net670));
 sky130_fd_sc_hd__dfxtp_4 s889 (.CLK(clknet_4_5_0_clk),
    .D(net57),
    .Q(net671));
 sky130_fd_sc_hd__dfxtp_4 s890 (.CLK(clknet_4_5_0_clk),
    .D(net58),
    .Q(net672));
 sky130_fd_sc_hd__dfxtp_4 s891 (.CLK(clknet_4_4_0_clk),
    .D(net64),
    .Q(net912));
 sky130_fd_sc_hd__dlclkp_1 s892 (.CLK(clknet_4_4_0_clk),
    .GATE(net65),
    .GCLK(net673));
 sky130_fd_sc_hd__dlclkp_2 s893 (.CLK(clknet_4_1_0_clk),
    .GATE(net69),
    .GCLK(net674));
 sky130_fd_sc_hd__dlclkp_4 s894 (.CLK(clknet_4_5_0_clk),
    .GATE(net80),
    .GCLK(net675));
 sky130_fd_sc_hd__dlxbn_1 s895 (.D(net82),
    .GATE_N(clknet_4_0_0_clk),
    .Q(net903),
    .Q_N(net676));
 sky130_fd_sc_hd__dlxbn_1 s896 (.D(net89),
    .GATE_N(clknet_4_1_0_clk),
    .Q(net678),
    .Q_N(net677));
 sky130_fd_sc_hd__dlxbp_1 s897 (.D(net92),
    .GATE(clknet_4_1_0_clk),
    .Q(net680),
    .Q_N(net679));
 sky130_fd_sc_hd__dlxtn_2 s898 (.D(net93),
    .GATE_N(clknet_4_1_0_clk),
    .Q(net681));
 sky130_fd_sc_hd__dlxtn_1 s899 (.D(net105),
    .GATE_N(clknet_4_0_0_clk),
    .Q(net682));
 sky130_fd_sc_hd__dlxtn_4 s900 (.D(net121),
    .GATE_N(clknet_4_0_0_clk),
    .Q(net683));
 sky130_fd_sc_hd__dlxtp_1 s901 (.D(net139),
    .GATE(clknet_4_7_0_clk),
    .Q(net684));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s902 (.D(net142),
    .SLEEP_B(clknet_4_7_0_clk),
    .Q(net685));
 sky130_fd_sc_hd__dfxbp_2 s903 (.CLK(clknet_4_7_0_clk),
    .D(net145),
    .Q(net687),
    .Q_N(net686));
 sky130_fd_sc_hd__dfxbp_2 s904 (.CLK(clknet_4_13_0_clk),
    .D(net146),
    .Q(net689),
    .Q_N(net688));
 sky130_fd_sc_hd__dfxtp_1 s905 (.CLK(clknet_4_7_0_clk),
    .D(net149),
    .Q(net690));
 sky130_fd_sc_hd__dfxtp_1 s906 (.CLK(clknet_4_7_0_clk),
    .D(net152),
    .Q(net691));
 sky130_fd_sc_hd__dfxtp_4 s907 (.CLK(clknet_4_7_0_clk),
    .D(net153),
    .Q(net692));
 sky130_fd_sc_hd__dlclkp_1 s908 (.CLK(clknet_4_4_0_clk),
    .GATE(net156),
    .GCLK(net693));
 sky130_fd_sc_hd__dlclkp_2 s909 (.CLK(clknet_4_6_0_clk),
    .GATE(net159),
    .GCLK(net694));
 sky130_fd_sc_hd__dlclkp_4 s910 (.CLK(clknet_4_7_0_clk),
    .GATE(net160),
    .GCLK(net695));
 sky130_fd_sc_hd__dlxbn_2 s911 (.D(net162),
    .GATE_N(clknet_4_6_0_clk),
    .Q(net697),
    .Q_N(net696));
 sky130_fd_sc_hd__dlxbn_2 s912 (.D(net163),
    .GATE_N(clknet_4_6_0_clk),
    .Q(net873),
    .Q_N(net698));
 sky130_fd_sc_hd__dlxbp_1 s913 (.D(net164),
    .GATE(clknet_4_9_0_clk),
    .Q(net700),
    .Q_N(net699));
 sky130_fd_sc_hd__dlxtn_2 s914 (.D(net170),
    .GATE_N(clknet_4_6_0_clk),
    .Q(net701));
 sky130_fd_sc_hd__dlxtn_1 s915 (.D(net172),
    .GATE_N(clknet_4_6_0_clk),
    .Q(net702));
 sky130_fd_sc_hd__dlxtn_2 s916 (.D(net176),
    .GATE_N(clknet_4_1_0_clk),
    .Q(net703));
 sky130_fd_sc_hd__dlxtp_1 s917 (.D(net183),
    .GATE(clknet_4_3_0_clk),
    .Q(net704));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s918 (.D(net189),
    .SLEEP_B(clknet_4_3_0_clk),
    .Q(net705));
 sky130_fd_sc_hd__dfxbp_1 s919 (.CLK(clknet_4_3_0_clk),
    .D(net195),
    .Q(net707),
    .Q_N(net706));
 sky130_fd_sc_hd__dfxbp_2 s920 (.CLK(clknet_4_2_0_clk),
    .D(net203),
    .Q(net709),
    .Q_N(net708));
 sky130_fd_sc_hd__dfxtp_1 s921 (.CLK(clknet_4_0_0_clk),
    .D(net204),
    .Q(net921));
 sky130_fd_sc_hd__dfxtp_1 s922 (.CLK(clknet_4_3_0_clk),
    .D(net205),
    .Q(net710));
 sky130_fd_sc_hd__dfxtp_2 s923 (.CLK(clknet_4_0_0_clk),
    .D(net217),
    .Q(net711));
 sky130_fd_sc_hd__dlclkp_1 s924 (.CLK(clknet_4_13_0_clk),
    .GATE(net244),
    .GCLK(net712));
 sky130_fd_sc_hd__dlclkp_2 s925 (.CLK(clknet_4_13_0_clk),
    .GATE(net249),
    .GCLK(net713));
 sky130_fd_sc_hd__dlclkp_4 s926 (.CLK(clknet_4_13_0_clk),
    .GATE(net256),
    .GCLK(net714));
 sky130_fd_sc_hd__dlxbn_1 s927 (.D(net259),
    .GATE_N(clknet_4_13_0_clk),
    .Q(net716),
    .Q_N(net715));
 sky130_fd_sc_hd__dlxbn_1 s928 (.D(net262),
    .GATE_N(clknet_4_12_0_clk),
    .Q(net718),
    .Q_N(net717));
 sky130_fd_sc_hd__dlxbp_1 s929 (.D(net264),
    .GATE(clknet_4_6_0_clk),
    .Q(net720),
    .Q_N(net719));
 sky130_fd_sc_hd__dlxtn_2 s930 (.D(net266),
    .GATE_N(clknet_4_12_0_clk),
    .Q(net721));
 sky130_fd_sc_hd__dlxtn_1 s931 (.D(net267),
    .GATE_N(clknet_4_12_0_clk),
    .Q(net722));
 sky130_fd_sc_hd__dlxtn_2 s932 (.D(net268),
    .GATE_N(clknet_4_12_0_clk),
    .Q(net723));
 sky130_fd_sc_hd__dlxtp_1 s933 (.D(net270),
    .GATE(clknet_4_6_0_clk),
    .Q(net724));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s934 (.D(net272),
    .SLEEP_B(clknet_4_12_0_clk),
    .Q(net725));
 sky130_fd_sc_hd__dfxbp_1 s935 (.CLK(clknet_4_12_0_clk),
    .D(net274),
    .Q(net727),
    .Q_N(net726));
 sky130_fd_sc_hd__dfxbp_1 s936 (.CLK(clknet_4_12_0_clk),
    .D(net275),
    .Q(net729),
    .Q_N(net728));
 sky130_fd_sc_hd__dfxtp_2 s937 (.CLK(clknet_4_12_0_clk),
    .D(net279),
    .Q(net730));
 sky130_fd_sc_hd__dfxtp_4 s938 (.CLK(clknet_4_9_0_clk),
    .D(net280),
    .Q(net731));
 sky130_fd_sc_hd__dfxtp_1 s939 (.CLK(clknet_4_9_0_clk),
    .D(net286),
    .Q(net732));
 sky130_fd_sc_hd__dlclkp_1 s940 (.CLK(clknet_4_9_0_clk),
    .GATE(net289),
    .GCLK(net733));
 sky130_fd_sc_hd__dlclkp_2 s941 (.CLK(clknet_4_3_0_clk),
    .GATE(net292),
    .GCLK(net734));
 sky130_fd_sc_hd__dlclkp_4 s942 (.CLK(clknet_4_3_0_clk),
    .GATE(net294),
    .GCLK(net735));
 sky130_fd_sc_hd__dlxbn_2 s943 (.D(net299),
    .GATE_N(clknet_4_9_0_clk),
    .Q(net737),
    .Q_N(net736));
 sky130_fd_sc_hd__dlxbn_2 s944 (.D(net301),
    .GATE_N(clknet_4_3_0_clk),
    .Q(net889),
    .Q_N(net738));
 sky130_fd_sc_hd__dlxbp_1 s945 (.D(net303),
    .GATE(clknet_4_9_0_clk),
    .Q(net740),
    .Q_N(net739));
 sky130_fd_sc_hd__dlxtn_4 s946 (.D(net305),
    .GATE_N(clknet_4_3_0_clk),
    .Q(net741));
 sky130_fd_sc_hd__dlxtn_1 s947 (.D(net313),
    .GATE_N(clknet_4_8_0_clk),
    .Q(net742));
 sky130_fd_sc_hd__dlxtn_2 s948 (.D(net315),
    .GATE_N(clknet_4_2_0_clk),
    .Q(net743));
 sky130_fd_sc_hd__dlxtp_1 s949 (.D(net319),
    .GATE(clknet_4_3_0_clk),
    .Q(net913));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s950 (.D(net323),
    .SLEEP_B(clknet_4_2_0_clk),
    .Q(net744));
 sky130_fd_sc_hd__dfxbp_1 s951 (.CLK(clknet_4_8_0_clk),
    .D(net338),
    .Q(net746),
    .Q_N(net745));
 sky130_fd_sc_hd__dfxbp_1 s952 (.CLK(clknet_4_13_0_clk),
    .D(net342),
    .Q(net748),
    .Q_N(net747));
 sky130_fd_sc_hd__dfxtp_4 s953 (.CLK(clknet_4_15_0_clk),
    .D(net365),
    .Q(net891));
 sky130_fd_sc_hd__dfxtp_1 s954 (.CLK(clknet_4_12_0_clk),
    .D(net376),
    .Q(net749));
 sky130_fd_sc_hd__dfxtp_2 s955 (.CLK(clknet_4_11_0_clk),
    .D(net389),
    .Q(net750));
 sky130_fd_sc_hd__dlclkp_1 s956 (.CLK(clknet_4_9_0_clk),
    .GATE(net391),
    .GCLK(net751));
 sky130_fd_sc_hd__dlclkp_2 s957 (.CLK(clknet_4_11_0_clk),
    .GATE(net398),
    .GCLK(net752));
 sky130_fd_sc_hd__dlclkp_4 s958 (.CLK(clknet_4_11_0_clk),
    .GATE(net404),
    .GCLK(net753));
 sky130_fd_sc_hd__dlxbn_1 s959 (.D(net406),
    .GATE_N(clknet_4_10_0_clk),
    .Q(net876),
    .Q_N(net754));
 sky130_fd_sc_hd__dlxbn_1 s960 (.D(net408),
    .GATE_N(clknet_4_9_0_clk),
    .Q(net756),
    .Q_N(net755));
 sky130_fd_sc_hd__dlxbp_1 s961 (.D(net421),
    .GATE(clknet_4_8_0_clk),
    .Q(net758),
    .Q_N(net757));
 sky130_fd_sc_hd__dlxtn_2 s962 (.D(net425),
    .GATE_N(clknet_4_8_0_clk),
    .Q(net759));
 sky130_fd_sc_hd__dlxtn_1 s963 (.D(net443),
    .GATE_N(clknet_4_8_0_clk),
    .Q(net760));
 sky130_fd_sc_hd__dlxtn_2 s964 (.D(net463),
    .GATE_N(clknet_4_15_0_clk),
    .Q(net761));
 sky130_fd_sc_hd__dlxtp_1 s965 (.D(net470),
    .GATE(clknet_4_15_0_clk),
    .Q(net762));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s966 (.D(net473),
    .SLEEP_B(clknet_4_15_0_clk),
    .Q(net763));
 sky130_fd_sc_hd__dfxbp_1 s967 (.CLK(clknet_4_14_0_clk),
    .D(net478),
    .Q(net765),
    .Q_N(net764));
 sky130_fd_sc_hd__dfxbp_1 s968 (.CLK(clknet_4_14_0_clk),
    .D(net482),
    .Q(net767),
    .Q_N(net766));
 sky130_fd_sc_hd__dfxtp_2 s969 (.CLK(clknet_4_14_0_clk),
    .D(net485),
    .Q(net768));
 sky130_fd_sc_hd__dfxtp_1 s970 (.CLK(clknet_4_14_0_clk),
    .D(net497),
    .Q(net769));
 sky130_fd_sc_hd__dfxtp_1 s971 (.CLK(clknet_4_11_0_clk),
    .D(net499),
    .Q(net770));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Right_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Right_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Right_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Right_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Right_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Right_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Right_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Right_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Right_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Right_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Right_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Right_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Right_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Right_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Right_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Right_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Right_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Right_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Right_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Right_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Right_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_161 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_162 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_163 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_164 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_165 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_166 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_167 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_168 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_169 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_170 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_171 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_172 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_173 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_174 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_175 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_176 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_177 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_178 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_179 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_180 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_181 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_182 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Left_183 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Left_184 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Left_185 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Left_186 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Left_187 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Left_188 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Left_189 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Left_190 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Left_191 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Left_192 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Left_193 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Left_194 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Left_195 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Left_196 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Left_197 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Left_198 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Left_199 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Left_200 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Left_201 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Left_202 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Left_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1347 ();
 sky130_fd_sc_hd__buf_4 input1 (.A(in0),
    .X(net484));
 sky130_fd_sc_hd__buf_4 input2 (.A(in1),
    .X(net771));
 sky130_fd_sc_hd__buf_2 input3 (.A(in10),
    .X(net772));
 sky130_fd_sc_hd__dlymetal6s2s_1 input4 (.A(in11),
    .X(net773));
 sky130_fd_sc_hd__buf_1 input5 (.A(in12),
    .X(net774));
 sky130_fd_sc_hd__buf_4 input6 (.A(in13),
    .X(net775));
 sky130_fd_sc_hd__buf_6 input7 (.A(in14),
    .X(net776));
 sky130_fd_sc_hd__buf_1 input8 (.A(in15),
    .X(net777));
 sky130_fd_sc_hd__clkbuf_4 input9 (.A(in16),
    .X(net778));
 sky130_fd_sc_hd__clkbuf_4 input10 (.A(in17),
    .X(net779));
 sky130_fd_sc_hd__buf_2 input11 (.A(in18),
    .X(net780));
 sky130_fd_sc_hd__buf_1 input12 (.A(in19),
    .X(net781));
 sky130_fd_sc_hd__dlymetal6s2s_1 input13 (.A(in2),
    .X(net782));
 sky130_fd_sc_hd__buf_1 input14 (.A(in20),
    .X(net783));
 sky130_fd_sc_hd__dlymetal6s2s_1 input15 (.A(in21),
    .X(net784));
 sky130_fd_sc_hd__buf_4 input16 (.A(in22),
    .X(net785));
 sky130_fd_sc_hd__buf_1 input17 (.A(in23),
    .X(net786));
 sky130_fd_sc_hd__buf_4 input18 (.A(in24),
    .X(net787));
 sky130_fd_sc_hd__clkbuf_2 input19 (.A(in25),
    .X(net788));
 sky130_fd_sc_hd__clkbuf_2 input20 (.A(in26),
    .X(net789));
 sky130_fd_sc_hd__buf_2 input21 (.A(in27),
    .X(net790));
 sky130_fd_sc_hd__clkbuf_2 input22 (.A(in28),
    .X(net791));
 sky130_fd_sc_hd__buf_2 input23 (.A(in29),
    .X(net792));
 sky130_fd_sc_hd__clkbuf_4 input24 (.A(in3),
    .X(net793));
 sky130_fd_sc_hd__buf_2 input25 (.A(in30),
    .X(net794));
 sky130_fd_sc_hd__buf_4 input26 (.A(in31),
    .X(net795));
 sky130_fd_sc_hd__buf_4 input27 (.A(in32),
    .X(net796));
 sky130_fd_sc_hd__clkbuf_4 input28 (.A(in33),
    .X(net797));
 sky130_fd_sc_hd__buf_4 input29 (.A(in34),
    .X(net798));
 sky130_fd_sc_hd__buf_2 input30 (.A(in35),
    .X(net799));
 sky130_fd_sc_hd__clkbuf_4 input31 (.A(in36),
    .X(net800));
 sky130_fd_sc_hd__buf_2 input32 (.A(in37),
    .X(net801));
 sky130_fd_sc_hd__clkbuf_2 input33 (.A(in38),
    .X(net802));
 sky130_fd_sc_hd__buf_1 input34 (.A(in39),
    .X(net803));
 sky130_fd_sc_hd__clkbuf_8 input35 (.A(in4),
    .X(net804));
 sky130_fd_sc_hd__buf_4 input36 (.A(in40),
    .X(net805));
 sky130_fd_sc_hd__clkbuf_4 input37 (.A(in41),
    .X(net806));
 sky130_fd_sc_hd__buf_2 input38 (.A(in42),
    .X(net807));
 sky130_fd_sc_hd__buf_4 input39 (.A(in43),
    .X(net808));
 sky130_fd_sc_hd__clkbuf_4 input40 (.A(in44),
    .X(net809));
 sky130_fd_sc_hd__buf_1 input41 (.A(in45),
    .X(net810));
 sky130_fd_sc_hd__clkbuf_2 input42 (.A(in46),
    .X(net811));
 sky130_fd_sc_hd__dlymetal6s2s_1 input43 (.A(in47),
    .X(net812));
 sky130_fd_sc_hd__clkbuf_2 input44 (.A(in48),
    .X(net813));
 sky130_fd_sc_hd__clkbuf_4 input45 (.A(in49),
    .X(net814));
 sky130_fd_sc_hd__buf_12 input46 (.A(in5),
    .X(net815));
 sky130_fd_sc_hd__clkbuf_2 input47 (.A(in50),
    .X(net816));
 sky130_fd_sc_hd__clkbuf_4 input48 (.A(in51),
    .X(net817));
 sky130_fd_sc_hd__buf_2 input49 (.A(in52),
    .X(net818));
 sky130_fd_sc_hd__clkbuf_2 input50 (.A(in53),
    .X(net819));
 sky130_fd_sc_hd__clkbuf_2 input51 (.A(in54),
    .X(net820));
 sky130_fd_sc_hd__clkbuf_4 input52 (.A(in55),
    .X(net821));
 sky130_fd_sc_hd__clkbuf_4 input53 (.A(in56),
    .X(net822));
 sky130_fd_sc_hd__buf_1 input54 (.A(in57),
    .X(net823));
 sky130_fd_sc_hd__buf_1 input55 (.A(in58),
    .X(net824));
 sky130_fd_sc_hd__buf_4 input56 (.A(in59),
    .X(net825));
 sky130_fd_sc_hd__clkbuf_4 input57 (.A(in6),
    .X(net826));
 sky130_fd_sc_hd__clkbuf_4 input58 (.A(in60),
    .X(net827));
 sky130_fd_sc_hd__buf_4 input59 (.A(in61),
    .X(net828));
 sky130_fd_sc_hd__clkbuf_2 input60 (.A(in62),
    .X(net829));
 sky130_fd_sc_hd__clkbuf_2 input61 (.A(in63),
    .X(net830));
 sky130_fd_sc_hd__clkbuf_2 input62 (.A(in64),
    .X(net831));
 sky130_fd_sc_hd__clkbuf_2 input63 (.A(in65),
    .X(net832));
 sky130_fd_sc_hd__clkbuf_2 input64 (.A(in66),
    .X(net833));
 sky130_fd_sc_hd__buf_1 input65 (.A(in67),
    .X(net834));
 sky130_fd_sc_hd__clkbuf_1 input66 (.A(in68),
    .X(net835));
 sky130_fd_sc_hd__buf_1 input67 (.A(in69),
    .X(net836));
 sky130_fd_sc_hd__buf_4 input68 (.A(in7),
    .X(net837));
 sky130_fd_sc_hd__clkbuf_4 input69 (.A(in70),
    .X(net838));
 sky130_fd_sc_hd__buf_1 input70 (.A(in71),
    .X(net839));
 sky130_fd_sc_hd__buf_2 input71 (.A(in72),
    .X(net840));
 sky130_fd_sc_hd__clkbuf_4 input72 (.A(in73),
    .X(net841));
 sky130_fd_sc_hd__clkbuf_2 input73 (.A(in74),
    .X(net842));
 sky130_fd_sc_hd__buf_1 input74 (.A(in75),
    .X(net843));
 sky130_fd_sc_hd__buf_1 input75 (.A(in76),
    .X(net844));
 sky130_fd_sc_hd__buf_1 input76 (.A(in77),
    .X(net845));
 sky130_fd_sc_hd__buf_1 input77 (.A(in78),
    .X(net846));
 sky130_fd_sc_hd__buf_1 input78 (.A(in79),
    .X(net847));
 sky130_fd_sc_hd__buf_1 input79 (.A(in8),
    .X(net848));
 sky130_fd_sc_hd__buf_1 input80 (.A(in80),
    .X(net849));
 sky130_fd_sc_hd__clkbuf_1 input81 (.A(in81),
    .X(net850));
 sky130_fd_sc_hd__buf_1 input82 (.A(in82),
    .X(net851));
 sky130_fd_sc_hd__buf_1 input83 (.A(in83),
    .X(net852));
 sky130_fd_sc_hd__buf_1 input84 (.A(in84),
    .X(net853));
 sky130_fd_sc_hd__buf_1 input85 (.A(in85),
    .X(net854));
 sky130_fd_sc_hd__buf_1 input86 (.A(in86),
    .X(net855));
 sky130_fd_sc_hd__buf_1 input87 (.A(in87),
    .X(net856));
 sky130_fd_sc_hd__buf_2 input88 (.A(in88),
    .X(net857));
 sky130_fd_sc_hd__clkbuf_2 input89 (.A(in89),
    .X(net858));
 sky130_fd_sc_hd__dlymetal6s2s_1 input90 (.A(in9),
    .X(net859));
 sky130_fd_sc_hd__buf_1 input91 (.A(in90),
    .X(net860));
 sky130_fd_sc_hd__buf_2 input92 (.A(in91),
    .X(net861));
 sky130_fd_sc_hd__dlymetal6s2s_1 input93 (.A(in92),
    .X(net862));
 sky130_fd_sc_hd__clkbuf_2 input94 (.A(in93),
    .X(net863));
 sky130_fd_sc_hd__buf_1 input95 (.A(in94),
    .X(net864));
 sky130_fd_sc_hd__clkbuf_2 input96 (.A(in95),
    .X(net865));
 sky130_fd_sc_hd__buf_1 input97 (.A(in96),
    .X(net866));
 sky130_fd_sc_hd__buf_2 input98 (.A(in97),
    .X(net867));
 sky130_fd_sc_hd__clkbuf_2 input99 (.A(in98),
    .X(net868));
 sky130_fd_sc_hd__buf_1 input100 (.A(in99),
    .X(net869));
 sky130_fd_sc_hd__clkbuf_1 output101 (.A(net870),
    .X(out0));
 sky130_fd_sc_hd__buf_2 output102 (.A(net871),
    .X(out1));
 sky130_fd_sc_hd__buf_2 output103 (.A(net976),
    .X(out10));
 sky130_fd_sc_hd__buf_2 output104 (.A(net873),
    .X(out11));
 sky130_fd_sc_hd__buf_2 output105 (.A(net874),
    .X(out13));
 sky130_fd_sc_hd__buf_2 output106 (.A(net875),
    .X(out14));
 sky130_fd_sc_hd__buf_2 output107 (.A(net876),
    .X(out15));
 sky130_fd_sc_hd__buf_2 output108 (.A(net877),
    .X(out16));
 sky130_fd_sc_hd__buf_2 output109 (.A(net878),
    .X(out17));
 sky130_fd_sc_hd__buf_2 output110 (.A(net879),
    .X(out18));
 sky130_fd_sc_hd__buf_2 output111 (.A(net880),
    .X(out21));
 sky130_fd_sc_hd__buf_2 output112 (.A(net881),
    .X(out22));
 sky130_fd_sc_hd__clkbuf_1 output113 (.A(net882),
    .X(out23));
 sky130_fd_sc_hd__buf_2 output114 (.A(net883),
    .X(out24));
 sky130_fd_sc_hd__clkbuf_1 output115 (.A(net884),
    .X(out25));
 sky130_fd_sc_hd__clkbuf_4 output116 (.A(net970),
    .X(out26));
 sky130_fd_sc_hd__clkbuf_1 output117 (.A(net886),
    .X(out28));
 sky130_fd_sc_hd__clkbuf_1 output118 (.A(clknet_1_0__leaf_net887),
    .X(out29));
 sky130_fd_sc_hd__buf_2 output119 (.A(net888),
    .X(out31));
 sky130_fd_sc_hd__buf_2 output120 (.A(net889),
    .X(out32));
 sky130_fd_sc_hd__clkbuf_1 output121 (.A(clknet_1_0__leaf_net890),
    .X(out34));
 sky130_fd_sc_hd__buf_2 output122 (.A(net891),
    .X(out35));
 sky130_fd_sc_hd__buf_2 output123 (.A(net892),
    .X(out36));
 sky130_fd_sc_hd__clkbuf_1 output124 (.A(clknet_1_1__leaf_net893),
    .X(out37));
 sky130_fd_sc_hd__clkbuf_1 output125 (.A(clknet_1_0__leaf_net894),
    .X(out39));
 sky130_fd_sc_hd__clkbuf_1 output126 (.A(clknet_1_1__leaf_net895),
    .X(out40));
 sky130_fd_sc_hd__buf_2 output127 (.A(net896),
    .X(out42));
 sky130_fd_sc_hd__buf_2 output128 (.A(net897),
    .X(out43));
 sky130_fd_sc_hd__clkbuf_1 output129 (.A(clknet_1_1__leaf_net898),
    .X(out44));
 sky130_fd_sc_hd__clkbuf_1 output130 (.A(net899),
    .X(out45));
 sky130_fd_sc_hd__clkbuf_1 output131 (.A(clknet_1_0__leaf_net900),
    .X(out46));
 sky130_fd_sc_hd__buf_2 output132 (.A(net901),
    .X(out47));
 sky130_fd_sc_hd__buf_2 output133 (.A(net902),
    .X(out48));
 sky130_fd_sc_hd__buf_2 output134 (.A(net903),
    .X(out49));
 sky130_fd_sc_hd__clkbuf_1 output135 (.A(clknet_1_1__leaf_net904),
    .X(out5));
 sky130_fd_sc_hd__clkbuf_1 output136 (.A(clknet_1_1__leaf_net905),
    .X(out51));
 sky130_fd_sc_hd__buf_2 output137 (.A(net906),
    .X(out53));
 sky130_fd_sc_hd__buf_2 output138 (.A(net907),
    .X(out54));
 sky130_fd_sc_hd__clkbuf_1 output139 (.A(clknet_1_0__leaf_net908),
    .X(out55));
 sky130_fd_sc_hd__buf_2 output140 (.A(net909),
    .X(out56));
 sky130_fd_sc_hd__buf_2 output141 (.A(net910),
    .X(out57));
 sky130_fd_sc_hd__buf_2 output142 (.A(net911),
    .X(out58));
 sky130_fd_sc_hd__buf_2 output143 (.A(net912),
    .X(out59));
 sky130_fd_sc_hd__buf_2 output144 (.A(net913),
    .X(out6));
 sky130_fd_sc_hd__buf_2 output145 (.A(net914),
    .X(out60));
 sky130_fd_sc_hd__buf_2 output146 (.A(net915),
    .X(out61));
 sky130_fd_sc_hd__clkbuf_1 output147 (.A(clknet_1_0__leaf_net916),
    .X(out64));
 sky130_fd_sc_hd__buf_2 output148 (.A(net917),
    .X(out65));
 sky130_fd_sc_hd__buf_2 output149 (.A(net918),
    .X(out66));
 sky130_fd_sc_hd__buf_2 output150 (.A(net919),
    .X(out67));
 sky130_fd_sc_hd__buf_2 output151 (.A(net920),
    .X(out68));
 sky130_fd_sc_hd__buf_2 output152 (.A(net989),
    .X(out69));
 sky130_fd_sc_hd__clkbuf_1 output153 (.A(clknet_1_0__leaf_net922),
    .X(out70));
 sky130_fd_sc_hd__clkbuf_1 output154 (.A(clknet_1_0__leaf_net923),
    .X(out71));
 sky130_fd_sc_hd__buf_2 output155 (.A(net924),
    .X(out72));
 sky130_fd_sc_hd__buf_2 output156 (.A(net925),
    .X(out73));
 sky130_fd_sc_hd__buf_2 output157 (.A(net926),
    .X(out75));
 sky130_fd_sc_hd__buf_2 output158 (.A(net927),
    .X(out76));
 sky130_fd_sc_hd__buf_2 output159 (.A(net928),
    .X(out78));
 sky130_fd_sc_hd__buf_2 output160 (.A(net929),
    .X(out79));
 sky130_fd_sc_hd__clkbuf_1 output161 (.A(net930),
    .X(out8));
 sky130_fd_sc_hd__buf_2 output162 (.A(net931),
    .X(out80));
 sky130_fd_sc_hd__clkbuf_4 output163 (.A(net932),
    .X(out81));
 sky130_fd_sc_hd__buf_2 output164 (.A(net933),
    .X(out82));
 sky130_fd_sc_hd__buf_2 output165 (.A(net934),
    .X(out83));
 sky130_fd_sc_hd__clkbuf_1 output166 (.A(clknet_1_1__leaf_net935),
    .X(out84));
 sky130_fd_sc_hd__clkbuf_1 output167 (.A(clknet_1_1__leaf_net936),
    .X(out85));
 sky130_fd_sc_hd__buf_2 output168 (.A(net937),
    .X(out88));
 sky130_fd_sc_hd__clkbuf_1 output169 (.A(clknet_1_1__leaf_net938),
    .X(out89));
 sky130_fd_sc_hd__clkbuf_1 output170 (.A(clknet_1_1__leaf_net939),
    .X(out9));
 sky130_fd_sc_hd__buf_2 output171 (.A(net940),
    .X(out90));
 sky130_fd_sc_hd__buf_2 output172 (.A(net941),
    .X(out91));
 sky130_fd_sc_hd__buf_2 output173 (.A(net942),
    .X(out93));
 sky130_fd_sc_hd__buf_2 output174 (.A(net943),
    .X(out95));
 sky130_fd_sc_hd__buf_2 output175 (.A(net944),
    .X(out96));
 sky130_fd_sc_hd__buf_2 output176 (.A(net945),
    .X(out97));
 sky130_fd_sc_hd__buf_2 output177 (.A(net946),
    .X(out98));
 sky130_fd_sc_hd__buf_2 output178 (.A(net947),
    .X(out99));
 sky130_fd_sc_hd__clkbuf_4 fanout179 (.A(net148),
    .X(net948));
 sky130_fd_sc_hd__buf_2 fanout180 (.A(net950),
    .X(net949));
 sky130_fd_sc_hd__clkbuf_2 fanout181 (.A(net951),
    .X(net950));
 sky130_fd_sc_hd__clkbuf_4 fanout182 (.A(net952),
    .X(net951));
 sky130_fd_sc_hd__clkbuf_4 fanout183 (.A(net131),
    .X(net952));
 sky130_fd_sc_hd__buf_4 fanout184 (.A(net54),
    .X(net953));
 sky130_fd_sc_hd__buf_4 fanout185 (.A(net53),
    .X(net954));
 sky130_fd_sc_hd__clkbuf_4 fanout186 (.A(net956),
    .X(net955));
 sky130_fd_sc_hd__clkbuf_4 fanout187 (.A(net957),
    .X(net956));
 sky130_fd_sc_hd__clkbuf_4 fanout188 (.A(net47),
    .X(net957));
 sky130_fd_sc_hd__clkbuf_4 fanout189 (.A(net897),
    .X(net958));
 sky130_fd_sc_hd__clkbuf_4 fanout190 (.A(net234),
    .X(net959));
 sky130_fd_sc_hd__clkbuf_4 fanout191 (.A(net961),
    .X(net960));
 sky130_fd_sc_hd__clkbuf_4 fanout192 (.A(net130),
    .X(net961));
 sky130_fd_sc_hd__clkbuf_4 fanout193 (.A(net143),
    .X(net962));
 sky130_fd_sc_hd__buf_4 fanout194 (.A(net37),
    .X(net963));
 sky130_fd_sc_hd__buf_8 fanout195 (.A(net127),
    .X(net964));
 sky130_fd_sc_hd__buf_12 fanout196 (.A(net966),
    .X(net965));
 sky130_fd_sc_hd__buf_8 fanout197 (.A(net125),
    .X(net966));
 sky130_fd_sc_hd__clkbuf_4 fanout198 (.A(net61),
    .X(net967));
 sky130_fd_sc_hd__buf_4 fanout199 (.A(net39),
    .X(net968));
 sky130_fd_sc_hd__buf_4 fanout200 (.A(net885),
    .X(net969));
 sky130_fd_sc_hd__clkbuf_2 fanout201 (.A(net885),
    .X(net970));
 sky130_fd_sc_hd__buf_4 fanout202 (.A(net1038),
    .X(net971));
 sky130_fd_sc_hd__buf_8 fanout203 (.A(net34),
    .X(net972));
 sky130_fd_sc_hd__buf_12 fanout204 (.A(net33),
    .X(net973));
 sky130_fd_sc_hd__clkbuf_4 fanout205 (.A(net32),
    .X(net974));
 sky130_fd_sc_hd__buf_12 fanout206 (.A(net872),
    .X(net975));
 sky130_fd_sc_hd__buf_2 fanout207 (.A(net1036),
    .X(net976));
 sky130_fd_sc_hd__buf_4 fanout208 (.A(net30),
    .X(net977));
 sky130_fd_sc_hd__clkbuf_8 fanout209 (.A(net29),
    .X(net978));
 sky130_fd_sc_hd__clkbuf_2 fanout210 (.A(net29),
    .X(net979));
 sky130_fd_sc_hd__buf_4 fanout211 (.A(net27),
    .X(net980));
 sky130_fd_sc_hd__buf_12 fanout212 (.A(net23),
    .X(net981));
 sky130_fd_sc_hd__clkbuf_4 fanout213 (.A(net22),
    .X(net982));
 sky130_fd_sc_hd__clkbuf_4 fanout214 (.A(net984),
    .X(net983));
 sky130_fd_sc_hd__buf_8 fanout215 (.A(net985),
    .X(net984));
 sky130_fd_sc_hd__buf_8 fanout216 (.A(net986),
    .X(net985));
 sky130_fd_sc_hd__buf_8 fanout217 (.A(net21),
    .X(net986));
 sky130_fd_sc_hd__clkbuf_4 fanout218 (.A(net19),
    .X(net987));
 sky130_fd_sc_hd__buf_4 fanout219 (.A(net722),
    .X(net988));
 sky130_fd_sc_hd__clkbuf_4 fanout220 (.A(net921),
    .X(net989));
 sky130_fd_sc_hd__buf_2 max_cap221 (.A(net705),
    .X(net990));
 sky130_fd_sc_hd__clkbuf_4 fanout222 (.A(net702),
    .X(net991));
 sky130_fd_sc_hd__clkbuf_2 fanout223 (.A(net702),
    .X(net992));
 sky130_fd_sc_hd__buf_4 fanout224 (.A(net691),
    .X(net993));
 sky130_fd_sc_hd__clkbuf_4 fanout225 (.A(net995),
    .X(net994));
 sky130_fd_sc_hd__buf_4 fanout226 (.A(net690),
    .X(net995));
 sky130_fd_sc_hd__buf_4 fanout227 (.A(net689),
    .X(net996));
 sky130_fd_sc_hd__buf_4 fanout228 (.A(net20),
    .X(net997));
 sky130_fd_sc_hd__buf_8 fanout229 (.A(net18),
    .X(net998));
 sky130_fd_sc_hd__clkbuf_4 fanout230 (.A(net1),
    .X(net999));
 sky130_fd_sc_hd__clkbuf_4 fanout231 (.A(net865),
    .X(net1000));
 sky130_fd_sc_hd__buf_4 fanout232 (.A(net859),
    .X(net1001));
 sky130_fd_sc_hd__buf_4 fanout233 (.A(net1004),
    .X(net1002));
 sky130_fd_sc_hd__buf_4 fanout234 (.A(net1004),
    .X(net1003));
 sky130_fd_sc_hd__buf_2 fanout235 (.A(net777),
    .X(net1004));
 sky130_fd_sc_hd__clkbuf_8 fanout236 (.A(net848),
    .X(net1005));
 sky130_fd_sc_hd__buf_8 fanout237 (.A(net776),
    .X(net1006));
 sky130_fd_sc_hd__buf_8 fanout238 (.A(net826),
    .X(net1007));
 sky130_fd_sc_hd__clkbuf_2 fanout239 (.A(net826),
    .X(net1008));
 sky130_fd_sc_hd__buf_4 fanout240 (.A(net1010),
    .X(net1009));
 sky130_fd_sc_hd__buf_2 fanout241 (.A(net774),
    .X(net1010));
 sky130_fd_sc_hd__buf_12 fanout242 (.A(net1013),
    .X(net1011));
 sky130_fd_sc_hd__clkbuf_2 fanout243 (.A(net1013),
    .X(net1012));
 sky130_fd_sc_hd__buf_12 fanout244 (.A(net815),
    .X(net1013));
 sky130_fd_sc_hd__clkbuf_4 fanout245 (.A(net814),
    .X(net1014));
 sky130_fd_sc_hd__buf_4 fanout246 (.A(net810),
    .X(net1015));
 sky130_fd_sc_hd__clkbuf_8 fanout247 (.A(net773),
    .X(net1016));
 sky130_fd_sc_hd__buf_4 fanout248 (.A(net772),
    .X(net1017));
 sky130_fd_sc_hd__clkbuf_4 fanout249 (.A(net792),
    .X(net1018));
 sky130_fd_sc_hd__buf_4 fanout250 (.A(net791),
    .X(net1019));
 sky130_fd_sc_hd__buf_2 fanout251 (.A(net791),
    .X(net1020));
 sky130_fd_sc_hd__clkbuf_4 fanout252 (.A(net789),
    .X(net1021));
 sky130_fd_sc_hd__buf_2 fanout253 (.A(net789),
    .X(net1022));
 sky130_fd_sc_hd__buf_4 fanout254 (.A(net784),
    .X(net1023));
 sky130_fd_sc_hd__buf_4 fanout255 (.A(net783),
    .X(net1024));
 sky130_fd_sc_hd__clkbuf_2 fanout256 (.A(net783),
    .X(net1025));
 sky130_fd_sc_hd__clkbuf_4 fanout257 (.A(net782),
    .X(net1026));
 sky130_fd_sc_hd__buf_4 fanout258 (.A(net781),
    .X(net1027));
 sky130_fd_sc_hd__buf_4 fanout259 (.A(net780),
    .X(net1028));
 sky130_fd_sc_hd__buf_4 fanout260 (.A(net779),
    .X(net1029));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net753 (.A(net753),
    .X(clknet_0_net753));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net753 (.A(clknet_0_net753),
    .X(clknet_1_0__leaf_net753));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net753 (.A(clknet_0_net753),
    .X(clknet_1_1__leaf_net753));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net517 (.A(net517),
    .X(clknet_0_net517));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net517 (.A(clknet_0_net517),
    .X(clknet_1_0__leaf_net517));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net517 (.A(clknet_0_net517),
    .X(clknet_1_1__leaf_net517));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net522 (.A(net522),
    .X(clknet_0_net522));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net522 (.A(clknet_0_net522),
    .X(clknet_1_0__leaf_net522));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net522 (.A(clknet_0_net522),
    .X(clknet_1_1__leaf_net522));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net412 (.A(net412),
    .X(clknet_0_net412));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net412 (.A(clknet_0_net412),
    .X(clknet_1_0__leaf_net412));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net412 (.A(clknet_0_net412),
    .X(clknet_1_1__leaf_net412));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net411 (.A(net411),
    .X(clknet_0_net411));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net411 (.A(clknet_0_net411),
    .X(clknet_1_0__leaf_net411));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net411 (.A(clknet_0_net411),
    .X(clknet_1_1__leaf_net411));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net407 (.A(net407),
    .X(clknet_0_net407));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net407 (.A(clknet_0_net407),
    .X(clknet_1_0__leaf_net407));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net407 (.A(clknet_0_net407),
    .X(clknet_1_1__leaf_net407));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net549 (.A(net549),
    .X(clknet_0_net549));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net549 (.A(clknet_0_net549),
    .X(clknet_1_0__leaf_net549));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net549 (.A(clknet_0_net549),
    .X(clknet_1_1__leaf_net549));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net752 (.A(net752),
    .X(clknet_0_net752));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net752 (.A(clknet_0_net752),
    .X(clknet_1_0__leaf_net752));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net752 (.A(clknet_0_net752),
    .X(clknet_1_1__leaf_net752));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net409 (.A(net409),
    .X(clknet_0_net409));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net409 (.A(clknet_0_net409),
    .X(clknet_1_0__leaf_net409));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net409 (.A(clknet_0_net409),
    .X(clknet_1_1__leaf_net409));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net403 (.A(net403),
    .X(clknet_0_net403));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net403 (.A(clknet_0_net403),
    .X(clknet_1_0__leaf_net403));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net403 (.A(clknet_0_net403),
    .X(clknet_1_1__leaf_net403));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net413 (.A(net413),
    .X(clknet_0_net413));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net413 (.A(clknet_0_net413),
    .X(clknet_1_0__leaf_net413));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net413 (.A(clknet_0_net413),
    .X(clknet_1_1__leaf_net413));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net751 (.A(net751),
    .X(clknet_0_net751));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net751 (.A(clknet_0_net751),
    .X(clknet_1_0__leaf_net751));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net751 (.A(clknet_0_net751),
    .X(clknet_1_1__leaf_net751));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net410 (.A(net410),
    .X(clknet_0_net410));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net410 (.A(clknet_0_net410),
    .X(clknet_1_0__leaf_net410));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net410 (.A(clknet_0_net410),
    .X(clknet_1_1__leaf_net410));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net392 (.A(net392),
    .X(clknet_0_net392));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net392 (.A(clknet_0_net392),
    .X(clknet_1_0__leaf_net392));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net392 (.A(clknet_0_net392),
    .X(clknet_1_1__leaf_net392));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net496 (.A(net496),
    .X(clknet_0_net496));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net496 (.A(clknet_0_net496),
    .X(clknet_1_0__leaf_net496));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net496 (.A(clknet_0_net496),
    .X(clknet_1_1__leaf_net496));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net939 (.A(net939),
    .X(clknet_0_net939));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net939 (.A(clknet_0_net939),
    .X(clknet_1_0__leaf_net939));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net939 (.A(clknet_0_net939),
    .X(clknet_1_1__leaf_net939));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net735 (.A(net735),
    .X(clknet_0_net735));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net735 (.A(clknet_0_net735),
    .X(clknet_1_0__leaf_net735));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net735 (.A(clknet_0_net735),
    .X(clknet_1_1__leaf_net735));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net310 (.A(net310),
    .X(clknet_0_net310));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net310 (.A(clknet_0_net310),
    .X(clknet_1_0__leaf_net310));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net310 (.A(clknet_0_net310),
    .X(clknet_1_1__leaf_net310));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net307 (.A(net307),
    .X(clknet_0_net307));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net307 (.A(clknet_0_net307),
    .X(clknet_1_0__leaf_net307));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net307 (.A(clknet_0_net307),
    .X(clknet_1_1__leaf_net307));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net905 (.A(net905),
    .X(clknet_0_net905));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net905 (.A(clknet_0_net905),
    .X(clknet_1_0__leaf_net905));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net905 (.A(clknet_0_net905),
    .X(clknet_1_1__leaf_net905));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net908 (.A(net908),
    .X(clknet_0_net908));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net908 (.A(clknet_0_net908),
    .X(clknet_1_0__leaf_net908));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net908 (.A(clknet_0_net908),
    .X(clknet_1_1__leaf_net908));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net296 (.A(net296),
    .X(clknet_0_net296));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net296 (.A(clknet_0_net296),
    .X(clknet_1_0__leaf_net296));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net296 (.A(clknet_0_net296),
    .X(clknet_1_1__leaf_net296));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net904 (.A(net904),
    .X(clknet_0_net904));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net904 (.A(clknet_0_net904),
    .X(clknet_1_0__leaf_net904));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net904 (.A(clknet_0_net904),
    .X(clknet_1_1__leaf_net904));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net394 (.A(net394),
    .X(clknet_0_net394));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net394 (.A(clknet_0_net394),
    .X(clknet_1_0__leaf_net394));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net394 (.A(clknet_0_net394),
    .X(clknet_1_1__leaf_net394));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net734 (.A(net734),
    .X(clknet_0_net734));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net734 (.A(clknet_0_net734),
    .X(clknet_1_0__leaf_net734));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net734 (.A(clknet_0_net734),
    .X(clknet_1_1__leaf_net734));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net733 (.A(net733),
    .X(clknet_0_net733));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net733 (.A(clknet_0_net733),
    .X(clknet_1_0__leaf_net733));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net733 (.A(clknet_0_net733),
    .X(clknet_1_1__leaf_net733));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net714 (.A(net714),
    .X(clknet_0_net714));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net714 (.A(clknet_0_net714),
    .X(clknet_1_0__leaf_net714));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net714 (.A(clknet_0_net714),
    .X(clknet_1_1__leaf_net714));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net460 (.A(net460),
    .X(clknet_0_net460));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net460 (.A(clknet_0_net460),
    .X(clknet_1_0__leaf_net460));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net460 (.A(clknet_0_net460),
    .X(clknet_1_1__leaf_net460));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net504 (.A(net504),
    .X(clknet_0_net504));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net504 (.A(clknet_0_net504),
    .X(clknet_1_0__leaf_net504));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net504 (.A(clknet_0_net504),
    .X(clknet_1_1__leaf_net504));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net462 (.A(net462),
    .X(clknet_0_net462));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net462 (.A(clknet_0_net462),
    .X(clknet_1_0__leaf_net462));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net462 (.A(clknet_0_net462),
    .X(clknet_1_1__leaf_net462));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net458 (.A(net458),
    .X(clknet_0_net458));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net458 (.A(clknet_0_net458),
    .X(clknet_1_0__leaf_net458));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net458 (.A(clknet_0_net458),
    .X(clknet_1_1__leaf_net458));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net641 (.A(net641),
    .X(clknet_0_net641));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net641 (.A(clknet_0_net641),
    .X(clknet_1_0__leaf_net641));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net641 (.A(clknet_0_net641),
    .X(clknet_1_1__leaf_net641));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net518 (.A(net518),
    .X(clknet_0_net518));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net518 (.A(clknet_0_net518),
    .X(clknet_1_0__leaf_net518));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net518 (.A(clknet_0_net518),
    .X(clknet_1_1__leaf_net518));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net509 (.A(net509),
    .X(clknet_0_net509));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net509 (.A(clknet_0_net509),
    .X(clknet_1_0__leaf_net509));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net509 (.A(clknet_0_net509),
    .X(clknet_1_1__leaf_net509));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net260 (.A(net260),
    .X(clknet_0_net260));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net260 (.A(clknet_0_net260),
    .X(clknet_1_0__leaf_net260));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net260 (.A(clknet_0_net260),
    .X(clknet_1_1__leaf_net260));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net893 (.A(net893),
    .X(clknet_0_net893));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net893 (.A(clknet_0_net893),
    .X(clknet_1_0__leaf_net893));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net893 (.A(clknet_0_net893),
    .X(clknet_1_1__leaf_net893));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net401 (.A(net401),
    .X(clknet_0_net401));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net401 (.A(clknet_0_net401),
    .X(clknet_1_0__leaf_net401));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net401 (.A(clknet_0_net401),
    .X(clknet_1_1__leaf_net401));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net713 (.A(net713),
    .X(clknet_0_net713));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net713 (.A(clknet_0_net713),
    .X(clknet_1_0__leaf_net713));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net713 (.A(clknet_0_net713),
    .X(clknet_1_1__leaf_net713));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net405 (.A(net405),
    .X(clknet_0_net405));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net405 (.A(clknet_0_net405),
    .X(clknet_1_0__leaf_net405));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net405 (.A(clknet_0_net405),
    .X(clknet_1_1__leaf_net405));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net336 (.A(net336),
    .X(clknet_0_net336));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net336 (.A(clknet_0_net336),
    .X(clknet_1_0__leaf_net336));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net336 (.A(clknet_0_net336),
    .X(clknet_1_1__leaf_net336));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net894 (.A(net894),
    .X(clknet_0_net894));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net894 (.A(clknet_0_net894),
    .X(clknet_1_0__leaf_net894));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net894 (.A(clknet_0_net894),
    .X(clknet_1_1__leaf_net894));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net277 (.A(net277),
    .X(clknet_0_net277));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net277 (.A(clknet_0_net277),
    .X(clknet_1_0__leaf_net277));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net277 (.A(clknet_0_net277),
    .X(clknet_1_1__leaf_net277));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net422 (.A(net422),
    .X(clknet_0_net422));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net422 (.A(clknet_0_net422),
    .X(clknet_1_0__leaf_net422));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net422 (.A(clknet_0_net422),
    .X(clknet_1_1__leaf_net422));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net373 (.A(net373),
    .X(clknet_0_net373));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net373 (.A(clknet_0_net373),
    .X(clknet_1_0__leaf_net373));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net373 (.A(clknet_0_net373),
    .X(clknet_1_1__leaf_net373));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net378 (.A(net378),
    .X(clknet_0_net378));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net378 (.A(clknet_0_net378),
    .X(clknet_1_0__leaf_net378));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net378 (.A(clknet_0_net378),
    .X(clknet_1_1__leaf_net378));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net898 (.A(net898),
    .X(clknet_0_net898));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net898 (.A(clknet_0_net898),
    .X(clknet_1_0__leaf_net898));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net898 (.A(clknet_0_net898),
    .X(clknet_1_1__leaf_net898));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net712 (.A(net712),
    .X(clknet_0_net712));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net712 (.A(clknet_0_net712),
    .X(clknet_1_0__leaf_net712));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net712 (.A(clknet_0_net712),
    .X(clknet_1_1__leaf_net712));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net512 (.A(net512),
    .X(clknet_0_net512));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net512 (.A(clknet_0_net512),
    .X(clknet_1_0__leaf_net512));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net512 (.A(clknet_0_net512),
    .X(clknet_1_1__leaf_net512));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net465 (.A(net465),
    .X(clknet_0_net465));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net465 (.A(clknet_0_net465),
    .X(clknet_1_0__leaf_net465));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net465 (.A(clknet_0_net465),
    .X(clknet_1_1__leaf_net465));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net346 (.A(net346),
    .X(clknet_0_net346));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net346 (.A(clknet_0_net346),
    .X(clknet_1_0__leaf_net346));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net346 (.A(clknet_0_net346),
    .X(clknet_1_1__leaf_net346));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net616 (.A(net616),
    .X(clknet_0_net616));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net616 (.A(clknet_0_net616),
    .X(clknet_1_0__leaf_net616));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net616 (.A(clknet_0_net616),
    .X(clknet_1_1__leaf_net616));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net354 (.A(net354),
    .X(clknet_0_net354));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net354 (.A(clknet_0_net354),
    .X(clknet_1_0__leaf_net354));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net354 (.A(clknet_0_net354),
    .X(clknet_1_1__leaf_net354));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net615 (.A(net615),
    .X(clknet_0_net615));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net615 (.A(clknet_0_net615),
    .X(clknet_1_0__leaf_net615));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net615 (.A(clknet_0_net615),
    .X(clknet_1_1__leaf_net615));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net390 (.A(net390),
    .X(clknet_0_net390));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net390 (.A(clknet_0_net390),
    .X(clknet_1_0__leaf_net390));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net390 (.A(clknet_0_net390),
    .X(clknet_1_1__leaf_net390));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net353 (.A(net353),
    .X(clknet_0_net353));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net353 (.A(clknet_0_net353),
    .X(clknet_1_0__leaf_net353));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net353 (.A(net1061),
    .X(clknet_1_1__leaf_net353));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net273 (.A(net273),
    .X(clknet_0_net273));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net273 (.A(clknet_0_net273),
    .X(clknet_1_0__leaf_net273));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net273 (.A(clknet_0_net273),
    .X(clknet_1_1__leaf_net273));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net379 (.A(net379),
    .X(clknet_0_net379));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net379 (.A(clknet_0_net379),
    .X(clknet_1_0__leaf_net379));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net379 (.A(clknet_0_net379),
    .X(clknet_1_1__leaf_net379));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net276 (.A(net276),
    .X(clknet_0_net276));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net276 (.A(clknet_0_net276),
    .X(clknet_1_0__leaf_net276));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net276 (.A(clknet_0_net276),
    .X(clknet_1_1__leaf_net276));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net247 (.A(net247),
    .X(clknet_0_net247));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net247 (.A(clknet_0_net247),
    .X(clknet_1_0__leaf_net247));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net247 (.A(clknet_0_net247),
    .X(clknet_1_1__leaf_net247));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net695 (.A(net695),
    .X(clknet_0_net695));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net695 (.A(clknet_0_net695),
    .X(clknet_1_0__leaf_net695));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net695 (.A(clknet_0_net695),
    .X(clknet_1_1__leaf_net695));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net377 (.A(net377),
    .X(clknet_0_net377));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net377 (.A(clknet_0_net377),
    .X(clknet_1_0__leaf_net377));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net377 (.A(clknet_0_net377),
    .X(clknet_1_1__leaf_net377));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net399 (.A(net399),
    .X(clknet_0_net399));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net399 (.A(clknet_0_net399),
    .X(clknet_1_0__leaf_net399));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net399 (.A(clknet_0_net399),
    .X(clknet_1_1__leaf_net399));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net502 (.A(net502),
    .X(clknet_0_net502));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net502 (.A(clknet_0_net502),
    .X(clknet_1_0__leaf_net502));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net502 (.A(clknet_0_net502),
    .X(clknet_1_1__leaf_net502));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net532 (.A(net532),
    .X(clknet_0_net532));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net532 (.A(clknet_0_net532),
    .X(clknet_1_0__leaf_net532));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net532 (.A(clknet_0_net532),
    .X(clknet_1_1__leaf_net532));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net535 (.A(net535),
    .X(clknet_0_net535));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net535 (.A(clknet_0_net535),
    .X(clknet_1_0__leaf_net535));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net535 (.A(clknet_0_net535),
    .X(clknet_1_1__leaf_net535));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net167 (.A(net167),
    .X(clknet_0_net167));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net167 (.A(clknet_0_net167),
    .X(clknet_1_0__leaf_net167));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net167 (.A(clknet_0_net167),
    .X(clknet_1_1__leaf_net167));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net191 (.A(net191),
    .X(clknet_0_net191));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net191 (.A(clknet_0_net191),
    .X(clknet_1_0__leaf_net191));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net191 (.A(clknet_0_net191),
    .X(clknet_1_1__leaf_net191));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net887 (.A(net887),
    .X(clknet_0_net887));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net887 (.A(clknet_0_net887),
    .X(clknet_1_0__leaf_net887));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net887 (.A(clknet_0_net887),
    .X(clknet_1_1__leaf_net887));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net312 (.A(net312),
    .X(clknet_0_net312));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net312 (.A(clknet_0_net312),
    .X(clknet_1_0__leaf_net312));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net312 (.A(clknet_0_net312),
    .X(clknet_1_1__leaf_net312));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net168 (.A(net168),
    .X(clknet_0_net168));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net168 (.A(clknet_0_net168),
    .X(clknet_1_0__leaf_net168));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net168 (.A(clknet_0_net168),
    .X(clknet_1_1__leaf_net168));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net161 (.A(net161),
    .X(clknet_0_net161));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net161 (.A(clknet_0_net161),
    .X(clknet_1_0__leaf_net161));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net161 (.A(clknet_0_net161),
    .X(clknet_1_1__leaf_net161));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net263 (.A(net263),
    .X(clknet_0_net263));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net263 (.A(clknet_0_net263),
    .X(clknet_1_0__leaf_net263));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net263 (.A(clknet_0_net263),
    .X(clknet_1_1__leaf_net263));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net166 (.A(net166),
    .X(clknet_0_net166));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net166 (.A(clknet_0_net166),
    .X(clknet_1_0__leaf_net166));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net166 (.A(clknet_0_net166),
    .X(clknet_1_1__leaf_net166));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net283 (.A(net283),
    .X(clknet_0_net283));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net283 (.A(clknet_0_net283),
    .X(clknet_1_0__leaf_net283));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net283 (.A(clknet_0_net283),
    .X(clknet_1_1__leaf_net283));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net302 (.A(net302),
    .X(clknet_0_net302));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net302 (.A(clknet_0_net302),
    .X(clknet_1_0__leaf_net302));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net302 (.A(clknet_0_net302),
    .X(clknet_1_1__leaf_net302));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net178 (.A(net178),
    .X(clknet_0_net178));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net178 (.A(clknet_0_net178),
    .X(clknet_1_0__leaf_net178));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net178 (.A(clknet_0_net178),
    .X(clknet_1_1__leaf_net178));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net505 (.A(net505),
    .X(clknet_0_net505));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net505 (.A(clknet_0_net505),
    .X(clknet_1_0__leaf_net505));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net505 (.A(clknet_0_net505),
    .X(clknet_1_1__leaf_net505));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net922 (.A(net922),
    .X(clknet_0_net922));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net922 (.A(clknet_0_net922),
    .X(clknet_1_0__leaf_net922));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net922 (.A(clknet_0_net922),
    .X(clknet_1_1__leaf_net922));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net179 (.A(net179),
    .X(clknet_0_net179));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net179 (.A(clknet_0_net179),
    .X(clknet_1_0__leaf_net179));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net179 (.A(clknet_0_net179),
    .X(clknet_1_1__leaf_net179));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net613 (.A(net613),
    .X(clknet_0_net613));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net613 (.A(clknet_0_net613),
    .X(clknet_1_0__leaf_net613));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net613 (.A(clknet_0_net613),
    .X(clknet_1_1__leaf_net613));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net218 (.A(net218),
    .X(clknet_0_net218));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net218 (.A(clknet_0_net218),
    .X(clknet_1_0__leaf_net218));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net218 (.A(clknet_0_net218),
    .X(clknet_1_1__leaf_net218));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net219 (.A(net219),
    .X(clknet_0_net219));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net219 (.A(clknet_0_net219),
    .X(clknet_1_0__leaf_net219));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net219 (.A(clknet_0_net219),
    .X(clknet_1_1__leaf_net219));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net694 (.A(net694),
    .X(clknet_0_net694));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net694 (.A(clknet_0_net694),
    .X(clknet_1_0__leaf_net694));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net694 (.A(clknet_0_net694),
    .X(clknet_1_1__leaf_net694));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net935 (.A(net935),
    .X(clknet_0_net935));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net935 (.A(clknet_0_net935),
    .X(clknet_1_0__leaf_net935));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net935 (.A(clknet_0_net935),
    .X(clknet_1_1__leaf_net935));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net693 (.A(net693),
    .X(clknet_0_net693));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net693 (.A(clknet_0_net693),
    .X(clknet_1_0__leaf_net693));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net693 (.A(clknet_0_net693),
    .X(clknet_1_1__leaf_net693));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net895 (.A(net895),
    .X(clknet_0_net895));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net895 (.A(clknet_0_net895),
    .X(clknet_1_0__leaf_net895));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net895 (.A(clknet_0_net895),
    .X(clknet_1_1__leaf_net895));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net157 (.A(net157),
    .X(clknet_0_net157));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net157 (.A(clknet_0_net157),
    .X(clknet_1_0__leaf_net157));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net157 (.A(clknet_0_net157),
    .X(clknet_1_1__leaf_net157));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net293 (.A(net293),
    .X(clknet_0_net293));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net293 (.A(clknet_0_net293),
    .X(clknet_1_0__leaf_net293));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net293 (.A(clknet_0_net293),
    .X(clknet_1_1__leaf_net293));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net295 (.A(net295),
    .X(clknet_0_net295));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net295 (.A(clknet_0_net295),
    .X(clknet_1_0__leaf_net295));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net295 (.A(clknet_0_net295),
    .X(clknet_1_1__leaf_net295));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net900 (.A(net900),
    .X(clknet_0_net900));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net900 (.A(clknet_0_net900),
    .X(clknet_1_0__leaf_net900));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net900 (.A(clknet_0_net900),
    .X(clknet_1_1__leaf_net900));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net675 (.A(net675),
    .X(clknet_0_net675));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net675 (.A(clknet_0_net675),
    .X(clknet_1_0__leaf_net675));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net675 (.A(clknet_0_net675),
    .X(clknet_1_1__leaf_net675));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net284 (.A(net284),
    .X(clknet_0_net284));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net284 (.A(clknet_0_net284),
    .X(clknet_1_0__leaf_net284));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net284 (.A(clknet_0_net284),
    .X(clknet_1_1__leaf_net284));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net104 (.A(net104),
    .X(clknet_0_net104));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net104 (.A(clknet_0_net104),
    .X(clknet_1_0__leaf_net104));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net104 (.A(clknet_0_net104),
    .X(clknet_1_1__leaf_net104));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net890 (.A(net890),
    .X(clknet_0_net890));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net890 (.A(clknet_0_net890),
    .X(clknet_1_0__leaf_net890));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net890 (.A(clknet_0_net890),
    .X(clknet_1_1__leaf_net890));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net231 (.A(net231),
    .X(clknet_0_net231));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net231 (.A(clknet_0_net231),
    .X(clknet_1_0__leaf_net231));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net231 (.A(clknet_0_net231),
    .X(clknet_1_1__leaf_net231));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net333 (.A(net333),
    .X(clknet_0_net333));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net333 (.A(clknet_0_net333),
    .X(clknet_1_0__leaf_net333));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net333 (.A(clknet_0_net333),
    .X(clknet_1_1__leaf_net333));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net221 (.A(net221),
    .X(clknet_0_net221));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net221 (.A(clknet_0_net221),
    .X(clknet_1_0__leaf_net221));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net221 (.A(clknet_0_net221),
    .X(clknet_1_1__leaf_net221));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net674 (.A(net674),
    .X(clknet_0_net674));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net674 (.A(clknet_0_net674),
    .X(clknet_1_0__leaf_net674));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net674 (.A(clknet_0_net674),
    .X(clknet_1_1__leaf_net674));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net318 (.A(net318),
    .X(clknet_0_net318));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net318 (.A(clknet_0_net318),
    .X(clknet_1_0__leaf_net318));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net318 (.A(clknet_0_net318),
    .X(clknet_1_1__leaf_net318));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net199 (.A(net199),
    .X(clknet_0_net199));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net199 (.A(clknet_0_net199),
    .X(clknet_1_0__leaf_net199));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net199 (.A(clknet_0_net199),
    .X(clknet_1_1__leaf_net199));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net98 (.A(net98),
    .X(clknet_0_net98));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net98 (.A(clknet_0_net98),
    .X(clknet_1_0__leaf_net98));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net98 (.A(clknet_0_net98),
    .X(clknet_1_1__leaf_net98));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net100 (.A(net100),
    .X(clknet_0_net100));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net100 (.A(clknet_0_net100),
    .X(clknet_1_0__leaf_net100));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net100 (.A(clknet_0_net100),
    .X(clknet_1_1__leaf_net100));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net193 (.A(net193),
    .X(clknet_0_net193));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net193 (.A(clknet_0_net193),
    .X(clknet_1_0__leaf_net193));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net193 (.A(clknet_0_net193),
    .X(clknet_1_1__leaf_net193));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net916 (.A(net916),
    .X(clknet_0_net916));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net916 (.A(clknet_0_net916),
    .X(clknet_1_0__leaf_net916));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net916 (.A(clknet_0_net916),
    .X(clknet_1_1__leaf_net916));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net73 (.A(net73),
    .X(clknet_0_net73));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net73 (.A(clknet_0_net73),
    .X(clknet_1_0__leaf_net73));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net73 (.A(clknet_0_net73),
    .X(clknet_1_1__leaf_net73));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net530 (.A(net530),
    .X(clknet_0_net530));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net530 (.A(clknet_0_net530),
    .X(clknet_1_0__leaf_net530));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net530 (.A(clknet_0_net530),
    .X(clknet_1_1__leaf_net530));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net76 (.A(net76),
    .X(clknet_0_net76));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net76 (.A(clknet_0_net76),
    .X(clknet_1_0__leaf_net76));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net76 (.A(clknet_0_net76),
    .X(clknet_1_1__leaf_net76));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net182 (.A(net182),
    .X(clknet_0_net182));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net182 (.A(clknet_0_net182),
    .X(clknet_1_0__leaf_net182));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net182 (.A(clknet_0_net182),
    .X(clknet_1_1__leaf_net182));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net186 (.A(net186),
    .X(clknet_0_net186));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net186 (.A(clknet_0_net186),
    .X(clknet_1_0__leaf_net186));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net186 (.A(clknet_0_net186),
    .X(clknet_1_1__leaf_net186));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net78 (.A(net78),
    .X(clknet_0_net78));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net78 (.A(clknet_0_net78),
    .X(clknet_1_0__leaf_net78));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net78 (.A(clknet_0_net78),
    .X(clknet_1_1__leaf_net78));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net84 (.A(net84),
    .X(clknet_0_net84));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net84 (.A(clknet_0_net84),
    .X(clknet_1_0__leaf_net84));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net84 (.A(clknet_0_net84),
    .X(clknet_1_1__leaf_net84));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net938 (.A(net938),
    .X(clknet_0_net938));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net938 (.A(clknet_0_net938),
    .X(clknet_1_0__leaf_net938));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net938 (.A(clknet_0_net938),
    .X(clknet_1_1__leaf_net938));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net109 (.A(net109),
    .X(clknet_0_net109));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net109 (.A(clknet_0_net109),
    .X(clknet_1_0__leaf_net109));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net109 (.A(clknet_0_net109),
    .X(clknet_1_1__leaf_net109));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net651 (.A(net651),
    .X(clknet_0_net651));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net651 (.A(clknet_0_net651),
    .X(clknet_1_0__leaf_net651));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net651 (.A(clknet_0_net651),
    .X(clknet_1_1__leaf_net651));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net328 (.A(net328),
    .X(clknet_0_net328));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net328 (.A(clknet_0_net328),
    .X(clknet_1_0__leaf_net328));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net328 (.A(clknet_0_net328),
    .X(clknet_1_1__leaf_net328));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net113 (.A(net113),
    .X(clknet_0_net113));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net113 (.A(clknet_0_net113),
    .X(clknet_1_0__leaf_net113));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net113 (.A(clknet_0_net113),
    .X(clknet_1_1__leaf_net113));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net116 (.A(net116),
    .X(clknet_0_net116));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net116 (.A(clknet_0_net116),
    .X(clknet_1_0__leaf_net116));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net116 (.A(clknet_0_net116),
    .X(clknet_1_1__leaf_net116));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net923 (.A(net923),
    .X(clknet_0_net923));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net923 (.A(clknet_0_net923),
    .X(clknet_1_0__leaf_net923));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net923 (.A(clknet_0_net923),
    .X(clknet_1_1__leaf_net923));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net111 (.A(net111),
    .X(clknet_0_net111));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net111 (.A(clknet_0_net111),
    .X(clknet_1_0__leaf_net111));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net111 (.A(clknet_0_net111),
    .X(clknet_1_1__leaf_net111));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net83 (.A(net83),
    .X(clknet_0_net83));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net83 (.A(clknet_0_net83),
    .X(clknet_1_0__leaf_net83));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net83 (.A(clknet_0_net83),
    .X(clknet_1_1__leaf_net83));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net936 (.A(net936),
    .X(clknet_0_net936));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net936 (.A(clknet_0_net936),
    .X(clknet_1_0__leaf_net936));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net936 (.A(clknet_0_net936),
    .X(clknet_1_1__leaf_net936));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net79 (.A(net79),
    .X(clknet_0_net79));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net79 (.A(clknet_0_net79),
    .X(clknet_1_0__leaf_net79));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net79 (.A(clknet_0_net79),
    .X(clknet_1_1__leaf_net79));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net70 (.A(net70),
    .X(clknet_0_net70));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net70 (.A(clknet_0_net70),
    .X(clknet_1_0__leaf_net70));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net70 (.A(clknet_0_net70),
    .X(clknet_1_1__leaf_net70));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net74 (.A(net74),
    .X(clknet_0_net74));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net74 (.A(clknet_0_net74),
    .X(clknet_1_0__leaf_net74));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net74 (.A(clknet_0_net74),
    .X(clknet_1_1__leaf_net74));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net285 (.A(net285),
    .X(clknet_0_net285));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net285 (.A(clknet_0_net285),
    .X(clknet_1_0__leaf_net285));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net285 (.A(clknet_0_net285),
    .X(clknet_1_1__leaf_net285));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net72 (.A(net72),
    .X(clknet_0_net72));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net72 (.A(clknet_0_net72),
    .X(clknet_1_0__leaf_net72));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net72 (.A(clknet_0_net72),
    .X(clknet_1_1__leaf_net72));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net202 (.A(net202),
    .X(clknet_0_net202));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net202 (.A(clknet_0_net202),
    .X(clknet_1_0__leaf_net202));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net202 (.A(clknet_0_net202),
    .X(clknet_1_1__leaf_net202));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net208 (.A(net208),
    .X(clknet_0_net208));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net208 (.A(clknet_0_net208),
    .X(clknet_1_0__leaf_net208));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net208 (.A(clknet_0_net208),
    .X(clknet_1_1__leaf_net208));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net75 (.A(net75),
    .X(clknet_0_net75));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net75 (.A(clknet_0_net75),
    .X(clknet_1_0__leaf_net75));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net75 (.A(clknet_0_net75),
    .X(clknet_1_1__leaf_net75));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net77 (.A(net77),
    .X(clknet_0_net77));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net77 (.A(clknet_0_net77),
    .X(clknet_1_0__leaf_net77));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net77 (.A(clknet_0_net77),
    .X(clknet_1_1__leaf_net77));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net184 (.A(net184),
    .X(clknet_0_net184));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net184 (.A(clknet_0_net184),
    .X(clknet_1_0__leaf_net184));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net184 (.A(clknet_0_net184),
    .X(clknet_1_1__leaf_net184));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net288 (.A(net288),
    .X(clknet_0_net288));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net288 (.A(clknet_0_net288),
    .X(clknet_1_0__leaf_net288));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net288 (.A(clknet_0_net288),
    .X(clknet_1_1__leaf_net288));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net175 (.A(net175),
    .X(clknet_0_net175));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net175 (.A(clknet_0_net175),
    .X(clknet_1_0__leaf_net175));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net175 (.A(clknet_0_net175),
    .X(clknet_1_1__leaf_net175));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net673 (.A(net673),
    .X(clknet_0_net673));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net673 (.A(clknet_0_net673),
    .X(clknet_1_0__leaf_net673));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net673 (.A(clknet_0_net673),
    .X(clknet_1_1__leaf_net673));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net66 (.A(net66),
    .X(clknet_0_net66));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net66 (.A(clknet_0_net66),
    .X(clknet_1_0__leaf_net66));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net66 (.A(clknet_0_net66),
    .X(clknet_1_1__leaf_net66));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net174 (.A(net174),
    .X(clknet_0_net174));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net174 (.A(clknet_0_net174),
    .X(clknet_1_0__leaf_net174));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net174 (.A(clknet_0_net174),
    .X(clknet_1_1__leaf_net174));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer1 (.A(net31),
    .X(net1030));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer2 (.A(net1030),
    .X(net1031));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer3 (.A(net1033),
    .X(net1032));
 sky130_fd_sc_hd__mux4_1 clone4 (.A0(net1046),
    .A1(net1023),
    .A2(net1034),
    .A3(net1037),
    .S0(net26),
    .S1(net983),
    .X(net1033));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer5 (.A(net1035),
    .X(net1034));
 sky130_fd_sc_hd__mux4_1 clone6 (.A0(net1017),
    .A1(net1085),
    .A2(net1083),
    .A3(net1057),
    .S0(net27),
    .S1(net1079),
    .X(net1035));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer7 (.A(net872),
    .X(net1036));
 sky130_fd_sc_hd__a2111o_1 clone8 (.A1(net1005),
    .A2(net981),
    .B1(net778),
    .C1(net983),
    .D1(net987),
    .X(net1037));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer9 (.A(net34),
    .X(net1038));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer10 (.A(net1055),
    .X(net1039));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer11 (.A(net31),
    .X(net1040));
 sky130_fd_sc_hd__clkbuf_1 clone12 (.A(net21),
    .X(net1041));
 sky130_fd_sc_hd__clkbuf_1 clone13 (.A(net815),
    .X(net1042));
 sky130_fd_sc_hd__dlygate4sd3_1 rebuffer14 (.A(net1044),
    .X(net1043));
 sky130_fd_sc_hd__clkbuf_1 clone15 (.A(net776),
    .X(net1044));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer16 (.A(net345),
    .X(net1045));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer17 (.A(net1054),
    .X(net1046));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer18 (.A(net1046),
    .X(net1047));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer19 (.A(net1047),
    .X(net1048));
 sky130_fd_sc_hd__clkbuf_1 clone20 (.A(net33),
    .X(net1049));
 sky130_fd_sc_hd__clkbuf_1 clone21 (.A(net127),
    .X(net1050));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer22 (.A(net127),
    .X(net1051));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer23 (.A(net1051),
    .X(net1052));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer24 (.A(net1052),
    .X(net1053));
 sky130_fd_sc_hd__clkbuf_1 clone25 (.A(net23),
    .X(net1054));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer26 (.A(net1090),
    .X(net1055));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer27 (.A(net1055),
    .X(net1056));
 sky130_fd_sc_hd__clkbuf_1 clone28 (.A(net18),
    .X(net1057));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer29 (.A(net966),
    .X(net1058));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer30 (.A(net1058),
    .X(net1059));
 sky130_fd_sc_hd__clkbuf_1 clone31 (.A(net1013),
    .X(net1060));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer32 (.A(clknet_0_net353),
    .X(net1061));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer33 (.A(net815),
    .X(net1062));
 sky130_fd_sc_hd__clkbuf_1 clone34 (.A(net966),
    .X(net1063));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer35 (.A(clknet_1_0__leaf_net353),
    .X(net1064));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer36 (.A(clknet_1_0__leaf_net353),
    .X(net1065));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer37 (.A(clknet_1_0__leaf_net353),
    .X(net1066));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(net768),
    .X(net1067));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(net747),
    .X(net1068));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(net620),
    .X(net1069));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(net685),
    .X(net1070));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(net242),
    .X(net1071));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(net348),
    .X(net1072));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(net351),
    .X(net1073));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(net684),
    .X(net1074));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(net688),
    .X(net1075));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(net253),
    .X(net1076));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(net708),
    .X(net1077));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(net372),
    .X(net1078));
 sky130_fd_sc_hd__clkbuf_2 fanout1 (.A(net983),
    .X(net1079));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout2 (.A(net987),
    .X(net1080));
 sky130_fd_sc_hd__clkdlybuf4s15_2 fanout3 (.A(net1023),
    .X(net1081));
 sky130_fd_sc_hd__clkbuf_1 fanout4 (.A(net1017),
    .X(net1082));
 sky130_fd_sc_hd__clkbuf_1 fanout5 (.A(net1005),
    .X(net1083));
 sky130_fd_sc_hd__buf_6 fanout6 (.A(net778),
    .X(net1084));
 sky130_fd_sc_hd__clkbuf_1 fanout7 (.A(net775),
    .X(net1085));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_A (.DIODE(clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(in0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(in1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(in10));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(in11));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(in12));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(in13));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(in14));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(in15));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(in16));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(in17));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(in18));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(in19));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(in2));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(in20));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(in21));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(in22));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(in23));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(in24));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(in25));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(in26));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(in27));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_A (.DIODE(in28));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_A (.DIODE(in29));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_A (.DIODE(in3));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_A (.DIODE(in30));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_A (.DIODE(in31));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_A (.DIODE(in32));
 sky130_fd_sc_hd__diode_2 ANTENNA_input28_A (.DIODE(in33));
 sky130_fd_sc_hd__diode_2 ANTENNA_input29_A (.DIODE(in34));
 sky130_fd_sc_hd__diode_2 ANTENNA_input30_A (.DIODE(in35));
 sky130_fd_sc_hd__diode_2 ANTENNA_input31_A (.DIODE(in36));
 sky130_fd_sc_hd__diode_2 ANTENNA_input32_A (.DIODE(in37));
 sky130_fd_sc_hd__diode_2 ANTENNA_input33_A (.DIODE(in38));
 sky130_fd_sc_hd__diode_2 ANTENNA_input34_A (.DIODE(in39));
 sky130_fd_sc_hd__diode_2 ANTENNA_input35_A (.DIODE(in4));
 sky130_fd_sc_hd__diode_2 ANTENNA_input36_A (.DIODE(in40));
 sky130_fd_sc_hd__diode_2 ANTENNA_input37_A (.DIODE(in41));
 sky130_fd_sc_hd__diode_2 ANTENNA_input38_A (.DIODE(in42));
 sky130_fd_sc_hd__diode_2 ANTENNA_input39_A (.DIODE(in43));
 sky130_fd_sc_hd__diode_2 ANTENNA_input40_A (.DIODE(in44));
 sky130_fd_sc_hd__diode_2 ANTENNA_input41_A (.DIODE(in45));
 sky130_fd_sc_hd__diode_2 ANTENNA_input42_A (.DIODE(in46));
 sky130_fd_sc_hd__diode_2 ANTENNA_input43_A (.DIODE(in47));
 sky130_fd_sc_hd__diode_2 ANTENNA_input44_A (.DIODE(in48));
 sky130_fd_sc_hd__diode_2 ANTENNA_input45_A (.DIODE(in49));
 sky130_fd_sc_hd__diode_2 ANTENNA_input46_A (.DIODE(in5));
 sky130_fd_sc_hd__diode_2 ANTENNA_input47_A (.DIODE(in50));
 sky130_fd_sc_hd__diode_2 ANTENNA_input48_A (.DIODE(in51));
 sky130_fd_sc_hd__diode_2 ANTENNA_input49_A (.DIODE(in52));
 sky130_fd_sc_hd__diode_2 ANTENNA_input50_A (.DIODE(in53));
 sky130_fd_sc_hd__diode_2 ANTENNA_input51_A (.DIODE(in54));
 sky130_fd_sc_hd__diode_2 ANTENNA_input52_A (.DIODE(in55));
 sky130_fd_sc_hd__diode_2 ANTENNA_input53_A (.DIODE(in56));
 sky130_fd_sc_hd__diode_2 ANTENNA_input54_A (.DIODE(in57));
 sky130_fd_sc_hd__diode_2 ANTENNA_input55_A (.DIODE(in58));
 sky130_fd_sc_hd__diode_2 ANTENNA_input56_A (.DIODE(in59));
 sky130_fd_sc_hd__diode_2 ANTENNA_input57_A (.DIODE(in6));
 sky130_fd_sc_hd__diode_2 ANTENNA_input58_A (.DIODE(in60));
 sky130_fd_sc_hd__diode_2 ANTENNA_input59_A (.DIODE(in61));
 sky130_fd_sc_hd__diode_2 ANTENNA_input60_A (.DIODE(in62));
 sky130_fd_sc_hd__diode_2 ANTENNA_input61_A (.DIODE(in63));
 sky130_fd_sc_hd__diode_2 ANTENNA_input62_A (.DIODE(in64));
 sky130_fd_sc_hd__diode_2 ANTENNA_input63_A (.DIODE(in65));
 sky130_fd_sc_hd__diode_2 ANTENNA_input64_A (.DIODE(in66));
 sky130_fd_sc_hd__diode_2 ANTENNA_input65_A (.DIODE(in67));
 sky130_fd_sc_hd__diode_2 ANTENNA_input66_A (.DIODE(in68));
 sky130_fd_sc_hd__diode_2 ANTENNA_input67_A (.DIODE(in69));
 sky130_fd_sc_hd__diode_2 ANTENNA_input68_A (.DIODE(in7));
 sky130_fd_sc_hd__diode_2 ANTENNA_input69_A (.DIODE(in70));
 sky130_fd_sc_hd__diode_2 ANTENNA_input70_A (.DIODE(in71));
 sky130_fd_sc_hd__diode_2 ANTENNA_input71_A (.DIODE(in72));
 sky130_fd_sc_hd__diode_2 ANTENNA_input72_A (.DIODE(in73));
 sky130_fd_sc_hd__diode_2 ANTENNA_input73_A (.DIODE(in74));
 sky130_fd_sc_hd__diode_2 ANTENNA_input74_A (.DIODE(in75));
 sky130_fd_sc_hd__diode_2 ANTENNA_input75_A (.DIODE(in76));
 sky130_fd_sc_hd__diode_2 ANTENNA_input76_A (.DIODE(in77));
 sky130_fd_sc_hd__diode_2 ANTENNA_input77_A (.DIODE(in78));
 sky130_fd_sc_hd__diode_2 ANTENNA_input78_A (.DIODE(in79));
 sky130_fd_sc_hd__diode_2 ANTENNA_input79_A (.DIODE(in8));
 sky130_fd_sc_hd__diode_2 ANTENNA_input80_A (.DIODE(in80));
 sky130_fd_sc_hd__diode_2 ANTENNA_input81_A (.DIODE(in81));
 sky130_fd_sc_hd__diode_2 ANTENNA_input82_A (.DIODE(in82));
 sky130_fd_sc_hd__diode_2 ANTENNA_input83_A (.DIODE(in83));
 sky130_fd_sc_hd__diode_2 ANTENNA_input84_A (.DIODE(in84));
 sky130_fd_sc_hd__diode_2 ANTENNA_input85_A (.DIODE(in85));
 sky130_fd_sc_hd__diode_2 ANTENNA_input86_A (.DIODE(in86));
 sky130_fd_sc_hd__diode_2 ANTENNA_input87_A (.DIODE(in87));
 sky130_fd_sc_hd__diode_2 ANTENNA_input88_A (.DIODE(in88));
 sky130_fd_sc_hd__diode_2 ANTENNA_input89_A (.DIODE(in89));
 sky130_fd_sc_hd__diode_2 ANTENNA_input90_A (.DIODE(in9));
 sky130_fd_sc_hd__diode_2 ANTENNA_input91_A (.DIODE(in90));
 sky130_fd_sc_hd__diode_2 ANTENNA_input92_A (.DIODE(in91));
 sky130_fd_sc_hd__diode_2 ANTENNA_input93_A (.DIODE(in92));
 sky130_fd_sc_hd__diode_2 ANTENNA_input94_A (.DIODE(in93));
 sky130_fd_sc_hd__diode_2 ANTENNA_input95_A (.DIODE(in94));
 sky130_fd_sc_hd__diode_2 ANTENNA_input96_A (.DIODE(in95));
 sky130_fd_sc_hd__diode_2 ANTENNA_input97_A (.DIODE(in96));
 sky130_fd_sc_hd__diode_2 ANTENNA_input98_A (.DIODE(in97));
 sky130_fd_sc_hd__diode_2 ANTENNA_input99_A (.DIODE(in98));
 sky130_fd_sc_hd__diode_2 ANTENNA_input100_A (.DIODE(in99));
 sky130_fd_sc_hd__diode_2 ANTENNA_c372_A1 (.DIODE(net0));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_A0 (.DIODE(net0));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_A2 (.DIODE(net0));
 sky130_fd_sc_hd__diode_2 ANTENNA_c108_A1 (.DIODE(net0));
 sky130_fd_sc_hd__diode_2 ANTENNA_c105_S1 (.DIODE(net0));
 sky130_fd_sc_hd__diode_2 ANTENNA_c100_X (.DIODE(net0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout230_A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_A0 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_c763_S0 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_A2 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_c101_X (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_c757_A1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_A3 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_A2 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_A2 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c239_Q (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c566_A1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c533_D (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_A0 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c408_A3 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c277_S0 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c269_C1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_B1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c265_A1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c264_X (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_A0 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_A2 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_c664_A2 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_c546_A2 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_A0 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_c408_A2 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_c286_S0 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_c272_RESET_B (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_c266_X (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_c530_A2 (.DIODE(net1091));
 sky130_fd_sc_hd__diode_2 ANTENNA_c533_RESET_B (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_c276_S1 (.DIODE(net1091));
 sky130_fd_sc_hd__diode_2 ANTENNA_c273_SCD (.DIODE(net1091));
 sky130_fd_sc_hd__diode_2 ANTENNA_c271_A1 (.DIODE(net1091));
 sky130_fd_sc_hd__diode_2 ANTENNA_c269_A1 (.DIODE(net1091));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_X (.DIODE(net1091));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_A0 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_c397_A2 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_A1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_S0 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_c274_D (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_c270_A2 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_c269_X (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_c676_A1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_c664_S0 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_c403_B1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_c401_D1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_A3 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_c272_Q_N (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_c670_A1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA_c412_A3 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_A0 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA_c276_A2 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA_c273_RESET_B (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA_c272_Q (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA_c311_A2 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_A2 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_A2 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_c273_Q_N (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_c427_A0 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c397_A1 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_A0 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c273_Q (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c676_A2 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_c545_S0 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_S1 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_c275_A2 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_c274_Q_N (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_c679_A3 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_c673_A0 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_c279_A1 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_c276_A0 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_c274_Q (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_A0 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_S0 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_A0 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_A2 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_A0 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_A0 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_c278_A1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_c276_S0 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_c275_X (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout193_A (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA_c536_C1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA_c665_A2 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA_c679_A2 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA_c680_A1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_X (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout179_A (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_A2 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_A2 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_A2 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_A3 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_X (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_A1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_A3 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_c430_S0 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_A3 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_A0 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_A2 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_X (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_A0 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_A1 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA_c437_A1 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_A1 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA_c297_A2 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_X (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_A0 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_S0 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_A0 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA_c297_A0 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_A2 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_X (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_A0 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA_c344_A1 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA_c323_A2 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA_c313_A1 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_X (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout218_A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c405_D (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c264_C1 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_A2 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_X (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_A0 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_S0 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_A2 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_A2 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_A2 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_A2 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_X (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_c371_A2 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_c370_A3 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_A0 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_A2 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_A2 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_A3 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_c241_A1 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_c103_X (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout228_A (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_A2 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA_c266_A3 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA_c275_A1 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA_c277_A1 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA_c134_X (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_A0 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_A0 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_c350_A1 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_X (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone12_A (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout217_A (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_A0 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_X (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_c531_A2 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout213_A (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_c537_C1 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_c136_X (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge878_RESET_B (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_X (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer26_A (.DIODE(net1090));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone25_A (.DIODE(net1099));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout212_A (.DIODE(net1099));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_A2 (.DIODE(net1099));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_X (.DIODE(net1099));
 sky130_fd_sc_hd__diode_2 ANTENNA_c687_A1 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_S0 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA_c681_A0 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA_c667_A3 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_A1 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_A2 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_A3 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA_c416_S0 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA_c398_D (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_X (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout190_A (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_c701_A3 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_c397_X (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_C1 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA_c446_A1 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_A1 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_A2 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA_c398_Q_N (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_A0 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c561_B1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c414_A0 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c400_D (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c398_Q (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c546_A1 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA_c544_A3 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA_c539_C1 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA_c532_RESET_B (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA_c400_SCE (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA_c399_X (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_A3 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_A2 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c405_SCD (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c400_Q_N (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_A0 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_A1 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_A0 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_c414_A1 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_c400_Q (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_A3 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_A1 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA_c533_SCD (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_A2 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA_c411_SCD (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA_c406_B1 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA_c405_Q_N (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA_c766_A0 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_A1 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA_c633_A3 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA_c539_B1 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA_c412_A2 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA_c409_D (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA_c408_A0 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA_c405_Q (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net247_A (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c406_X (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_A3 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_A0 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_A0 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_A1 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_c544_A0 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_c534_RESET_B (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_c402_RESET_B (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_c269_D1 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_A0 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_X (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_A2 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_A3 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA_c409_Q_N (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_A1 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA_c415_A0 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA_c409_Q (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA_c587_A3 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_A0 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_A3 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_SCD (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA_c411_Q_N (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_A0 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_A1 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_A0 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA_c413_D (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA_c411_Q (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_A0 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_A1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_A1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA_c413_Q (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone4_S0 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_A0 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c416_A0 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c400_RESET_B (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c266_S0 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c265_A2 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_S0 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_A3 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_A2 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_A1 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c140_X (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone6_S0 (.DIODE(net1087));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout211_A (.DIODE(net1087));
 sky130_fd_sc_hd__diode_2 ANTENNA_c143_S0 (.DIODE(net1087));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_A1 (.DIODE(net1087));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_B1 (.DIODE(net1087));
 sky130_fd_sc_hd__diode_2 ANTENNA_c404_S1 (.DIODE(net1087));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_X (.DIODE(net1087));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_A0 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_A3 (.DIODE(net1086));
 sky130_fd_sc_hd__diode_2 ANTENNA_c148_A1 (.DIODE(net1086));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_A2 (.DIODE(net1086));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_A2 (.DIODE(net1086));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_A3 (.DIODE(net1086));
 sky130_fd_sc_hd__diode_2 ANTENNA_c143_X (.DIODE(net1086));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout210_A (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout209_A (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_X (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_c762_A0 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_S1 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_A3 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c231_A1 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c230_A2 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c108_A0 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c104_X (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout208_A (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_A1 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_A1 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_X (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net310_A (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_X (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout205_A (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_A1 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_A1 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_S0 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_c148_X (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone20_A (.DIODE(net1088));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout204_A (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_A0 (.DIODE(net1088));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_A1 (.DIODE(net1088));
 sky130_fd_sc_hd__diode_2 ANTENNA_c765_A0 (.DIODE(net1088));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_X (.DIODE(net1088));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net346_A (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA_c531_X (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_A2 (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA_c662_B1 (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA_c541_SCD (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA_c535_C1 (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA_c533_Q_N (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_A2 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_A1 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_A2 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_A2 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_c670_D1 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_c537_B1 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_c529_SCE (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_c404_A0 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_A0 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_S0 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_X (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_A0 (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_A3 (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_A2 (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA_c660_A2 (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA_c537_A1 (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA_c533_Q (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA_c427_A1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c410_D (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c401_A2 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_A3 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c272_D (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c269_B1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c159_D1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_B1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_S1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_A1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_X (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_S0 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA_c668_S0 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA_c666_D1 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA_c549_S0 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA_c548_SCE (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA_c547_A1 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA_c546_D1 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA_c544_S0 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA_c543_B1 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA_c541_Q_N (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA_c767_B1 (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA_c760_B1 (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_A0 (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_A3 (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_A1 (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A2 (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_S0 (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_A1 (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA_c545_A1 (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA_c542_A1 (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA_c541_Q (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout194_A (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_A3 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c720_A1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_S0 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_X (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold49_A (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_A2 (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_Q_N (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_A2 (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA_c691_A1 (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_A3 (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_A0 (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA_c554_A1 (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_X (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_A0 (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA_c610_A3 (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_B1 (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_A1 (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA_c560_Q (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout199_A (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_A2 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_A1 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_X (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_c434_A0 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_A1 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_S0 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_A2 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_c158_A0 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_X (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_c743_A0 (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_A2 (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_A1 (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA_c586_A2 (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_A1 (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_X (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA_c742_A1 (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_A1 (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_A3 (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_A1 (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_A2 (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_X (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_A0 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_S0 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_S1 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_A1 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_A0 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_A1 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_S0 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_A1 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_X (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_c565_A2 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_c559_A2 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_c216_A3 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_c198_B1 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_Q_N (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge869_GCLK (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA_c613_X (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA_c577_A1 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_A1 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_A1 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_A1 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_Q (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout188_A (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_A1 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_X (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_A1 (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_A0 (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_A2 (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_S0 (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_S1 (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA_c676_X (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_A0 (.DIODE(net474));
 sky130_fd_sc_hd__diode_2 ANTENNA_c693_A2 (.DIODE(net474));
 sky130_fd_sc_hd__diode_2 ANTENNA_c680_A0 (.DIODE(net474));
 sky130_fd_sc_hd__diode_2 ANTENNA_c679_A1 (.DIODE(net474));
 sky130_fd_sc_hd__diode_2 ANTENNA_c678_X (.DIODE(net474));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_S0 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_c184_A3 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_c180_A1 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_A3 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_A3 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_Q_N (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_c742_A0 (.DIODE(net488));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_A2 (.DIODE(net488));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_A2 (.DIODE(net488));
 sky130_fd_sc_hd__diode_2 ANTENNA_c703_A1 (.DIODE(net488));
 sky130_fd_sc_hd__diode_2 ANTENNA_c695_A3 (.DIODE(net488));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_X (.DIODE(net488));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_A2 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_c424_A0 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_A0 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_A1 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_A1 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_Q (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_c767_A1 (.DIODE(net495));
 sky130_fd_sc_hd__diode_2 ANTENNA_c765_S0 (.DIODE(net495));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_A0 (.DIODE(net495));
 sky130_fd_sc_hd__diode_2 ANTENNA_c701_A1 (.DIODE(net495));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_X (.DIODE(net495));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_A0 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_A0 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_A0 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_c109_S1 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_c108_S1 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_c107_A0 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_c106_X (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge856_D (.DIODE(net507));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_X (.DIODE(net507));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout185_A (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_S0 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_X (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout184_A (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_A0 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_A1 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_X (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge797_Q (.DIODE(net570));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_S1 (.DIODE(net570));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_A2 (.DIODE(net570));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_A2 (.DIODE(net570));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_A3 (.DIODE(net570));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_S1 (.DIODE(net570));
 sky130_fd_sc_hd__diode_2 ANTENNA_c218_C1 (.DIODE(net570));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_D1 (.DIODE(net570));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge799_Q_N (.DIODE(net572));
 sky130_fd_sc_hd__diode_2 ANTENNA_c256_S1 (.DIODE(net572));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_S0 (.DIODE(net572));
 sky130_fd_sc_hd__diode_2 ANTENNA_c232_S0 (.DIODE(net572));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_S0 (.DIODE(net572));
 sky130_fd_sc_hd__diode_2 ANTENNA_c184_S0 (.DIODE(net572));
 sky130_fd_sc_hd__diode_2 ANTENNA_c182_S0 (.DIODE(net572));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge799_Q (.DIODE(net573));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_A2 (.DIODE(net573));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_A3 (.DIODE(net573));
 sky130_fd_sc_hd__diode_2 ANTENNA_c261_S1 (.DIODE(net573));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_S1 (.DIODE(net573));
 sky130_fd_sc_hd__diode_2 ANTENNA_c194_S0 (.DIODE(net573));
 sky130_fd_sc_hd__diode_2 ANTENNA_c190_S1 (.DIODE(net573));
 sky130_fd_sc_hd__diode_2 ANTENNA_c180_S1 (.DIODE(net573));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge801_Q (.DIODE(net576));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_A3 (.DIODE(net576));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_B1 (.DIODE(net576));
 sky130_fd_sc_hd__diode_2 ANTENNA_c283_A3 (.DIODE(net576));
 sky130_fd_sc_hd__diode_2 ANTENNA_c279_S0 (.DIODE(net576));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge805_Q (.DIODE(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_S1 (.DIODE(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA_c560_SCE (.DIODE(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_C1 (.DIODE(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA_c543_D1 (.DIODE(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA_c541_SET_B (.DIODE(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA_c540_SCE (.DIODE(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge811_Q (.DIODE(net586));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_C1 (.DIODE(net586));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_S1 (.DIODE(net586));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_S1 (.DIODE(net586));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_D1 (.DIODE(net586));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_D1 (.DIODE(net586));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge826_Q (.DIODE(net604));
 sky130_fd_sc_hd__diode_2 ANTENNA_c564_A3 (.DIODE(net604));
 sky130_fd_sc_hd__diode_2 ANTENNA_c559_C1 (.DIODE(net604));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_A3 (.DIODE(net604));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_A3 (.DIODE(net604));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_A2 (.DIODE(net604));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_A3 (.DIODE(net604));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_S0 (.DIODE(net604));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_A2 (.DIODE(net604));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge827_Q (.DIODE(net605));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_S0 (.DIODE(net605));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_A3 (.DIODE(net605));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_A3 (.DIODE(net605));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_A3 (.DIODE(net605));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_S0 (.DIODE(net605));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge829_Q (.DIODE(net607));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_S0 (.DIODE(net607));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_S0 (.DIODE(net607));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_S0 (.DIODE(net607));
 sky130_fd_sc_hd__diode_2 ANTENNA_c238_S1 (.DIODE(net607));
 sky130_fd_sc_hd__diode_2 ANTENNA_c232_S1 (.DIODE(net607));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_S1 (.DIODE(net607));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_S1 (.DIODE(net607));
 sky130_fd_sc_hd__diode_2 ANTENNA_c220_S1 (.DIODE(net607));
 sky130_fd_sc_hd__diode_2 ANTENNA_c218_D1 (.DIODE(net607));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout198_A (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_A3 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_X (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge839_Q_N (.DIODE(net617));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_A3 (.DIODE(net617));
 sky130_fd_sc_hd__diode_2 ANTENNA_c700_S0 (.DIODE(net617));
 sky130_fd_sc_hd__diode_2 ANTENNA_c698_A3 (.DIODE(net617));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge839_Q (.DIODE(net618));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_S0 (.DIODE(net618));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_S0 (.DIODE(net618));
 sky130_fd_sc_hd__diode_2 ANTENNA_c544_S1 (.DIODE(net618));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge840_Q_N (.DIODE(net619));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_S0 (.DIODE(net619));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_A2 (.DIODE(net619));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_S0 (.DIODE(net619));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_A1 (.DIODE(net619));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_A2 (.DIODE(net619));
 sky130_fd_sc_hd__diode_2 ANTENNA_c218_A1 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_A2 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_A3 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA_c183_A2 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_A1 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA_c180_A2 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_X (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_A3 (.DIODE(net623));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_S0 (.DIODE(net623));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_S0 (.DIODE(net623));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_A3 (.DIODE(net623));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_A2 (.DIODE(net623));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_S0 (.DIODE(net623));
 sky130_fd_sc_hd__diode_2 ANTENNA_c216_S1 (.DIODE(net623));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_S1 (.DIODE(net623));
 sky130_fd_sc_hd__diode_2 ANTENNA_c184_S1 (.DIODE(net623));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_D1 (.DIODE(net623));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_S1 (.DIODE(net623));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_A3 (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_S0 (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_A3 (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_A3 (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA_c212_C1 (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_D1 (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_S1 (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_S1 (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_S0 (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_S1 (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_S1 (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_S1 (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_SET_B (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge851_Q (.DIODE(net633));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_A3 (.DIODE(net633));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_S0 (.DIODE(net633));
 sky130_fd_sc_hd__diode_2 ANTENNA_c373_S0 (.DIODE(net633));
 sky130_fd_sc_hd__diode_2 ANTENNA_c369_C1 (.DIODE(net633));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge858_Q_N (.DIODE(net639));
 sky130_fd_sc_hd__diode_2 ANTENNA_c757_S0 (.DIODE(net639));
 sky130_fd_sc_hd__diode_2 ANTENNA_c743_A2 (.DIODE(net639));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_S0 (.DIODE(net639));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge863_Q (.DIODE(net645));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_A2 (.DIODE(net645));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_S0 (.DIODE(net645));
 sky130_fd_sc_hd__diode_2 ANTENNA_c582_S1 (.DIODE(net645));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_A2 (.DIODE(net645));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_A3 (.DIODE(net645));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_A3 (.DIODE(net645));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge864_Q (.DIODE(net646));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_S1 (.DIODE(net646));
 sky130_fd_sc_hd__diode_2 ANTENNA_c613_S0 (.DIODE(net646));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_A3 (.DIODE(net646));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_A3 (.DIODE(net646));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_A2 (.DIODE(net646));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_A2 (.DIODE(net646));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge865_Q (.DIODE(net647));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_A2 (.DIODE(net647));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_A3 (.DIODE(net647));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_A3 (.DIODE(net647));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_S0 (.DIODE(net647));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_A3 (.DIODE(net647));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_S0 (.DIODE(net647));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_S0 (.DIODE(net647));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_S0 (.DIODE(net647));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge881_SET_B (.DIODE(net652));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge872_X (.DIODE(net652));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge873_Q_N (.DIODE(net653));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_S0 (.DIODE(net653));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_A2 (.DIODE(net653));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_S0 (.DIODE(net653));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge877_Q (.DIODE(net658));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_A3 (.DIODE(net658));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_S1 (.DIODE(net658));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_A3 (.DIODE(net658));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_S1 (.DIODE(net658));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_A3 (.DIODE(net658));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_S0 (.DIODE(net658));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge881_Q (.DIODE(net663));
 sky130_fd_sc_hd__diode_2 ANTENNA_c769_S1 (.DIODE(net663));
 sky130_fd_sc_hd__diode_2 ANTENNA_c767_D1 (.DIODE(net663));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_A3 (.DIODE(net663));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_A3 (.DIODE(net663));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_S0 (.DIODE(net663));
 sky130_fd_sc_hd__diode_2 ANTENNA_c674_S1 (.DIODE(net663));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge883_Q (.DIODE(net664));
 sky130_fd_sc_hd__diode_2 ANTENNA_c744_A3 (.DIODE(net664));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_S0 (.DIODE(net664));
 sky130_fd_sc_hd__diode_2 ANTENNA_c691_S0 (.DIODE(net664));
 sky130_fd_sc_hd__diode_2 ANTENNA_c677_S0 (.DIODE(net664));
 sky130_fd_sc_hd__diode_2 ANTENNA_c676_S0 (.DIODE(net664));
 sky130_fd_sc_hd__diode_2 ANTENNA_c675_C1 (.DIODE(net664));
 sky130_fd_sc_hd__diode_2 ANTENNA_s887_Q_N (.DIODE(net668));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_A3 (.DIODE(net668));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_S0 (.DIODE(net668));
 sky130_fd_sc_hd__diode_2 ANTENNA_c561_C1 (.DIODE(net668));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_S0 (.DIODE(net668));
 sky130_fd_sc_hd__diode_2 ANTENNA_s887_Q (.DIODE(net669));
 sky130_fd_sc_hd__diode_2 ANTENNA_c743_A3 (.DIODE(net669));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_S0 (.DIODE(net669));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_A3 (.DIODE(net669));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_S0 (.DIODE(net669));
 sky130_fd_sc_hd__diode_2 ANTENNA_s889_Q (.DIODE(net671));
 sky130_fd_sc_hd__diode_2 ANTENNA_c496_S1 (.DIODE(net671));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_S1 (.DIODE(net671));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_A2 (.DIODE(net671));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_A3 (.DIODE(net671));
 sky130_fd_sc_hd__diode_2 ANTENNA_c234_S0 (.DIODE(net671));
 sky130_fd_sc_hd__diode_2 ANTENNA_c221_S0 (.DIODE(net671));
 sky130_fd_sc_hd__diode_2 ANTENNA_c203_D1 (.DIODE(net671));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_S1 (.DIODE(net671));
 sky130_fd_sc_hd__diode_2 ANTENNA_s890_Q (.DIODE(net672));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_S0 (.DIODE(net672));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_A3 (.DIODE(net672));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_S0 (.DIODE(net672));
 sky130_fd_sc_hd__diode_2 ANTENNA_c562_SET_B (.DIODE(net672));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_S0 (.DIODE(net672));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_S0 (.DIODE(net672));
 sky130_fd_sc_hd__diode_2 ANTENNA_c221_S1 (.DIODE(net672));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_S1 (.DIODE(net672));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net675_A (.DIODE(net675));
 sky130_fd_sc_hd__diode_2 ANTENNA_s894_GCLK (.DIODE(net675));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_A1 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_A1 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_A0 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_A1 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c191_S0 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_A0 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c184_X (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_s898_Q (.DIODE(net681));
 sky130_fd_sc_hd__diode_2 ANTENNA_c762_A3 (.DIODE(net681));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_S1 (.DIODE(net681));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_S0 (.DIODE(net681));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_A3 (.DIODE(net681));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_D1 (.DIODE(net681));
 sky130_fd_sc_hd__diode_2 ANTENNA_s900_Q (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_S0 (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_S0 (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_S0 (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_S0 (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_A3 (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_S1 (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_S0 (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold45_A (.DIODE(net684));
 sky130_fd_sc_hd__diode_2 ANTENNA_s901_Q (.DIODE(net684));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_S0 (.DIODE(net684));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_S0 (.DIODE(net684));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_S0 (.DIODE(net684));
 sky130_fd_sc_hd__diode_2 ANTENNA_c279_S1 (.DIODE(net684));
 sky130_fd_sc_hd__diode_2 ANTENNA_c277_S1 (.DIODE(net684));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold41_A (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA_s902_Q (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_C1 (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_S0 (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_A3 (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA_c283_S0 (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_S1 (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA_s903_Q_N (.DIODE(net686));
 sky130_fd_sc_hd__diode_2 ANTENNA_c424_A3 (.DIODE(net686));
 sky130_fd_sc_hd__diode_2 ANTENNA_c399_D1 (.DIODE(net686));
 sky130_fd_sc_hd__diode_2 ANTENNA_c398_SET_B (.DIODE(net686));
 sky130_fd_sc_hd__diode_2 ANTENNA_c397_D1 (.DIODE(net686));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_A3 (.DIODE(net686));
 sky130_fd_sc_hd__diode_2 ANTENNA_c295_S1 (.DIODE(net686));
 sky130_fd_sc_hd__diode_2 ANTENNA_s903_Q (.DIODE(net687));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_A2 (.DIODE(net687));
 sky130_fd_sc_hd__diode_2 ANTENNA_c538_SET_B (.DIODE(net687));
 sky130_fd_sc_hd__diode_2 ANTENNA_c532_SET_B (.DIODE(net687));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_A2 (.DIODE(net687));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_S0 (.DIODE(net687));
 sky130_fd_sc_hd__diode_2 ANTENNA_c283_S1 (.DIODE(net687));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold46_A (.DIODE(net688));
 sky130_fd_sc_hd__diode_2 ANTENNA_s904_Q_N (.DIODE(net688));
 sky130_fd_sc_hd__diode_2 ANTENNA_c673_S0 (.DIODE(net688));
 sky130_fd_sc_hd__diode_2 ANTENNA_c668_S1 (.DIODE(net688));
 sky130_fd_sc_hd__diode_2 ANTENNA_c663_C1 (.DIODE(net688));
 sky130_fd_sc_hd__diode_2 ANTENNA_c660_D1 (.DIODE(net688));
 sky130_fd_sc_hd__diode_2 ANTENNA_c554_S1 (.DIODE(net688));
 sky130_fd_sc_hd__diode_2 ANTENNA_c531_C1 (.DIODE(net688));
 sky130_fd_sc_hd__diode_2 ANTENNA_c529_SET_B (.DIODE(net688));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_A3 (.DIODE(net688));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout227_A (.DIODE(net689));
 sky130_fd_sc_hd__diode_2 ANTENNA_c680_A3 (.DIODE(net689));
 sky130_fd_sc_hd__diode_2 ANTENNA_s904_Q (.DIODE(net689));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout224_A (.DIODE(net691));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_S0 (.DIODE(net691));
 sky130_fd_sc_hd__diode_2 ANTENNA_s906_Q (.DIODE(net691));
 sky130_fd_sc_hd__diode_2 ANTENNA_s907_Q (.DIODE(net692));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_S0 (.DIODE(net692));
 sky130_fd_sc_hd__diode_2 ANTENNA_c556_S1 (.DIODE(net692));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_D1 (.DIODE(net692));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_S0 (.DIODE(net692));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_S0 (.DIODE(net692));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_A2 (.DIODE(net692));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_S0 (.DIODE(net692));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net693_A (.DIODE(net693));
 sky130_fd_sc_hd__diode_2 ANTENNA_s908_GCLK (.DIODE(net693));
 sky130_fd_sc_hd__diode_2 ANTENNA_s911_Q (.DIODE(net697));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_S0 (.DIODE(net697));
 sky130_fd_sc_hd__diode_2 ANTENNA_c561_D1 (.DIODE(net697));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_S0 (.DIODE(net697));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_S1 (.DIODE(net697));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_S1 (.DIODE(net697));
 sky130_fd_sc_hd__diode_2 ANTENNA_s912_Q_N (.DIODE(net698));
 sky130_fd_sc_hd__diode_2 ANTENNA_c586_S1 (.DIODE(net698));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_S1 (.DIODE(net698));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_S0 (.DIODE(net698));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_S1 (.DIODE(net698));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_S1 (.DIODE(net698));
 sky130_fd_sc_hd__diode_2 ANTENNA_s913_Q_N (.DIODE(net699));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_S0 (.DIODE(net699));
 sky130_fd_sc_hd__diode_2 ANTENNA_c703_S0 (.DIODE(net699));
 sky130_fd_sc_hd__diode_2 ANTENNA_c555_A3 (.DIODE(net699));
 sky130_fd_sc_hd__diode_2 ANTENNA_s913_Q (.DIODE(net700));
 sky130_fd_sc_hd__diode_2 ANTENNA_c744_S1 (.DIODE(net700));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_S0 (.DIODE(net700));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_C1 (.DIODE(net700));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_S1 (.DIODE(net700));
 sky130_fd_sc_hd__diode_2 ANTENNA_s914_Q (.DIODE(net701));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_A3 (.DIODE(net701));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_S0 (.DIODE(net701));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_S0 (.DIODE(net701));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_S0 (.DIODE(net701));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_S0 (.DIODE(net701));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_S1 (.DIODE(net701));
 sky130_fd_sc_hd__diode_2 ANTENNA_c313_S0 (.DIODE(net701));
 sky130_fd_sc_hd__diode_2 ANTENNA_c311_S1 (.DIODE(net701));
 sky130_fd_sc_hd__diode_2 ANTENNA_s916_Q (.DIODE(net703));
 sky130_fd_sc_hd__diode_2 ANTENNA_c364_S1 (.DIODE(net703));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_S0 (.DIODE(net703));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_S0 (.DIODE(net703));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_S1 (.DIODE(net703));
 sky130_fd_sc_hd__diode_2 ANTENNA_c323_S1 (.DIODE(net703));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_S1 (.DIODE(net703));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_S1 (.DIODE(net703));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_S1 (.DIODE(net703));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_S1 (.DIODE(net703));
 sky130_fd_sc_hd__diode_2 ANTENNA_s917_Q (.DIODE(net704));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_S0 (.DIODE(net704));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_S1 (.DIODE(net704));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_S1 (.DIODE(net704));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_S1 (.DIODE(net704));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_S1 (.DIODE(net704));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap221_A (.DIODE(net705));
 sky130_fd_sc_hd__diode_2 ANTENNA_s918_Q (.DIODE(net705));
 sky130_fd_sc_hd__diode_2 ANTENNA_c615_A3 (.DIODE(net705));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_S1 (.DIODE(net705));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_A3 (.DIODE(net705));
 sky130_fd_sc_hd__diode_2 ANTENNA_s919_Q (.DIODE(net707));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_S0 (.DIODE(net707));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_S1 (.DIODE(net707));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_S1 (.DIODE(net707));
 sky130_fd_sc_hd__diode_2 ANTENNA_c350_S0 (.DIODE(net707));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold48_A (.DIODE(net708));
 sky130_fd_sc_hd__diode_2 ANTENNA_s920_Q_N (.DIODE(net708));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_S1 (.DIODE(net708));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_S1 (.DIODE(net708));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_S0 (.DIODE(net708));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_S0 (.DIODE(net708));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_A1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_A0 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_A3 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_A1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_c238_A3 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_c215_A1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_c190_A0 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_A2 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_X (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_s922_Q (.DIODE(net710));
 sky130_fd_sc_hd__diode_2 ANTENNA_c611_A3 (.DIODE(net710));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_S1 (.DIODE(net710));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_S1 (.DIODE(net710));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_S1 (.DIODE(net710));
 sky130_fd_sc_hd__diode_2 ANTENNA_s923_Q (.DIODE(net711));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_S0 (.DIODE(net711));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_S0 (.DIODE(net711));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_S1 (.DIODE(net711));
 sky130_fd_sc_hd__diode_2 ANTENNA_c366_S1 (.DIODE(net711));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_S1 (.DIODE(net711));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_S1 (.DIODE(net711));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net713_A (.DIODE(net713));
 sky130_fd_sc_hd__diode_2 ANTENNA_s925_GCLK (.DIODE(net713));
 sky130_fd_sc_hd__diode_2 ANTENNA_s928_Q (.DIODE(net718));
 sky130_fd_sc_hd__diode_2 ANTENNA_c723_S1 (.DIODE(net718));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_S1 (.DIODE(net718));
 sky130_fd_sc_hd__diode_2 ANTENNA_c702_S1 (.DIODE(net718));
 sky130_fd_sc_hd__diode_2 ANTENNA_s929_Q (.DIODE(net720));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_S1 (.DIODE(net720));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_S1 (.DIODE(net720));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_S0 (.DIODE(net720));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_S1 (.DIODE(net720));
 sky130_fd_sc_hd__diode_2 ANTENNA_s930_Q (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_S1 (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_A3 (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_A2 (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA_c555_S1 (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_S1 (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_A1 (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA_c431_S0 (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA_s932_Q (.DIODE(net723));
 sky130_fd_sc_hd__diode_2 ANTENNA_c611_S0 (.DIODE(net723));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_S1 (.DIODE(net723));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_S1 (.DIODE(net723));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_S1 (.DIODE(net723));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_S0 (.DIODE(net723));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_S0 (.DIODE(net723));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_S0 (.DIODE(net723));
 sky130_fd_sc_hd__diode_2 ANTENNA_s933_Q (.DIODE(net724));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_S0 (.DIODE(net724));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_S0 (.DIODE(net724));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_S1 (.DIODE(net724));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_A3 (.DIODE(net724));
 sky130_fd_sc_hd__diode_2 ANTENNA_c427_S1 (.DIODE(net724));
 sky130_fd_sc_hd__diode_2 ANTENNA_s934_Q (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_S1 (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA_c437_A3 (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA_c430_S1 (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_S1 (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net73_A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_X (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_s937_Q (.DIODE(net730));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_S0 (.DIODE(net730));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_S0 (.DIODE(net730));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_S0 (.DIODE(net730));
 sky130_fd_sc_hd__diode_2 ANTENNA_c686_S0 (.DIODE(net730));
 sky130_fd_sc_hd__diode_2 ANTENNA_c564_S0 (.DIODE(net730));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_D1 (.DIODE(net730));
 sky130_fd_sc_hd__diode_2 ANTENNA_c437_S1 (.DIODE(net730));
 sky130_fd_sc_hd__diode_2 ANTENNA_s938_Q (.DIODE(net731));
 sky130_fd_sc_hd__diode_2 ANTENNA_c747_S1 (.DIODE(net731));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_S1 (.DIODE(net731));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_S1 (.DIODE(net731));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_S1 (.DIODE(net731));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_S0 (.DIODE(net731));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_S0 (.DIODE(net731));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_S1 (.DIODE(net731));
 sky130_fd_sc_hd__diode_2 ANTENNA_s943_Q_N (.DIODE(net736));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_S0 (.DIODE(net736));
 sky130_fd_sc_hd__diode_2 ANTENNA_c615_S0 (.DIODE(net736));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_A3 (.DIODE(net736));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_S0 (.DIODE(net736));
 sky130_fd_sc_hd__diode_2 ANTENNA_s943_Q (.DIODE(net737));
 sky130_fd_sc_hd__diode_2 ANTENNA_c766_S0 (.DIODE(net737));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_S1 (.DIODE(net737));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_S0 (.DIODE(net737));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_S1 (.DIODE(net737));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_S1 (.DIODE(net737));
 sky130_fd_sc_hd__diode_2 ANTENNA_s945_Q_N (.DIODE(net739));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_S1 (.DIODE(net739));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_S1 (.DIODE(net739));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_S1 (.DIODE(net739));
 sky130_fd_sc_hd__diode_2 ANTENNA_s945_Q (.DIODE(net740));
 sky130_fd_sc_hd__diode_2 ANTENNA_c762_S1 (.DIODE(net740));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_S1 (.DIODE(net740));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_S1 (.DIODE(net740));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_S0 (.DIODE(net740));
 sky130_fd_sc_hd__diode_2 ANTENNA_s946_Q (.DIODE(net741));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_S1 (.DIODE(net741));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_S1 (.DIODE(net741));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_S1 (.DIODE(net741));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_S1 (.DIODE(net741));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_S1 (.DIODE(net741));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_S1 (.DIODE(net741));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_S1 (.DIODE(net741));
 sky130_fd_sc_hd__diode_2 ANTENNA_s952_Q (.DIODE(net748));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_S1 (.DIODE(net748));
 sky130_fd_sc_hd__diode_2 ANTENNA_c560_SET_B (.DIODE(net748));
 sky130_fd_sc_hd__diode_2 ANTENNA_s955_Q (.DIODE(net750));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_S1 (.DIODE(net750));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_S0 (.DIODE(net750));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_S1 (.DIODE(net750));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_S1 (.DIODE(net750));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_S0 (.DIODE(net750));
 sky130_fd_sc_hd__diode_2 ANTENNA_s964_Q (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_c724_S0 (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_S0 (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_S0 (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_S1 (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_c680_S0 (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_c679_S1 (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_s966_Q (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_S1 (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_S1 (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA_c724_S1 (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_S1 (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA_c680_S1 (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA_c678_S1 (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA_s971_Q (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_S1 (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c739_S1 (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_S1 (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_S1 (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net79_A (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_X (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_A0 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_S1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_A2 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_A1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_c216_A2 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_S1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_S1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_c206_A1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_A2 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_c198_X (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net84_A (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_X (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_c482_A0 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_A1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_S1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_A3 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_A2 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_c208_A1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_c203_X (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_A0 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_A3 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_A1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_Q (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_A0 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_A2 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_c614_A2 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_c502_A3 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_A1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_A3 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_c206_X (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_A0 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_A3 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_c212_A1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_B1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_X (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_c373_A2 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_c364_A0 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_A3 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_A1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_c221_A0 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_C1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_c218_B1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_S1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_c216_A1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_X (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_X (.DIODE(net484));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_A3 (.DIODE(net484));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_A3 (.DIODE(net484));
 sky130_fd_sc_hd__diode_2 ANTENNA_c554_S0 (.DIODE(net484));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_A2 (.DIODE(net484));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_A2 (.DIODE(net484));
 sky130_fd_sc_hd__diode_2 ANTENNA_c259_A1 (.DIODE(net484));
 sky130_fd_sc_hd__diode_2 ANTENNA_c208_A0 (.DIODE(net484));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_A2 (.DIODE(net484));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_A1 (.DIODE(net484));
 sky130_fd_sc_hd__diode_2 ANTENNA_c112_A2 (.DIODE(net484));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_X (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_A0 (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_A2 (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_A1 (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_A1 (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_c270_A1 (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_c267_A1 (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_c266_A1 (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_S0 (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_A2 (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_c140_A3 (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout248_A (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_X (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_A0 (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_c271_S0 (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout247_A (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_X (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA_c760_A1 (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_A3 (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout7_A (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_X (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_c529_D (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone15_A (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout237_A (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_X (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A0 (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_S0 (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_S0 (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout235_A (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_X (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout6_A (.DIODE(net778));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone8_B1 (.DIODE(net778));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_X (.DIODE(net778));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout260_A (.DIODE(net779));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_X (.DIODE(net779));
 sky130_fd_sc_hd__diode_2 ANTENNA_c685_S1 (.DIODE(net779));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_A3 (.DIODE(net779));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_A2 (.DIODE(net779));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_A2 (.DIODE(net779));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout259_A (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_X (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_A2 (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA_c587_A2 (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA_c399_A1 (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA_c398_SCD (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout258_A (.DIODE(net781));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_X (.DIODE(net781));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_A2 (.DIODE(net781));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_A3 (.DIODE(net781));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout257_A (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_X (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_c685_S0 (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout256_A (.DIODE(net783));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout255_A (.DIODE(net783));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_X (.DIODE(net783));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout254_A (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_X (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA_c745_S0 (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_A0 (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_X (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_A1 (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_A0 (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_A3 (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_A2 (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_A1 (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_c230_A3 (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_A3 (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_C1 (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_c114_A (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_X (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c763_A2 (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A2 (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_A1 (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_A1 (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c198_D1 (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_A0 (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_B1 (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_D1 (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_X (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_A0 (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_A3 (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA_c182_A1 (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_A2 (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_A1 (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout253_A (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout252_A (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_X (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_X (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA_c262_A0 (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA_c180_A3 (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_A1 (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_D1 (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA_c120_C1 (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA_c115_B1 (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout251_A (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout250_A (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_X (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout249_A (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_X (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_c614_A0 (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_X (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_A0 (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_A1 (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_A1 (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c264_A1 (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c182_A0 (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_A1 (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_A3 (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_B1 (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c134_A2 (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_B1 (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_X (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_A0 (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_c158_A3 (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_A2 (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_c121_A2 (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_c120_A1 (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_X (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_A0 (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_A1 (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_A1 (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_A3 (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_A1 (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_c286_A3 (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_A0 (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_A2 (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_SCD (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_S0 (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_X (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_A0 (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_A3 (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA_c565_S0 (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_A0 (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_S0 (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_A3 (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA_c261_A0 (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA_c117_D1 (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA_c102_A2 (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA_input28_X (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA_c633_A2 (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_A1 (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_A3 (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_A0 (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_A0 (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_A1 (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_A2 (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA_input29_X (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA_c494_A1 (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_A0 (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_A2 (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA_c321_A2 (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_S0 (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_A2 (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_C1 (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_A0 (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA_c127_A2 (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA_input30_X (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c557_A1 (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_A0 (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c431_A1 (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_A1 (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_A1 (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_input31_X (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_A2 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_A0 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_A3 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_A2 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_B1 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c159_A1 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_input32_X (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_A0 (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_A1 (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_A2 (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_A0 (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_c239_D (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_c232_A1 (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_input34_X (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_A0 (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_A1 (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA_c159_A2 (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA_input35_X (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_A2 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A3 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_A2 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_A3 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c582_S0 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_A2 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_A3 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c340_A2 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c278_A0 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_S0 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_input36_X (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_A1 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_A2 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_c502_S1 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_A3 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_A2 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_A3 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_A2 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_SCE (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_A1 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_B1 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_input37_X (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_A2 (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_A2 (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA_c494_A3 (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA_c434_A1 (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_A3 (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_A2 (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_S0 (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA_input38_X (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_c263_A3 (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_A0 (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_c215_A3 (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_A2 (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_c122_A1 (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_c121_S1 (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_input39_X (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_A3 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_A0 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_A1 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_A0 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_A3 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c556_S0 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_A3 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_input40_X (.DIODE(net809));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A1 (.DIODE(net809));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_A1 (.DIODE(net809));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_A1 (.DIODE(net809));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_A2 (.DIODE(net809));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_A3 (.DIODE(net809));
 sky130_fd_sc_hd__diode_2 ANTENNA_c203_A1 (.DIODE(net809));
 sky130_fd_sc_hd__diode_2 ANTENNA_c198_C1 (.DIODE(net809));
 sky130_fd_sc_hd__diode_2 ANTENNA_input42_X (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_c586_A0 (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_A3 (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_A2 (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_A0 (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_c180_A0 (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_input43_X (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_A0 (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_S1 (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_S1 (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_input44_X (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_A0 (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c220_A1 (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_A1 (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c182_A2 (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c109_A3 (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout245_A (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_input45_X (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_S0 (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_c586_S0 (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_A2 (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_A1 (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer33_A (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone13_A (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout244_A (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_input46_X (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_input48_X (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_A1 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_A0 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_A1 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c198_A2 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c127_S1 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c110_A2 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_input49_X (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_A2 (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_A0 (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c577_A3 (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_A0 (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_A2 (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_input50_X (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_S0 (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_A1 (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_S1 (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_input51_X (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_c190_S0 (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_A1 (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_A2 (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_A1 (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_input52_X (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_A1 (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_A0 (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_A1 (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_A2 (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_S0 (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_c482_A2 (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_S0 (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_input53_X (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_A0 (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_A1 (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_A3 (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_c323_A3 (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_c262_S1 (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_c104_S1 (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_input56_X (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_c368_A2 (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_A3 (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_A0 (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_c261_A3 (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_c258_S0 (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_c183_S0 (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_c122_A2 (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_c119_B1 (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_c111_A1 (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_input58_X (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_A0 (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_A2 (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_c232_A2 (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_A2 (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_c208_S0 (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_A1 (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_B1 (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_c100_A3 (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_input59_X (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_S0 (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_A1 (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_A3 (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_A2 (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_A1 (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_C1 (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_c114_B (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_c103_A2 (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_input61_X (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA_c346_A0 (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_A0 (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_A1 (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_A3 (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_A3 (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_A2 (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA_input62_X (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_A0 (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c221_A3 (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_A3 (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_B1 (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c106_S1 (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c105_A1 (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_input64_X (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_A0 (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_A3 (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_A3 (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_S0 (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_c102_A1 (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_c100_A2 (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_input67_X (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_A3 (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_A0 (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_A2 (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA_input68_X (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c369_B1 (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_A0 (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_A1 (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_A2 (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c271_A0 (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c228_A2 (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c136_A2 (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c112_A1 (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c110_B1 (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c107_S0 (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_input69_X (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_A1 (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_A0 (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_A3 (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_A0 (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_c231_A3 (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_A1 (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_A2 (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_c105_A2 (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_c103_A3 (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_c101_S0 (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_input71_X (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_A0 (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_A2 (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_c257_A2 (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_c205_A1 (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_c108_S0 (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_input72_X (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_S0 (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_A0 (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_A1 (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_A2 (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_A0 (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_A2 (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_A2 (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_c203_A2 (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_input73_X (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_A2 (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_A0 (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_A2 (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_A2 (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_input75_X (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_A0 (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_A3 (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_C1 (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_input80_X (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_C1 (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_D (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_input83_X (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_A1 (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_A0 (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_input85_X (.DIODE(net854));
 sky130_fd_sc_hd__diode_2 ANTENNA_c236_A0 (.DIODE(net854));
 sky130_fd_sc_hd__diode_2 ANTENNA_c206_B1 (.DIODE(net854));
 sky130_fd_sc_hd__diode_2 ANTENNA_input87_X (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_A3 (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_A0 (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_input88_X (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A1 (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_A1 (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_c107_S1 (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_c102_A0 (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_input89_X (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_A2 (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_A3 (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_A1 (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_c238_A2 (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_c105_A0 (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout232_A (.DIODE(net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_input90_X (.DIODE(net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_c765_A1 (.DIODE(net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_A2 (.DIODE(net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_input92_X (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_A2 (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_c633_S0 (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_A2 (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_A1 (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_c234_A3 (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_A2 (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_c100_A0 (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_input93_X (.DIODE(net862));
 sky130_fd_sc_hd__diode_2 ANTENNA_c237_A2 (.DIODE(net862));
 sky130_fd_sc_hd__diode_2 ANTENNA_c222_A2 (.DIODE(net862));
 sky130_fd_sc_hd__diode_2 ANTENNA_c120_B1 (.DIODE(net862));
 sky130_fd_sc_hd__diode_2 ANTENNA_c104_A1 (.DIODE(net862));
 sky130_fd_sc_hd__diode_2 ANTENNA_input94_X (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_c129_A0 (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_c116_B1 (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_c111_C1 (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_c109_A0 (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_c100_S1 (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout231_A (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_input96_X (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c130_A3 (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c128_A3 (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c121_S0 (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c119_C1 (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_input98_X (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A0 (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_A1 (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c365_A0 (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c100_A1 (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_input99_X (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_A3 (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_A0 (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_A1 (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_c104_A0 (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_output104_A (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_s912_Q (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_S1 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_S0 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_S1 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_S1 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_S1 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_output105_A (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_A1 (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_A1 (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_Q (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_output107_A (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA_s959_Q (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_S0 (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA_output108_A (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge856_Q (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_S0 (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_A3 (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_A3 (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_output114_A (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_s888_Q (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_S1 (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_S0 (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_S1 (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_output119_A (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_A0 (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_c563_A2 (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_c562_Q (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_output120_A (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_s944_Q (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_A3 (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_S1 (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_S1 (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_output122_A (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_s953_Q (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_S1 (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_S1 (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c548_SET_B (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c547_S1 (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c545_S1 (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_output127_A (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c482_A1 (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_A2 (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_A2 (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_X (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout189_A (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_output128_A (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_A1 (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c286_A1 (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c158_X (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net898_A (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c434_X (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_output132_A (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge882_Q (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_S0 (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_A3 (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_S1 (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_S0 (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_S0 (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_A3 (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_S0 (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_output133_A (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge795_Q (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_A2 (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_A3 (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_S1 (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_output134_A (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_s895_Q (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_S1 (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_c231_S1 (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net904_A (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_X (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net905_A (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_X (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_output138_A (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge830_Q (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_S0 (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_A3 (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_c260_S1 (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_output140_A (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge803_Q (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_S1 (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_A3 (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_S0 (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_A3 (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_A3 (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_A3 (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_A3 (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_A3 (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_output142_A (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge885_Q (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_A3 (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_A3 (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_S0 (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_output143_A (.DIODE(net912));
 sky130_fd_sc_hd__diode_2 ANTENNA_s891_Q (.DIODE(net912));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_S0 (.DIODE(net912));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_S1 (.DIODE(net912));
 sky130_fd_sc_hd__diode_2 ANTENNA_c350_A2 (.DIODE(net912));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_S0 (.DIODE(net912));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_S0 (.DIODE(net912));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_S1 (.DIODE(net912));
 sky130_fd_sc_hd__diode_2 ANTENNA_c183_S1 (.DIODE(net912));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_S1 (.DIODE(net912));
 sky130_fd_sc_hd__diode_2 ANTENNA_output144_A (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA_s949_Q (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA_c743_S1 (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_S1 (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_S1 (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA_c482_S1 (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA_output146_A (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge878_Q (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_S0 (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_A3 (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_c724_A3 (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_c372_S1 (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_c366_A3 (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_output148_A (.DIODE(net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_c369_A1 (.DIODE(net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_c364_A2 (.DIODE(net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_c111_B1 (.DIODE(net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_c102_X (.DIODE(net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_output150_A (.DIODE(net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge868_Q (.DIODE(net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_c373_S1 (.DIODE(net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_c372_S0 (.DIODE(net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_c371_S1 (.DIODE(net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_A3 (.DIODE(net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_A2 (.DIODE(net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_output151_A (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge884_Q (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_c344_S0 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_S0 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_c340_S1 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_output158_A (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c263_S1 (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c262_S0 (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c261_S0 (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c259_A3 (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c256_A2 (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c237_A1 (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c231_X (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_output159_A (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge862_Q (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_S0 (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_A3 (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_S0 (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_S0 (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_A2 (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_output162_A (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_c760_C1 (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_A3 (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_A3 (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_A3 (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_output165_A (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_S1 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_A1 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c340_A1 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c260_A1 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c258_A1 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_S0 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_A0 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_S0 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_X (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net935_A (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_X (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net938_A (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge870_GCLK (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net939_A (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c571_X (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_output171_A (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge884_Q_N (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_S0 (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_A2 (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_c241_S1 (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout179_X (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c415_A2 (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_A1 (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_A3 (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_A3 (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_A2 (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_A0 (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c340_S0 (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_A3 (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_A2 (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_A3 (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout180_X (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c272_SCE (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c407_C1 (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c273_SET_B (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_S0 (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c279_A0 (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c276_A3 (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c274_SET_B (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_A1 (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c277_A3 (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c278_A3 (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout181_X (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_c283_A2 (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_c402_SCE (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_c398_RESET_B (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout180_A (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_A3 (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_A0 (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout182_X (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_c405_SET_B (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_c677_A1 (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_c565_A3 (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_RESET_B (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_c542_D1 (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_c533_SCE (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_c528_S1 (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_c411_RESET_B (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_c529_SCD (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout181_A (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout183_X (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout182_A (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c761_A1 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_A2 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_A2 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_A1 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_A2 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_A1 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout184_X (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_A2 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c582_A1 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c558_S0 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c235_A1 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_A3 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_A2 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_A1 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_A0 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_S0 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_S0 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout185_X (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c431_A3 (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c424_A1 (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_A2 (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c311_A0 (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_S0 (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_A0 (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c502_A1 (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_S0 (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c350_A0 (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_S0 (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout186_X (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_S0 (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_A3 (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_S0 (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_A2 (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_c180_S0 (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_S0 (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_A3 (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_A0 (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_RESET_B (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_A3 (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout187_X (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_A2 (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout186_A (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_S1 (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_c238_S0 (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_c236_S1 (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_S1 (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_c222_A3 (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_SET_B (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_A3 (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_S0 (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout188_X (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_A1 (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_A2 (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_A2 (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c560_SCD (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c554_A3 (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_A3 (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c765_A3 (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_A1 (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_A2 (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout187_A (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout189_X (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_A3 (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_SCE (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_S1 (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_SET_B (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c159_C1 (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_A1 (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c222_A1 (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_A1 (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c183_A3 (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_A2 (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout190_X (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_c700_A0 (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_c691_A3 (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_A1 (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_c678_A1 (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_c532_D (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_c528_S0 (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_c416_A3 (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_c409_RESET_B (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_c406_A2 (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_c399_A2 (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout191_X (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c413_SCD (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c403_C1 (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c399_B1 (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c279_A3 (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_A2 (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c278_A2 (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c276_A1 (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c272_SCD (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c271_A2 (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c274_SCE (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout192_X (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_B1 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c528_A0 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout191_A (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_A2 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_A1 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_A0 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout193_X (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c295_A1 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_A1 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_A1 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c283_A1 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_A0 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c763_A1 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_A2 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_A2 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_A1 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_A1 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout194_X (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_A3 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_A0 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_S0 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c702_A3 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_A1 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_A1 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c231_A0 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_A3 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_S1 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_A0 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_C1 (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout195_X (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c564_A1 (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_A3 (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_A2 (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c275_A0 (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone34_A (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer29_A (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout197_X (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_A2 (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c562_SCD (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c560_D (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_S0 (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout196_A (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout198_X (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_A1 (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_A2 (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_A1 (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_A1 (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_A3 (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_A1 (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_A0 (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_A3 (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_A2 (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_A0 (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout199_X (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_S0 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_A1 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_S0 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_A1 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_A2 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_A1 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_A2 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_A2 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c340_A3 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_S1 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_D1 (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout200_X (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_c275_A3 (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_c273_SCE (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_A0 (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_A0 (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_A1 (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_A3 (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_A1 (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_c257_A3 (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_c229_S0 (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout201_X (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_output116_A (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_c537_D1 (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_c536_A2 (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_c530_B1 (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_A2 (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout202_X (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_S1 (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_S1 (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_A3 (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_c769_A0 (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_A2 (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_A2 (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_A2 (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_c323_A0 (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_c206_C1 (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_D1 (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_c265_C1 (.DIODE(net1093));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout203_X (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c685_A1 (.DIODE(net1093));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_S1 (.DIODE(net1093));
 sky130_fd_sc_hd__diode_2 ANTENNA_c669_C1 (.DIODE(net1093));
 sky130_fd_sc_hd__diode_2 ANTENNA_c543_A2 (.DIODE(net1093));
 sky130_fd_sc_hd__diode_2 ANTENNA_c286_A0 (.DIODE(net1093));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_C1 (.DIODE(net1093));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_D1 (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout204_X (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_A1 (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_A2 (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_A2 (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_A1 (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout205_X (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_c270_B1 (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_A0 (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_A3 (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_A2 (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_A1 (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_A2 (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_A0 (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_c434_S0 (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_c297_A1 (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_c190_A2 (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout206_X (.DIODE(net1092));
 sky130_fd_sc_hd__diode_2 ANTENNA_c566_A3 (.DIODE(net1092));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_A2 (.DIODE(net1092));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_A3 (.DIODE(net1092));
 sky130_fd_sc_hd__diode_2 ANTENNA_c258_A2 (.DIODE(net1092));
 sky130_fd_sc_hd__diode_2 ANTENNA_c257_S0 (.DIODE(net1092));
 sky130_fd_sc_hd__diode_2 ANTENNA_c236_A1 (.DIODE(net1092));
 sky130_fd_sc_hd__diode_2 ANTENNA_c229_A1 (.DIODE(net1092));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_S1 (.DIODE(net1092));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_D1 (.DIODE(net1092));
 sky130_fd_sc_hd__diode_2 ANTENNA_c148_A0 (.DIODE(net1092));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout207_X (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_output103_A (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A2 (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_c739_S0 (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_A0 (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_c665_B1 (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout208_X (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_A1 (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_A2 (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_c685_A3 (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_c397_C1 (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_B1 (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_A2 (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_S1 (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_c295_A0 (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_A2 (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_c206_D1 (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_c267_D1 (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout209_X (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_A2 (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_S0 (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_A0 (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_c321_A3 (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_SCE (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_RESET_B (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_A0 (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_c148_S0 (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_A2 (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout210_X (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c759_A2 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_A1 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c746_S0 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c660_B1 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c610_A2 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout211_X (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c272_SET_B (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_B1 (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_S0 (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_A3 (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_A1 (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_A0 (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_A1 (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_A1 (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c222_S1 (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c220_A3 (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone8_A2 (.DIODE(net1098));
 sky130_fd_sc_hd__diode_2 ANTENNA_c138_A2 (.DIODE(net1098));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout212_X (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_A0 (.DIODE(net1098));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_A0 (.DIODE(net1098));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_A0 (.DIODE(net1098));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout213_X (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c530_D1 (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_A1 (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c401_A1 (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_A2 (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_A1 (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_A3 (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_A3 (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_A1 (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_A2 (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_A3 (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1_A (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone8_C1 (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone4_S1 (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout214_X (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c140_S1 (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout216_X (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_C1 (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_A1 (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_S0 (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_A2 (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout215_A (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout217_X (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_A0 (.DIODE(net1089));
 sky130_fd_sc_hd__diode_2 ANTENNA_c662_A2 (.DIODE(net1089));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_S1 (.DIODE(net1089));
 sky130_fd_sc_hd__diode_2 ANTENNA_c532_SCE (.DIODE(net1089));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout216_A (.DIODE(net1089));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout2_A (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone8_D1 (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout218_X (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout219_X (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_A2 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_S1 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c424_S1 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_S0 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_S1 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_S0 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_S1 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_S1 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_S1 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_S1 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout220_X (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_S1 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_S0 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c346_S1 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_S1 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_output152_A (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_S1 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_S0 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_S1 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_S1 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_S1 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap221_X (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_S1 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_S0 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_S1 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_S1 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_S0 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c494_S1 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c346_A3 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout222_X (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_S1 (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_S1 (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c323_S0 (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_S1 (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_S0 (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_S1 (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_S1 (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c313_S1 (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c482_S0 (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_S1 (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout223_X (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c611_A1 (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_S1 (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_S0 (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_S1 (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_S1 (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_S1 (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout224_X (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c695_S0 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_S0 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_S0 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_A3 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_S0 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_S0 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_A2 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_S0 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_S1 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_S1 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout226_X (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c743_S0 (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c742_S1 (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_S0 (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c587_S0 (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_C1 (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_S0 (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c313_A3 (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout225_A (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_S0 (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout227_X (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_B1 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_D1 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_S1 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_S1 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_S1 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_S1 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_S0 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_A3 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_S1 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_S0 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout228_X (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_A2 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c136_D1 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_S0 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_C1 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_C1 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_A0 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_A2 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c215_A0 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c212_A2 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c206_A2 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout230_X (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_A1 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_A2 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_A1 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_A2 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c231_A2 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_A3 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c106_S0 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c104_S0 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c103_S1 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c494_A2 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c265_D1 (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_A2 (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout232_X (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_A2 (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_A3 (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_A2 (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_A1 (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_A1 (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c229_A3 (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_A2 (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c158_A2 (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout233_X (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c267_B1 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c264_D1 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_A3 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c134_C1 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c205_A3 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c118_D1 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c115_D1 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c113_D1 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c112_B1 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c110_D1 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout234_X (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c543_C1 (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_A1 (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c403_D1 (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c402_SCD (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_D1 (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c766_A3 (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c761_A3 (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_A2 (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_A1 (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_S0 (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout235_X (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c660_C1 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c668_A3 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c671_D1 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout234_A (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_S0 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout233_A (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout5_A (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone8_A1 (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout236_X (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_A2 (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout237_X (.DIODE(net1097));
 sky130_fd_sc_hd__diode_2 ANTENNA_c571_A3 (.DIODE(net1097));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_A1 (.DIODE(net1097));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_A1 (.DIODE(net1097));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_A3 (.DIODE(net1097));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_C_N (.DIODE(net1097));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout238_X (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_c535_B1 (.DIODE(net1096));
 sky130_fd_sc_hd__diode_2 ANTENNA_c532_SCD (.DIODE(net1096));
 sky130_fd_sc_hd__diode_2 ANTENNA_c427_A2 (.DIODE(net1096));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_A0 (.DIODE(net1096));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_S1 (.DIODE(net1096));
 sky130_fd_sc_hd__diode_2 ANTENNA_c140_S0 (.DIODE(net1096));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_A0 (.DIODE(net1096));
 sky130_fd_sc_hd__diode_2 ANTENNA_c134_D1 (.DIODE(net1096));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_C1 (.DIODE(net1096));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_B (.DIODE(net1096));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout240_X (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_A1 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c136_A1 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c257_A0 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_S0 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_A0 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_A2 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_C1 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c127_S0 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c124_S1 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c115_A1 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout241_X (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_c661_C1 (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_c536_D1 (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_c405_SCE (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_A2 (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout240_A (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout242_X (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_A1 (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_D1 (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_S0 (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_D_N (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_c112_D1 (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout243_X (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c286_S1 (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_A2 (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_A2 (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_SCD (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_A3 (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone31_A (.DIODE(net1095));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout244_X (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_A1 (.DIODE(net1095));
 sky130_fd_sc_hd__diode_2 ANTENNA_c531_B1 (.DIODE(net1095));
 sky130_fd_sc_hd__diode_2 ANTENNA_c530_C1 (.DIODE(net1095));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout242_A (.DIODE(net1095));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout243_A (.DIODE(net1095));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout245_X (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_A1 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_A3 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c215_S0 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_A2 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c184_A2 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c131_A3 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c129_S1 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c116_D1 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c112_C1 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c111_A2 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout246_X (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_A3 (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_S0 (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_A1 (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_A3 (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_A2 (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_S0 (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c221_A2 (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_S1 (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_A3 (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_A1 (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout247_X (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_A0 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_A3 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_A2 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_A1 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_A0 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_A2 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_S0 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c264_B1 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c237_A0 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_A3 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout4_A (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone6_A0 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout248_X (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout249_X (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_S1 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c556_A3 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_A1 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_A3 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_A2 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_A1 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_A1 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c286_A2 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_A2 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_A2 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout250_X (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c428_A2 (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_A2 (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_S1 (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_A3 (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c229_A0 (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_D1 (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c129_S0 (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c121_A3 (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c113_C1 (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c111_D1 (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout251_X (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_c768_S1 (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_A1 (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_c696_A2 (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_A2 (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_c687_S1 (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_A3 (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_A0 (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_c563_C1 (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout252_X (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_A3 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c313_A2 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_A2 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_A1 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c230_A1 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c226_A1 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c191_A2 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_C1 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c158_S1 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c105_S0 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout253_X (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_A1 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c555_A1 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_A1 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c424_A2 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_S0 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_A0 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c295_A3 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout255_X (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_S0 (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_c557_B1 (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_A2 (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_c400_SCD (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_c397_B1 (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_A3 (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_c271_S1 (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_A2 (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_c267_A2 (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_S1 (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout256_X (.DIODE(net1025));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_A3 (.DIODE(net1025));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_A0 (.DIODE(net1025));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_A2 (.DIODE(net1025));
 sky130_fd_sc_hd__diode_2 ANTENNA_c686_A0 (.DIODE(net1025));
 sky130_fd_sc_hd__diode_2 ANTENNA_c668_A0 (.DIODE(net1025));
 sky130_fd_sc_hd__diode_2 ANTENNA_c582_A3 (.DIODE(net1025));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_A1 (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout257_X (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_A2 (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_A0 (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c677_A2 (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_A0 (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_A0 (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c274_RESET_B (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_S1 (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c134_B1 (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_A1 (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout258_X (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c686_A3 (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c675_A2 (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c667_A0 (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c664_A1 (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c587_A0 (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_A2 (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c401_B1 (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_A2 (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_A0 (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c134_A1 (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout259_X (.DIODE(net1028));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_A2 (.DIODE(net1028));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_A0 (.DIODE(net1028));
 sky130_fd_sc_hd__diode_2 ANTENNA_c148_A3 (.DIODE(net1028));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_A0 (.DIODE(net1028));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_A1 (.DIODE(net1028));
 sky130_fd_sc_hd__diode_2 ANTENNA_c502_A2 (.DIODE(net1028));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_S0 (.DIODE(net1028));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_S0 (.DIODE(net1028));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_S0 (.DIODE(net1028));
 sky130_fd_sc_hd__diode_2 ANTENNA_c215_A2 (.DIODE(net1028));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_B1 (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout260_X (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_A3 (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_A3 (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_A2 (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_c270_D1 (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_c266_A0 (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_c260_A0 (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_B1 (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_c119_A1 (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_c116_C1 (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_15_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_14_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_13_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_12_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_11_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_10_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_9_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_8_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_7_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_6_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_5_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_4_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_3_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_2_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_1_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_0_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_X (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c239_CLK_N (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge794_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge830_GATE (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge833_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge849_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge871_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge884_GATE_N (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s895_GATE_N (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s899_GATE_N (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s900_GATE_N (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s921_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s923_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_0_0_clk_X (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge797_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge799_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge829_GATE (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge870_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s893_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s896_GATE_N (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s897_GATE (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s898_GATE_N (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s916_GATE_N (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_1_0_clk_X (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge832_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge851_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge860_GATE (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge862_GATE_N (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge867_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge868_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge880_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge882_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s920_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s948_GATE_N (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s950_SLEEP_B (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_2_0_clk_X (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge835_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge861_GATE_N (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s917_GATE (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s918_SLEEP_B (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s919_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s922_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s941_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s942_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s944_GATE_N (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s946_GATE_N (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s949_GATE (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_3_0_clk_X (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c273_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c274_CLK_N (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c402_CLK_N (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge801_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge840_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s901_GATE (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s902_SLEEP_B (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s903_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s905_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s906_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s907_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s910_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_7_0_clk_X (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge795_CLK_N (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge838_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge842_CLK_N (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge853_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge864_GATE (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge877_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s947_GATE_N (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s951_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s961_GATE (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s962_GATE_N (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s963_GATE_N (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_8_0_clk_X (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c560_CLK_N (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge863_GATE_N (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s913_GATE (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s938_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s939_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s940_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s943_GATE_N (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s945_GATE (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s956_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s960_GATE_N (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_9_0_clk_X (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge850_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge856_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge857_GATE_N (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge866_GATE (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge874_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge875_CLK_N (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge876_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge878_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s959_GATE_N (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_10_0_clk_X (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge824_GATE_N (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge827_GATE (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge844_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge858_GATE_N (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge886_GATE (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s955_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s957_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s958_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s971_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_11_0_clk_X (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c398_CLK_N (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c562_CLK_N (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge814_GATE (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge826_GATE_N (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s928_GATE_N (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s930_GATE_N (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s931_GATE_N (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s932_GATE_N (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s934_SLEEP_B (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s935_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s936_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s937_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s954_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_12_0_clk_X (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c272_CLK_N (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c400_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c405_CLK_N (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c409_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c410_CLK_N (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c411_CLK_N (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c413_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c529_CLK_N (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c533_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c534_CLK_N (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge813_GATE_N (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s904_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s924_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s925_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s926_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s927_GATE_N (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s952_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_13_0_clk_X (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c548_CLK_N (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge796_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge798_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge837_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge839_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge859_GATE (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge879_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s967_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s968_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s969_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s970_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_14_0_clk_X (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c532_CLK_N (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c538_CLK_N (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c540_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c541_CLK_N (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge804_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge805_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge818_GATE (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge869_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge873_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge881_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge883_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s953_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s964_GATE_N (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s965_GATE (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s966_SLEEP_B (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_15_0_clk_X (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_A1 (.DIODE(clknet_1_0__leaf_net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_A2 (.DIODE(clknet_1_0__leaf_net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_A3 (.DIODE(clknet_1_0__leaf_net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_S0 (.DIODE(clknet_1_0__leaf_net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net939_X (.DIODE(clknet_1_0__leaf_net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_A2 (.DIODE(clknet_1_0__leaf_net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_A2 (.DIODE(clknet_1_0__leaf_net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_A0 (.DIODE(clknet_1_0__leaf_net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_A1 (.DIODE(clknet_1_0__leaf_net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_A2 (.DIODE(clknet_1_0__leaf_net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_A3 (.DIODE(clknet_1_0__leaf_net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_A1 (.DIODE(clknet_1_0__leaf_net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net904_X (.DIODE(clknet_1_0__leaf_net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_A1 (.DIODE(clknet_1_1__leaf_net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_A3 (.DIODE(clknet_1_1__leaf_net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_A3 (.DIODE(clknet_1_1__leaf_net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_output135_A (.DIODE(clknet_1_1__leaf_net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net904_X (.DIODE(clknet_1_1__leaf_net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net893_A (.DIODE(clknet_0_net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net893_A (.DIODE(clknet_0_net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net893_X (.DIODE(clknet_0_net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_A2 (.DIODE(clknet_1_0__leaf_net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_A2 (.DIODE(clknet_1_0__leaf_net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_S0 (.DIODE(clknet_1_0__leaf_net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_S0 (.DIODE(clknet_1_0__leaf_net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net893_X (.DIODE(clknet_1_0__leaf_net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_A1 (.DIODE(clknet_1_1__leaf_net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c528_A1 (.DIODE(clknet_1_1__leaf_net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_A2 (.DIODE(clknet_1_1__leaf_net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_output124_A (.DIODE(clknet_1_1__leaf_net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net893_X (.DIODE(clknet_1_1__leaf_net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net713_A (.DIODE(clknet_0_net713));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net713_A (.DIODE(clknet_0_net713));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net713_X (.DIODE(clknet_0_net713));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_A3 (.DIODE(clknet_1_0__leaf_net713));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_S0 (.DIODE(clknet_1_0__leaf_net713));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_S0 (.DIODE(clknet_1_0__leaf_net713));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_A3 (.DIODE(clknet_1_0__leaf_net713));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_S1 (.DIODE(clknet_1_0__leaf_net713));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_A2 (.DIODE(clknet_1_0__leaf_net713));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_S0 (.DIODE(clknet_1_0__leaf_net713));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net713_X (.DIODE(clknet_1_0__leaf_net713));
 sky130_fd_sc_hd__diode_2 ANTENNA_c434_A3 (.DIODE(clknet_1_0__leaf_net277));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_A2 (.DIODE(clknet_1_0__leaf_net277));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_A0 (.DIODE(clknet_1_0__leaf_net277));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net277_X (.DIODE(clknet_1_0__leaf_net277));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_A2 (.DIODE(clknet_1_0__leaf_net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_A2 (.DIODE(clknet_1_0__leaf_net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_A2 (.DIODE(clknet_1_0__leaf_net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net898_X (.DIODE(clknet_1_0__leaf_net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_A2 (.DIODE(clknet_1_1__leaf_net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c437_A2 (.DIODE(clknet_1_1__leaf_net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_output129_A (.DIODE(clknet_1_1__leaf_net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net898_X (.DIODE(clknet_1_1__leaf_net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c406_D1 (.DIODE(clknet_1_0__leaf_net712));
 sky130_fd_sc_hd__diode_2 ANTENNA_c407_D1 (.DIODE(clknet_1_0__leaf_net712));
 sky130_fd_sc_hd__diode_2 ANTENNA_c408_S1 (.DIODE(clknet_1_0__leaf_net712));
 sky130_fd_sc_hd__diode_2 ANTENNA_c410_SCE (.DIODE(clknet_1_0__leaf_net712));
 sky130_fd_sc_hd__diode_2 ANTENNA_c413_SET_B (.DIODE(clknet_1_0__leaf_net712));
 sky130_fd_sc_hd__diode_2 ANTENNA_c415_S0 (.DIODE(clknet_1_0__leaf_net712));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_S0 (.DIODE(clknet_1_0__leaf_net712));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_A3 (.DIODE(clknet_1_0__leaf_net712));
 sky130_fd_sc_hd__diode_2 ANTENNA_c531_D1 (.DIODE(clknet_1_0__leaf_net712));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net712_X (.DIODE(clknet_1_0__leaf_net712));
 sky130_fd_sc_hd__diode_2 ANTENNA_c534_SET_B (.DIODE(clknet_1_1__leaf_net712));
 sky130_fd_sc_hd__diode_2 ANTENNA_c667_S1 (.DIODE(clknet_1_1__leaf_net712));
 sky130_fd_sc_hd__diode_2 ANTENNA_c669_D1 (.DIODE(clknet_1_1__leaf_net712));
 sky130_fd_sc_hd__diode_2 ANTENNA_c681_S1 (.DIODE(clknet_1_1__leaf_net712));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_S0 (.DIODE(clknet_1_1__leaf_net712));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_A3 (.DIODE(clknet_1_1__leaf_net712));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_S1 (.DIODE(clknet_1_1__leaf_net712));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net712_X (.DIODE(clknet_1_1__leaf_net712));
 sky130_fd_sc_hd__diode_2 ANTENNA_c409_SCD (.DIODE(clknet_1_0__leaf_net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c430_A1 (.DIODE(clknet_1_0__leaf_net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c528_A2 (.DIODE(clknet_1_0__leaf_net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c534_SCD (.DIODE(clknet_1_0__leaf_net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_A1 (.DIODE(clknet_1_0__leaf_net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net247_X (.DIODE(clknet_1_0__leaf_net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c674_A1 (.DIODE(clknet_1_1__leaf_net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c695_A2 (.DIODE(clknet_1_1__leaf_net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c723_A1 (.DIODE(clknet_1_1__leaf_net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_A3 (.DIODE(clknet_1_1__leaf_net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c739_A3 (.DIODE(clknet_1_1__leaf_net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c761_A0 (.DIODE(clknet_1_1__leaf_net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net247_X (.DIODE(clknet_1_1__leaf_net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_S0 (.DIODE(clknet_1_1__leaf_net695));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_A3 (.DIODE(clknet_1_1__leaf_net695));
 sky130_fd_sc_hd__diode_2 ANTENNA_c555_A2 (.DIODE(clknet_1_1__leaf_net695));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_S0 (.DIODE(clknet_1_1__leaf_net695));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net695_X (.DIODE(clknet_1_1__leaf_net695));
 sky130_fd_sc_hd__diode_2 ANTENNA_c446_A3 (.DIODE(clknet_1_0__leaf_net263));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_A0 (.DIODE(clknet_1_0__leaf_net263));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net263_X (.DIODE(clknet_1_0__leaf_net263));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_A0 (.DIODE(clknet_1_0__leaf_net166));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_A2 (.DIODE(clknet_1_0__leaf_net166));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_A0 (.DIODE(clknet_1_0__leaf_net166));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net166_X (.DIODE(clknet_1_0__leaf_net166));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_S1 (.DIODE(clknet_1_0__leaf_net694));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_S0 (.DIODE(clknet_1_0__leaf_net694));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_S0 (.DIODE(clknet_1_0__leaf_net694));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_S0 (.DIODE(clknet_1_0__leaf_net694));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_S1 (.DIODE(clknet_1_0__leaf_net694));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_S0 (.DIODE(clknet_1_0__leaf_net694));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net694_X (.DIODE(clknet_1_0__leaf_net694));
 sky130_fd_sc_hd__diode_2 ANTENNA_c577_S1 (.DIODE(clknet_1_1__leaf_net694));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_S0 (.DIODE(clknet_1_1__leaf_net694));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_S0 (.DIODE(clknet_1_1__leaf_net694));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net694_X (.DIODE(clknet_1_1__leaf_net694));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_A2 (.DIODE(clknet_1_0__leaf_net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_A0 (.DIODE(clknet_1_0__leaf_net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net935_X (.DIODE(clknet_1_0__leaf_net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_SCE (.DIODE(clknet_1_1__leaf_net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_output166_A (.DIODE(clknet_1_1__leaf_net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net935_X (.DIODE(clknet_1_1__leaf_net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net693_A (.DIODE(clknet_0_net693));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net693_A (.DIODE(clknet_0_net693));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net693_X (.DIODE(clknet_0_net693));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_S1 (.DIODE(clknet_1_0__leaf_net693));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_S1 (.DIODE(clknet_1_0__leaf_net693));
 sky130_fd_sc_hd__diode_2 ANTENNA_c297_S1 (.DIODE(clknet_1_0__leaf_net693));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_S0 (.DIODE(clknet_1_0__leaf_net693));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_A3 (.DIODE(clknet_1_0__leaf_net693));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_A3 (.DIODE(clknet_1_0__leaf_net693));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_A3 (.DIODE(clknet_1_0__leaf_net693));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_S0 (.DIODE(clknet_1_0__leaf_net693));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_A3 (.DIODE(clknet_1_0__leaf_net693));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net693_X (.DIODE(clknet_1_0__leaf_net693));
 sky130_fd_sc_hd__diode_2 ANTENNA_c364_S0 (.DIODE(clknet_1_1__leaf_net693));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_A3 (.DIODE(clknet_1_1__leaf_net693));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_S1 (.DIODE(clknet_1_1__leaf_net693));
 sky130_fd_sc_hd__diode_2 ANTENNA_c693_A3 (.DIODE(clknet_1_1__leaf_net693));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_S0 (.DIODE(clknet_1_1__leaf_net693));
 sky130_fd_sc_hd__diode_2 ANTENNA_c762_S0 (.DIODE(clknet_1_1__leaf_net693));
 sky130_fd_sc_hd__diode_2 ANTENNA_c763_S1 (.DIODE(clknet_1_1__leaf_net693));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net693_X (.DIODE(clknet_1_1__leaf_net693));
 sky130_fd_sc_hd__diode_2 ANTENNA_c295_S0 (.DIODE(clknet_1_0__leaf_net157));
 sky130_fd_sc_hd__diode_2 ANTENNA_c430_A3 (.DIODE(clknet_1_0__leaf_net157));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_A2 (.DIODE(clknet_1_0__leaf_net157));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_A0 (.DIODE(clknet_1_0__leaf_net157));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net157_X (.DIODE(clknet_1_0__leaf_net157));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net900_A (.DIODE(clknet_0_net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net900_A (.DIODE(clknet_0_net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net900_X (.DIODE(clknet_0_net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_S0 (.DIODE(clknet_1_0__leaf_net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_A1 (.DIODE(clknet_1_0__leaf_net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_A2 (.DIODE(clknet_1_0__leaf_net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_A3 (.DIODE(clknet_1_0__leaf_net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_output131_A (.DIODE(clknet_1_0__leaf_net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net900_X (.DIODE(clknet_1_0__leaf_net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_A0 (.DIODE(clknet_1_1__leaf_net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_A1 (.DIODE(clknet_1_1__leaf_net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_A1 (.DIODE(clknet_1_1__leaf_net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_A1 (.DIODE(clknet_1_1__leaf_net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_A2 (.DIODE(clknet_1_1__leaf_net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_A3 (.DIODE(clknet_1_1__leaf_net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net900_X (.DIODE(clknet_1_1__leaf_net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net675_A (.DIODE(clknet_0_net675));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net675_A (.DIODE(clknet_0_net675));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net675_X (.DIODE(clknet_0_net675));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_S1 (.DIODE(clknet_1_0__leaf_net675));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_A3 (.DIODE(clknet_1_0__leaf_net675));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_A3 (.DIODE(clknet_1_0__leaf_net675));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_A3 (.DIODE(clknet_1_0__leaf_net675));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net675_X (.DIODE(clknet_1_0__leaf_net675));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_S0 (.DIODE(clknet_1_1__leaf_net675));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_S1 (.DIODE(clknet_1_1__leaf_net675));
 sky130_fd_sc_hd__diode_2 ANTENNA_c744_S0 (.DIODE(clknet_1_1__leaf_net675));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_S1 (.DIODE(clknet_1_1__leaf_net675));
 sky130_fd_sc_hd__diode_2 ANTENNA_c761_S1 (.DIODE(clknet_1_1__leaf_net675));
 sky130_fd_sc_hd__diode_2 ANTENNA_c762_A2 (.DIODE(clknet_1_1__leaf_net675));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net675_X (.DIODE(clknet_1_1__leaf_net675));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_S1 (.DIODE(clknet_1_0__leaf_net674));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_S1 (.DIODE(clknet_1_0__leaf_net674));
 sky130_fd_sc_hd__diode_2 ANTENNA_c215_S1 (.DIODE(clknet_1_0__leaf_net674));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_S0 (.DIODE(clknet_1_0__leaf_net674));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net674_X (.DIODE(clknet_1_0__leaf_net674));
 sky130_fd_sc_hd__diode_2 ANTENNA_c371_A1 (.DIODE(clknet_1_0__leaf_net199));
 sky130_fd_sc_hd__diode_2 ANTENNA_c769_A1 (.DIODE(clknet_1_0__leaf_net199));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net199_X (.DIODE(clknet_1_0__leaf_net199));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_A2 (.DIODE(clknet_1_1__leaf_net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A0 (.DIODE(clknet_1_1__leaf_net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net100_X (.DIODE(clknet_1_1__leaf_net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net73_A (.DIODE(clknet_0_net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net73_A (.DIODE(clknet_0_net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net73_X (.DIODE(clknet_0_net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_A2 (.DIODE(clknet_1_0__leaf_net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_c205_A2 (.DIODE(clknet_1_0__leaf_net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_A1 (.DIODE(clknet_1_0__leaf_net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net73_X (.DIODE(clknet_1_0__leaf_net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_SCD (.DIODE(clknet_1_0__leaf_net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_c208_A3 (.DIODE(clknet_1_0__leaf_net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_A1 (.DIODE(clknet_1_0__leaf_net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_A1 (.DIODE(clknet_1_0__leaf_net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_A3 (.DIODE(clknet_1_0__leaf_net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_A1 (.DIODE(clknet_1_0__leaf_net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net84_X (.DIODE(clknet_1_0__leaf_net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_c228_C1 (.DIODE(clknet_1_0__leaf_net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_c229_S1 (.DIODE(clknet_1_0__leaf_net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_A2 (.DIODE(clknet_1_0__leaf_net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net938_X (.DIODE(clknet_1_0__leaf_net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_RESET_B (.DIODE(clknet_1_1__leaf_net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_A2 (.DIODE(clknet_1_1__leaf_net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_c761_A2 (.DIODE(clknet_1_1__leaf_net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net83_X (.DIODE(clknet_1_1__leaf_net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_A1 (.DIODE(clknet_1_1__leaf_net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c226_A3 (.DIODE(clknet_1_1__leaf_net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c256_A1 (.DIODE(clknet_1_1__leaf_net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_output167_A (.DIODE(clknet_1_1__leaf_net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net936_X (.DIODE(clknet_1_1__leaf_net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c216_A0 (.DIODE(clknet_1_0__leaf_net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_c220_A2 (.DIODE(clknet_1_0__leaf_net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_A3 (.DIODE(clknet_1_0__leaf_net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_A3 (.DIODE(clknet_1_0__leaf_net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_A0 (.DIODE(clknet_1_0__leaf_net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net79_X (.DIODE(clknet_1_0__leaf_net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_A2 (.DIODE(clknet_1_1__leaf_net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_A3 (.DIODE(clknet_1_1__leaf_net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_A0 (.DIODE(clknet_1_1__leaf_net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_A0 (.DIODE(clknet_1_1__leaf_net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net79_X (.DIODE(clknet_1_1__leaf_net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_A1 (.DIODE(clknet_1_0__leaf_net70));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_A0 (.DIODE(clknet_1_0__leaf_net70));
 sky130_fd_sc_hd__diode_2 ANTENNA_c240_A3 (.DIODE(clknet_1_0__leaf_net70));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net70_X (.DIODE(clknet_1_0__leaf_net70));
 sky130_fd_sc_hd__diode_2 ANTENNA_c190_A1 (.DIODE(clknet_1_1__leaf_net70));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_A1 (.DIODE(clknet_1_1__leaf_net70));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_A0 (.DIODE(clknet_1_1__leaf_net70));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net70_X (.DIODE(clknet_1_1__leaf_net70));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_A1 (.DIODE(clknet_1_0__leaf_net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_A0 (.DIODE(clknet_1_0__leaf_net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net74_X (.DIODE(clknet_1_0__leaf_net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_c191_A1 (.DIODE(clknet_1_0__leaf_net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_A1 (.DIODE(clknet_1_0__leaf_net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net72_X (.DIODE(clknet_1_0__leaf_net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_A2 (.DIODE(clknet_1_1__leaf_net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_c344_A2 (.DIODE(clknet_1_1__leaf_net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_c446_A0 (.DIODE(clknet_1_1__leaf_net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net72_X (.DIODE(clknet_1_1__leaf_net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_A1 (.DIODE(clknet_1_0__leaf_net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_A2 (.DIODE(clknet_1_0__leaf_net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_A1 (.DIODE(clknet_1_0__leaf_net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_c371_A0 (.DIODE(clknet_1_0__leaf_net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net75_X (.DIODE(clknet_1_0__leaf_net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_A2 (.DIODE(clknet_1_1__leaf_net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_c194_A2 (.DIODE(clknet_1_1__leaf_net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_A1 (.DIODE(clknet_1_1__leaf_net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net75_X (.DIODE(clknet_1_1__leaf_net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_A2 (.DIODE(clknet_1_0__leaf_net288));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_A1 (.DIODE(clknet_1_0__leaf_net288));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_A3 (.DIODE(clknet_1_0__leaf_net288));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_A0 (.DIODE(clknet_1_0__leaf_net288));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net288_X (.DIODE(clknet_1_0__leaf_net288));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net673_A (.DIODE(clknet_0_net673));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net673_A (.DIODE(clknet_0_net673));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net673_X (.DIODE(clknet_0_net673));
 sky130_fd_sc_hd__diode_2 ANTENNA_c182_S1 (.DIODE(clknet_1_0__leaf_net673));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_S0 (.DIODE(clknet_1_0__leaf_net673));
 sky130_fd_sc_hd__diode_2 ANTENNA_c191_S1 (.DIODE(clknet_1_0__leaf_net673));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_S1 (.DIODE(clknet_1_0__leaf_net673));
 sky130_fd_sc_hd__diode_2 ANTENNA_c194_S1 (.DIODE(clknet_1_0__leaf_net673));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_S1 (.DIODE(clknet_1_0__leaf_net673));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net673_X (.DIODE(clknet_1_0__leaf_net673));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer2_A (.DIODE(net1030));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_A3 (.DIODE(net1030));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer1_X (.DIODE(net1030));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer3_A (.DIODE(net1033));
 sky130_fd_sc_hd__diode_2 ANTENNA_c667_A1 (.DIODE(net1033));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_A1 (.DIODE(net1033));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_A2 (.DIODE(net1033));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone4_X (.DIODE(net1033));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone4_A2 (.DIODE(net1034));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer5_X (.DIODE(net1034));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_A1 (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_A3 (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_A3 (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer5_A (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_A3 (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone6_X (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout207_A (.DIODE(net1036));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer7_X (.DIODE(net1036));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_A1 (.DIODE(net1037));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_A1 (.DIODE(net1037));
 sky130_fd_sc_hd__diode_2 ANTENNA_c660_A1 (.DIODE(net1037));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone4_A3 (.DIODE(net1037));
 sky130_fd_sc_hd__diode_2 ANTENNA_c669_B1 (.DIODE(net1037));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone8_X (.DIODE(net1037));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout202_A (.DIODE(net1038));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer9_X (.DIODE(net1038));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_S0 (.DIODE(net1040));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer11_X (.DIODE(net1040));
 sky130_fd_sc_hd__diode_2 ANTENNA_c544_A2 (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_c558_A2 (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_c701_S0 (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_c663_B1 (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_A0 (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone12_X (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_A1 (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_A1 (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_A0 (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_c665_C1 (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_c398_SCE (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone13_X (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer14_A (.DIODE(net1044));
 sky130_fd_sc_hd__diode_2 ANTENNA_c402_D (.DIODE(net1044));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_A0 (.DIODE(net1044));
 sky130_fd_sc_hd__diode_2 ANTENNA_c431_A2 (.DIODE(net1044));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone15_X (.DIODE(net1044));
 sky130_fd_sc_hd__diode_2 ANTENNA_c428_A3 (.DIODE(net1049));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_A3 (.DIODE(net1049));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_A3 (.DIODE(net1049));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_A2 (.DIODE(net1049));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_A3 (.DIODE(net1049));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone20_X (.DIODE(net1049));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer23_A (.DIODE(net1051));
 sky130_fd_sc_hd__diode_2 ANTENNA_c538_SCE (.DIODE(net1051));
 sky130_fd_sc_hd__diode_2 ANTENNA_c411_SCE (.DIODE(net1051));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer22_X (.DIODE(net1051));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_S0 (.DIODE(net1054));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_A3 (.DIODE(net1054));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_A0 (.DIODE(net1054));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer17_A (.DIODE(net1054));
 sky130_fd_sc_hd__diode_2 ANTENNA_c370_A2 (.DIODE(net1054));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone25_X (.DIODE(net1054));
 sky130_fd_sc_hd__diode_2 ANTENNA_c143_A3 (.DIODE(net1057));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_A2 (.DIODE(net1057));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_A3 (.DIODE(net1057));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_A1 (.DIODE(net1057));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone6_A3 (.DIODE(net1057));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone28_X (.DIODE(net1057));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_A2 (.DIODE(net1058));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer30_A (.DIODE(net1058));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_A1 (.DIODE(net1058));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_A1 (.DIODE(net1058));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer29_X (.DIODE(net1058));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_B1 (.DIODE(net1060));
 sky130_fd_sc_hd__diode_2 ANTENNA_c110_C1 (.DIODE(net1060));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_A0 (.DIODE(net1060));
 sky130_fd_sc_hd__diode_2 ANTENNA_c125_B1 (.DIODE(net1060));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_A0 (.DIODE(net1060));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone31_X (.DIODE(net1060));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_A3 (.DIODE(net1062));
 sky130_fd_sc_hd__diode_2 ANTENNA_c757_A2 (.DIODE(net1062));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer33_X (.DIODE(net1062));
 sky130_fd_sc_hd__diode_2 ANTENNA_c403_A2 (.DIODE(net1063));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_A1 (.DIODE(net1063));
 sky130_fd_sc_hd__diode_2 ANTENNA_c311_A1 (.DIODE(net1063));
 sky130_fd_sc_hd__diode_2 ANTENNA_c278_S0 (.DIODE(net1063));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_A1 (.DIODE(net1063));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone34_X (.DIODE(net1063));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1_X (.DIODE(net1079));
 sky130_fd_sc_hd__diode_2 ANTENNA_c136_B1 (.DIODE(net1079));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_A3 (.DIODE(net1079));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_D1 (.DIODE(net1079));
 sky130_fd_sc_hd__diode_2 ANTENNA_c138_C1 (.DIODE(net1079));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_S1 (.DIODE(net1079));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_C1 (.DIODE(net1079));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_S1 (.DIODE(net1079));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_S1 (.DIODE(net1079));
 sky130_fd_sc_hd__diode_2 ANTENNA_c143_S1 (.DIODE(net1079));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone6_S1 (.DIODE(net1079));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout2_X (.DIODE(net1080));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_C1 (.DIODE(net1080));
 sky130_fd_sc_hd__diode_2 ANTENNA_c138_D1 (.DIODE(net1080));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_A1 (.DIODE(net1080));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_S0 (.DIODE(net1080));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_A0 (.DIODE(net1080));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_A1 (.DIODE(net1080));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_A2 (.DIODE(net1080));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_A3 (.DIODE(net1080));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_A1 (.DIODE(net1080));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_A2 (.DIODE(net1080));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout3_X (.DIODE(net1081));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_A2 (.DIODE(net1081));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_A1 (.DIODE(net1081));
 sky130_fd_sc_hd__diode_2 ANTENNA_c611_A0 (.DIODE(net1081));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_S0 (.DIODE(net1081));
 sky130_fd_sc_hd__diode_2 ANTENNA_c277_A2 (.DIODE(net1081));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_D (.DIODE(net1081));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_B1 (.DIODE(net1081));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_A1 (.DIODE(net1081));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_A3 (.DIODE(net1081));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_A2 (.DIODE(net1081));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout4_X (.DIODE(net1082));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_C1 (.DIODE(net1082));
 sky130_fd_sc_hd__diode_2 ANTENNA_c143_A0 (.DIODE(net1082));
 sky130_fd_sc_hd__diode_2 ANTENNA_c140_A1 (.DIODE(net1082));
 sky130_fd_sc_hd__diode_2 ANTENNA_c494_S0 (.DIODE(net1082));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_A2 (.DIODE(net1082));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_A1 (.DIODE(net1082));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_A1 (.DIODE(net1082));
 sky130_fd_sc_hd__diode_2 ANTENNA_c203_C1 (.DIODE(net1082));
 sky130_fd_sc_hd__diode_2 ANTENNA_c107_A2 (.DIODE(net1082));
 sky130_fd_sc_hd__diode_2 ANTENNA_c101_A3 (.DIODE(net1082));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout5_X (.DIODE(net1083));
 sky130_fd_sc_hd__diode_2 ANTENNA_c666_B1 (.DIODE(net1083));
 sky130_fd_sc_hd__diode_2 ANTENNA_c404_A1 (.DIODE(net1083));
 sky130_fd_sc_hd__diode_2 ANTENNA_c138_A1 (.DIODE(net1083));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone6_A2 (.DIODE(net1083));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_A3 (.DIODE(net1083));
 sky130_fd_sc_hd__diode_2 ANTENNA_c183_A0 (.DIODE(net1083));
 sky130_fd_sc_hd__diode_2 ANTENNA_c159_B1 (.DIODE(net1083));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_S0 (.DIODE(net1083));
 sky130_fd_sc_hd__diode_2 ANTENNA_c143_A2 (.DIODE(net1083));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_A2 (.DIODE(net1083));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout6_X (.DIODE(net1084));
 sky130_fd_sc_hd__diode_2 ANTENNA_c407_A1 (.DIODE(net1084));
 sky130_fd_sc_hd__diode_2 ANTENNA_c404_S0 (.DIODE(net1084));
 sky130_fd_sc_hd__diode_2 ANTENNA_c266_A2 (.DIODE(net1084));
 sky130_fd_sc_hd__diode_2 ANTENNA_c265_B1 (.DIODE(net1084));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_A3 (.DIODE(net1084));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_A2 (.DIODE(net1084));
 sky130_fd_sc_hd__diode_2 ANTENNA_c140_A0 (.DIODE(net1084));
 sky130_fd_sc_hd__diode_2 ANTENNA_c138_B1 (.DIODE(net1084));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_A2 (.DIODE(net1084));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_A (.DIODE(net1084));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout7_X (.DIODE(net1085));
 sky130_fd_sc_hd__diode_2 ANTENNA_c412_A0 (.DIODE(net1085));
 sky130_fd_sc_hd__diode_2 ANTENNA_c401_C1 (.DIODE(net1085));
 sky130_fd_sc_hd__diode_2 ANTENNA_c399_C1 (.DIODE(net1085));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone6_A1 (.DIODE(net1085));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_A0 (.DIODE(net1085));
 sky130_fd_sc_hd__diode_2 ANTENNA_c277_A0 (.DIODE(net1085));
 sky130_fd_sc_hd__diode_2 ANTENNA_c275_S0 (.DIODE(net1085));
 sky130_fd_sc_hd__diode_2 ANTENNA_c269_A2 (.DIODE(net1085));
 sky130_fd_sc_hd__diode_2 ANTENNA_c148_A2 (.DIODE(net1085));
 sky130_fd_sc_hd__diode_2 ANTENNA_c143_A1 (.DIODE(net1085));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(net0));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(clknet_1_0__leaf_net73));
 sky130_fd_sc_hd__mux4_1 clone1 (.A0(net1082),
    .A1(net1085),
    .A2(net1083),
    .A3(net1057),
    .S0(net27),
    .S1(net1079),
    .X(net1086));
 sky130_fd_sc_hd__mux4_1 clone2 (.A0(net998),
    .A1(net26),
    .A2(net19),
    .A3(net1006),
    .S0(net24),
    .S1(net984),
    .X(net1087));
 sky130_fd_sc_hd__a2111o_1 clone3 (.A1(net31),
    .A2(net1001),
    .B1(net1081),
    .C1(net1094),
    .D1(net1079),
    .X(net1088));
 sky130_fd_sc_hd__clkbuf_1 clone5 (.A(net21),
    .X(net1089));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer6 (.A(net23),
    .X(net1090));
 sky130_fd_sc_hd__a2111o_1 clone7 (.A1(net1057),
    .A2(net1024),
    .B1(net124),
    .C1(net969),
    .D1(net964),
    .X(net1091));
 sky130_fd_sc_hd__clkbuf_1 clone9 (.A(net872),
    .X(net1092));
 sky130_fd_sc_hd__clkbuf_1 clone10 (.A(net34),
    .X(net1093));
 sky130_fd_sc_hd__clkbuf_1 clone11 (.A(net872),
    .X(net1094));
 sky130_fd_sc_hd__clkbuf_1 clone14 (.A(net815),
    .X(net1095));
 sky130_fd_sc_hd__clkbuf_1 clone16 (.A(net826),
    .X(net1096));
 sky130_fd_sc_hd__clkbuf_1 clone17 (.A(net776),
    .X(net1097));
 sky130_fd_sc_hd__clkbuf_1 clone18 (.A(net23),
    .X(net1098));
 sky130_fd_sc_hd__a2111o_1 clone19 (.A1(net984),
    .A2(net1026),
    .B1(net998),
    .C1(net1080),
    .D1(net1011),
    .X(net1099));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(net762),
    .X(net1108));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_413 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_5 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_103 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_19 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_191 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_256 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_423 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_230 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_90 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_245 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_71 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_130 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_366 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_452 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_6 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_143 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_163 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_452 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_479 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_546 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_471 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_469 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_275 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_67 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_102 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_480 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_422 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_198 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_443 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_59 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_143 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_163 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_497 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_539 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_423 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_510 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_525 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_168 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_226 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_10 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_186 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_395 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_497 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_412 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_487 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_171 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_441 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_5 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_163 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_525 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_115 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_146 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_310 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_525 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_448 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_507 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_227 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_407 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_270 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_10 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_525 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_403 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_440 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_5 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_395 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_499 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_511 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_5 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_546 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_480 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_5 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_10 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_617 ();
endmodule
