module netlist_1 (clk,
    in0,
    in1,
    in10,
    in11,
    in12,
    in13,
    in14,
    in15,
    in16,
    in17,
    in18,
    in19,
    in2,
    in20,
    in21,
    in22,
    in23,
    in24,
    in25,
    in26,
    in27,
    in28,
    in29,
    in3,
    in30,
    in31,
    in32,
    in33,
    in34,
    in35,
    in36,
    in37,
    in38,
    in39,
    in4,
    in40,
    in41,
    in42,
    in43,
    in44,
    in45,
    in46,
    in47,
    in48,
    in49,
    in5,
    in50,
    in51,
    in52,
    in53,
    in54,
    in55,
    in56,
    in57,
    in58,
    in59,
    in6,
    in60,
    in61,
    in62,
    in63,
    in64,
    in65,
    in66,
    in67,
    in68,
    in69,
    in7,
    in70,
    in71,
    in72,
    in73,
    in74,
    in75,
    in76,
    in77,
    in78,
    in79,
    in8,
    in80,
    in81,
    in82,
    in83,
    in84,
    in85,
    in86,
    in87,
    in88,
    in89,
    in9,
    in90,
    in91,
    in92,
    in93,
    in94,
    in95,
    in96,
    in97,
    in98,
    in99,
    out0,
    out1,
    out10,
    out11,
    out12,
    out13,
    out14,
    out15,
    out16,
    out17,
    out18,
    out19,
    out2,
    out20,
    out21,
    out22,
    out23,
    out24,
    out25,
    out26,
    out27,
    out28,
    out29,
    out3,
    out30,
    out31,
    out32,
    out33,
    out34,
    out35,
    out36,
    out37,
    out38,
    out39,
    out4,
    out40,
    out41,
    out42,
    out43,
    out44,
    out45,
    out46,
    out47,
    out48,
    out49,
    out5,
    out50,
    out51,
    out52,
    out53,
    out54,
    out55,
    out56,
    out57,
    out58,
    out59,
    out6,
    out60,
    out61,
    out62,
    out63,
    out64,
    out65,
    out66,
    out67,
    out68,
    out69,
    out7,
    out70,
    out71,
    out72,
    out73,
    out74,
    out75,
    out76,
    out77,
    out78,
    out79,
    out8,
    out80,
    out81,
    out82,
    out83,
    out84,
    out85,
    out86,
    out87,
    out88,
    out89,
    out9,
    out90,
    out91,
    out92,
    out93,
    out94,
    out95,
    out96,
    out97,
    out98,
    out99,
    rst);
 input clk;
 input in0;
 input in1;
 input in10;
 input in11;
 input in12;
 input in13;
 input in14;
 input in15;
 input in16;
 input in17;
 input in18;
 input in19;
 input in2;
 input in20;
 input in21;
 input in22;
 input in23;
 input in24;
 input in25;
 input in26;
 input in27;
 input in28;
 input in29;
 input in3;
 input in30;
 input in31;
 input in32;
 input in33;
 input in34;
 input in35;
 input in36;
 input in37;
 input in38;
 input in39;
 input in4;
 input in40;
 input in41;
 input in42;
 input in43;
 input in44;
 input in45;
 input in46;
 input in47;
 input in48;
 input in49;
 input in5;
 input in50;
 input in51;
 input in52;
 input in53;
 input in54;
 input in55;
 input in56;
 input in57;
 input in58;
 input in59;
 input in6;
 input in60;
 input in61;
 input in62;
 input in63;
 input in64;
 input in65;
 input in66;
 input in67;
 input in68;
 input in69;
 input in7;
 input in70;
 input in71;
 input in72;
 input in73;
 input in74;
 input in75;
 input in76;
 input in77;
 input in78;
 input in79;
 input in8;
 input in80;
 input in81;
 input in82;
 input in83;
 input in84;
 input in85;
 input in86;
 input in87;
 input in88;
 input in89;
 input in9;
 input in90;
 input in91;
 input in92;
 input in93;
 input in94;
 input in95;
 input in96;
 input in97;
 input in98;
 input in99;
 output out0;
 output out1;
 output out10;
 output out11;
 output out12;
 output out13;
 output out14;
 output out15;
 output out16;
 output out17;
 output out18;
 output out19;
 output out2;
 output out20;
 output out21;
 output out22;
 output out23;
 output out24;
 output out25;
 output out26;
 output out27;
 output out28;
 output out29;
 output out3;
 output out30;
 output out31;
 output out32;
 output out33;
 output out34;
 output out35;
 output out36;
 output out37;
 output out38;
 output out39;
 output out4;
 output out40;
 output out41;
 output out42;
 output out43;
 output out44;
 output out45;
 output out46;
 output out47;
 output out48;
 output out49;
 output out5;
 output out50;
 output out51;
 output out52;
 output out53;
 output out54;
 output out55;
 output out56;
 output out57;
 output out58;
 output out59;
 output out6;
 output out60;
 output out61;
 output out62;
 output out63;
 output out64;
 output out65;
 output out66;
 output out67;
 output out68;
 output out69;
 output out7;
 output out70;
 output out71;
 output out72;
 output out73;
 output out74;
 output out75;
 output out76;
 output out77;
 output out78;
 output out79;
 output out8;
 output out80;
 output out81;
 output out82;
 output out83;
 output out84;
 output out85;
 output out86;
 output out87;
 output out88;
 output out89;
 output out9;
 output out90;
 output out91;
 output out92;
 output out93;
 output out94;
 output out95;
 output out96;
 output out97;
 output out98;
 output out99;
 input rst;

 wire net0;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net63;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net64;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net65;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net66;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net67;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net68;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net69;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net7;
 wire net70;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net71;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net72;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net73;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net74;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net75;
 wire net750;
 wire net751;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net194;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_0_net734;
 wire clknet_1_0__leaf_net734;
 wire clknet_1_1__leaf_net734;
 wire clknet_0_net733;
 wire clknet_1_0__leaf_net733;
 wire clknet_1_1__leaf_net733;
 wire clknet_0_net732;
 wire clknet_1_0__leaf_net732;
 wire clknet_1_1__leaf_net732;
 wire clknet_0_net429;
 wire clknet_1_0__leaf_net429;
 wire clknet_1_1__leaf_net429;
 wire clknet_0_net715;
 wire clknet_1_0__leaf_net715;
 wire clknet_1_1__leaf_net715;
 wire clknet_0_net380;
 wire clknet_1_0__leaf_net380;
 wire clknet_1_1__leaf_net380;
 wire clknet_0_net377;
 wire clknet_1_0__leaf_net377;
 wire clknet_1_1__leaf_net377;
 wire clknet_0_net375;
 wire clknet_1_0__leaf_net375;
 wire clknet_1_1__leaf_net375;
 wire clknet_0_net714;
 wire clknet_1_0__leaf_net714;
 wire clknet_1_1__leaf_net714;
 wire clknet_0_net407;
 wire clknet_1_0__leaf_net407;
 wire clknet_1_1__leaf_net407;
 wire clknet_0_net713;
 wire clknet_1_0__leaf_net713;
 wire clknet_1_1__leaf_net713;
 wire clknet_0_net372;
 wire clknet_1_0__leaf_net372;
 wire clknet_1_1__leaf_net372;
 wire clknet_0_net695;
 wire clknet_1_0__leaf_net695;
 wire clknet_1_1__leaf_net695;
 wire clknet_0_net310;
 wire clknet_1_0__leaf_net310;
 wire clknet_1_1__leaf_net310;
 wire clknet_0_net527;
 wire clknet_1_0__leaf_net527;
 wire clknet_1_1__leaf_net527;
 wire clknet_0_net694;
 wire clknet_1_0__leaf_net694;
 wire clknet_1_1__leaf_net694;
 wire clknet_0_net868;
 wire clknet_1_0__leaf_net868;
 wire clknet_1_1__leaf_net868;
 wire clknet_0_net302;
 wire clknet_1_0__leaf_net302;
 wire clknet_1_1__leaf_net302;
 wire clknet_0_net882;
 wire clknet_1_0__leaf_net882;
 wire clknet_1_1__leaf_net882;
 wire clknet_0_net693;
 wire clknet_1_0__leaf_net693;
 wire clknet_1_1__leaf_net693;
 wire clknet_0_net675;
 wire clknet_1_0__leaf_net675;
 wire clknet_1_1__leaf_net675;
 wire clknet_0_net913;
 wire clknet_1_0__leaf_net913;
 wire clknet_1_1__leaf_net913;
 wire clknet_0_net521;
 wire clknet_1_0__leaf_net521;
 wire clknet_1_1__leaf_net521;
 wire clknet_0_net495;
 wire clknet_1_0__leaf_net495;
 wire clknet_1_1__leaf_net495;
 wire clknet_0_net451;
 wire clknet_1_0__leaf_net451;
 wire clknet_1_1__leaf_net451;
 wire clknet_0_net469;
 wire clknet_1_0__leaf_net469;
 wire clknet_1_1__leaf_net469;
 wire clknet_0_net455;
 wire clknet_1_0__leaf_net455;
 wire clknet_1_1__leaf_net455;
 wire clknet_0_net499;
 wire clknet_1_0__leaf_net499;
 wire clknet_1_1__leaf_net499;
 wire clknet_0_net502;
 wire clknet_1_0__leaf_net502;
 wire clknet_1_1__leaf_net502;
 wire clknet_0_net489;
 wire clknet_1_0__leaf_net489;
 wire clknet_1_1__leaf_net489;
 wire clknet_0_net458;
 wire clknet_1_0__leaf_net458;
 wire clknet_1_1__leaf_net458;
 wire clknet_0_net457;
 wire clknet_1_0__leaf_net457;
 wire clknet_1_1__leaf_net457;
 wire clknet_0_net463;
 wire clknet_1_0__leaf_net463;
 wire clknet_1_1__leaf_net463;
 wire clknet_0_net250;
 wire clknet_1_0__leaf_net250;
 wire clknet_1_1__leaf_net250;
 wire clknet_0_net456;
 wire clknet_1_0__leaf_net456;
 wire clknet_1_1__leaf_net456;
 wire clknet_0_net446;
 wire clknet_1_0__leaf_net446;
 wire clknet_1_1__leaf_net446;
 wire clknet_0_net481;
 wire clknet_1_0__leaf_net481;
 wire clknet_1_1__leaf_net481;
 wire clknet_0_net447;
 wire clknet_1_0__leaf_net447;
 wire clknet_1_1__leaf_net447;
 wire clknet_0_net443;
 wire clknet_1_0__leaf_net443;
 wire clknet_1_1__leaf_net443;
 wire clknet_0_net349;
 wire clknet_1_0__leaf_net349;
 wire clknet_1_1__leaf_net349;
 wire clknet_0_net674;
 wire clknet_1_0__leaf_net674;
 wire clknet_1_1__leaf_net674;
 wire clknet_0_net352;
 wire clknet_1_0__leaf_net352;
 wire clknet_1_1__leaf_net352;
 wire clknet_0_net523;
 wire clknet_1_0__leaf_net523;
 wire clknet_1_1__leaf_net523;
 wire clknet_0_net643;
 wire clknet_1_0__leaf_net643;
 wire clknet_1_1__leaf_net643;
 wire clknet_0_net528;
 wire clknet_1_0__leaf_net528;
 wire clknet_1_1__leaf_net528;
 wire clknet_0_net877;
 wire clknet_1_0__leaf_net877;
 wire clknet_1_1__leaf_net877;
 wire clknet_0_net358;
 wire clknet_1_0__leaf_net358;
 wire clknet_1_1__leaf_net358;
 wire clknet_0_net492;
 wire clknet_1_0__leaf_net492;
 wire clknet_1_1__leaf_net492;
 wire clknet_0_net509;
 wire clknet_1_0__leaf_net509;
 wire clknet_1_1__leaf_net509;
 wire clknet_0_net357;
 wire clknet_1_0__leaf_net357;
 wire clknet_1_1__leaf_net357;
 wire clknet_0_net353;
 wire clknet_1_0__leaf_net353;
 wire clknet_1_1__leaf_net353;
 wire clknet_0_net348;
 wire clknet_1_0__leaf_net348;
 wire clknet_1_1__leaf_net348;
 wire clknet_0_net370;
 wire clknet_1_0__leaf_net370;
 wire clknet_1_1__leaf_net370;
 wire clknet_0_net403;
 wire clknet_1_0__leaf_net403;
 wire clknet_1_1__leaf_net403;
 wire clknet_0_net366;
 wire clknet_1_0__leaf_net366;
 wire clknet_1_1__leaf_net366;
 wire clknet_0_net342;
 wire clknet_1_0__leaf_net342;
 wire clknet_1_1__leaf_net342;
 wire clknet_0_net444;
 wire clknet_1_0__leaf_net444;
 wire clknet_1_1__leaf_net444;
 wire clknet_0_net347;
 wire clknet_1_0__leaf_net347;
 wire clknet_1_1__leaf_net347;
 wire clknet_0_net343;
 wire clknet_1_0__leaf_net343;
 wire clknet_1_1__leaf_net343;
 wire clknet_0_net246;
 wire clknet_1_0__leaf_net246;
 wire clknet_1_1__leaf_net246;
 wire clknet_0_net673;
 wire clknet_1_0__leaf_net673;
 wire clknet_1_1__leaf_net673;
 wire clknet_0_net341;
 wire clknet_1_0__leaf_net341;
 wire clknet_1_1__leaf_net341;
 wire clknet_0_net367;
 wire clknet_1_0__leaf_net367;
 wire clknet_1_1__leaf_net367;
 wire clknet_0_net658;
 wire clknet_1_0__leaf_net658;
 wire clknet_1_1__leaf_net658;
 wire clknet_0_net907;
 wire clknet_1_0__leaf_net907;
 wire clknet_1_1__leaf_net907;
 wire clknet_0_net107;
 wire clknet_1_0__leaf_net107;
 wire clknet_1_1__leaf_net107;
 wire clknet_0_net318;
 wire clknet_1_0__leaf_net318;
 wire clknet_1_1__leaf_net318;
 wire clknet_0_net205;
 wire clknet_1_0__leaf_net205;
 wire clknet_1_1__leaf_net205;
 wire clknet_0_net109;
 wire clknet_1_0__leaf_net109;
 wire clknet_1_1__leaf_net109;
 wire clknet_0_net105;
 wire clknet_1_0__leaf_net105;
 wire clknet_1_1__leaf_net105;
 wire clknet_0_net921;
 wire clknet_1_0__leaf_net921;
 wire clknet_1_1__leaf_net921;
 wire clknet_0_net657;
 wire clknet_1_0__leaf_net657;
 wire clknet_1_1__leaf_net657;
 wire clknet_0_net656;
 wire clknet_1_0__leaf_net656;
 wire clknet_1_1__leaf_net656;
 wire clknet_0_net316;
 wire clknet_1_0__leaf_net316;
 wire clknet_1_1__leaf_net316;
 wire clknet_0_net644;
 wire clknet_1_0__leaf_net644;
 wire clknet_1_1__leaf_net644;
 wire clknet_0_net216;
 wire clknet_1_0__leaf_net216;
 wire clknet_1_1__leaf_net216;
 wire clknet_0_net912;
 wire clknet_1_0__leaf_net912;
 wire clknet_1_1__leaf_net912;
 wire clknet_0_net887;
 wire clknet_1_0__leaf_net887;
 wire clknet_1_1__leaf_net887;
 wire clknet_0_net319;
 wire clknet_1_0__leaf_net319;
 wire clknet_1_1__leaf_net319;
 wire clknet_0_net203;
 wire clknet_1_0__leaf_net203;
 wire clknet_1_1__leaf_net203;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;

 sky130_fd_sc_hd__mux4_2 c100 (.A0(net841),
    .A1(net843),
    .A2(net838),
    .A3(net1025),
    .S0(net848),
    .S1(net819),
    .X(net0));
 sky130_fd_sc_hd__mux4_1 c101 (.A0(net835),
    .A1(net848),
    .A2(net843),
    .A3(net841),
    .S0(net842),
    .S1(net819),
    .X(net1));
 sky130_fd_sc_hd__mux4_2 c102 (.A0(net1021),
    .A1(net842),
    .A2(net843),
    .A3(net815),
    .S0(net833),
    .S1(net848),
    .X(net903));
 sky130_fd_sc_hd__mux4_2 c103 (.A0(net843),
    .A1(net835),
    .A2(net842),
    .A3(net848),
    .S0(net844),
    .S1(net801),
    .X(net925));
 sky130_fd_sc_hd__mux4_1 c104 (.A0(net1),
    .A1(net822),
    .A2(net838),
    .A3(net848),
    .S0(net834),
    .S1(net825),
    .X(net2));
 sky130_fd_sc_hd__mux4_2 c105 (.A0(net848),
    .A1(net843),
    .A2(net2),
    .A3(net842),
    .S0(net844),
    .S1(net1003),
    .X(net3));
 sky130_fd_sc_hd__mux4_1 c106 (.A0(net839),
    .A1(net844),
    .A2(net3),
    .A3(net822),
    .S0(net799),
    .S1(net1024),
    .X(net4));
 sky130_fd_sc_hd__mux4_2 c107 (.A0(net842),
    .A1(net4),
    .A2(net822),
    .A3(net841),
    .S0(net817),
    .S1(net848),
    .X(net890));
 sky130_fd_sc_hd__mux4_1 c108 (.A0(net2),
    .A1(net767),
    .A2(net849),
    .A3(net844),
    .S0(net821),
    .S1(net890),
    .X(net5));
 sky130_fd_sc_hd__mux4_2 c109 (.A0(net850),
    .A1(net822),
    .A2(net5),
    .A3(net3),
    .S0(net770),
    .S1(net890),
    .X(net905));
 sky130_fd_sc_hd__mux4_1 c110 (.A0(net1),
    .A1(net841),
    .A2(net804),
    .A3(net903),
    .S0(net801),
    .S1(net1014),
    .X(net6));
 sky130_fd_sc_hd__a41o_1 c111 (.A1(net776),
    .A2(net817),
    .A3(net805),
    .A4(net6),
    .B1(net994),
    .X(net7));
 sky130_fd_sc_hd__a41o_1 c112 (.A1(net801),
    .A2(net828),
    .A3(net770),
    .A4(net1),
    .B1(net1014),
    .X(net8));
 sky130_fd_sc_hd__a41o_2 c113 (.A1(net839),
    .A2(net819),
    .A3(net833),
    .A4(net795),
    .B1(net805),
    .X(net901));
 sky130_fd_sc_hd__a41o_1 c114 (.A1(net8),
    .A2(net2),
    .A3(net795),
    .A4(net995),
    .B1(net833),
    .X(net915));
 sky130_fd_sc_hd__mux4_1 c115 (.A0(net841),
    .A1(net817),
    .A2(net901),
    .A3(net844),
    .S0(net1014),
    .S1(net995),
    .X(net924));
 sky130_fd_sc_hd__a41o_1 c116 (.A1(net770),
    .A2(net7),
    .A3(net925),
    .A4(net924),
    .B1(net773),
    .X(net914));
 sky130_fd_sc_hd__mux4_1 c117 (.A0(net830),
    .A1(net846),
    .A2(net8),
    .A3(net996),
    .S0(net915),
    .S1(net804),
    .X(net9));
 sky130_fd_sc_hd__mux4_2 c118 (.A0(net819),
    .A1(net801),
    .A2(net924),
    .A3(net914),
    .S0(net1014),
    .S1(net8),
    .X(net10));
 sky130_fd_sc_hd__a41o_1 c119 (.A1(net1014),
    .A2(net10),
    .A3(net817),
    .A4(net1006),
    .B1(net804),
    .X(net11));
 sky130_fd_sc_hd__a41o_1 c120 (.A1(net770),
    .A2(net901),
    .A3(net995),
    .A4(net804),
    .B1(net819),
    .X(net927));
 sky130_fd_sc_hd__a41o_1 c121 (.A1(net833),
    .A2(net11),
    .A3(net787),
    .A4(net830),
    .B1(net847),
    .X(net926));
 sky130_fd_sc_hd__a41o_1 c122 (.A1(net809),
    .A2(net798),
    .A3(net927),
    .A4(net795),
    .B1(net1014),
    .X(net917));
 sky130_fd_sc_hd__a41o_1 c123 (.A1(net6),
    .A2(net10),
    .A3(net917),
    .A4(net11),
    .B1(net927),
    .X(net928));
 sky130_fd_sc_hd__mux4_2 c124 (.A0(net995),
    .A1(net770),
    .A2(net11),
    .A3(net804),
    .S0(net845),
    .S1(net1014),
    .X(net909));
 sky130_fd_sc_hd__mux4_2 c125 (.A0(net846),
    .A1(net848),
    .A2(net795),
    .A3(net828),
    .S0(net833),
    .S1(net770),
    .X(net899));
 sky130_fd_sc_hd__mux4_1 c126 (.A0(net9),
    .A1(net11),
    .A2(net803),
    .A3(net801),
    .S0(net825),
    .S1(net915),
    .X(net12));
 sky130_fd_sc_hd__mux4_1 c127 (.A0(net795),
    .A1(net917),
    .A2(net899),
    .A3(net833),
    .S0(net846),
    .S1(net928),
    .X(net871));
 sky130_fd_sc_hd__a41o_1 c128 (.A1(net12),
    .A2(net901),
    .A3(net917),
    .A4(net871),
    .B1(net839),
    .X(net929));
 sky130_fd_sc_hd__a41o_1 c129 (.A1(net828),
    .A2(net901),
    .A3(net899),
    .A4(net11),
    .B1(net805),
    .X(net13));
 sky130_fd_sc_hd__mux4_1 c130 (.A0(net13),
    .A1(net830),
    .A2(net929),
    .A3(net9),
    .S0(net10),
    .S1(net12),
    .X(net919));
 sky130_fd_sc_hd__mux4_1 c131 (.A0(net10),
    .A1(net899),
    .A2(net847),
    .A3(net890),
    .S0(net909),
    .S1(net919),
    .X(net14));
 sky130_fd_sc_hd__a41o_4 c132 (.A1(net998),
    .A2(net1024),
    .A3(net1007),
    .A4(net994),
    .B1(net1011),
    .X(net15));
 sky130_fd_sc_hd__a41o_4 c133 (.A1(net15),
    .A2(net1135),
    .A3(net1134),
    .A4(net993),
    .B1(net1021),
    .X(net16));
 sky130_fd_sc_hd__a31o_4 c134 (.A1(net1134),
    .A2(net756),
    .A3(net1135),
    .B1(net1010),
    .X(net922));
 sky130_fd_sc_hd__a41o_4 c135 (.A1(net991),
    .A2(net994),
    .A3(net756),
    .A4(net1024),
    .B1(net996),
    .X(net17));
 sky130_fd_sc_hd__a41o_4 c136 (.A1(net17),
    .A2(net980),
    .A3(net1006),
    .A4(net1010),
    .B1(net1016),
    .X(net18));
 sky130_fd_sc_hd__a31o_4 c137 (.A1(net999),
    .A2(net15),
    .A3(net1001),
    .B1(net1010),
    .X(net19));
 sky130_fd_sc_hd__a41o_4 c138 (.A1(net17),
    .A2(net1134),
    .A3(net1003),
    .A4(net993),
    .B1(net980),
    .X(net851));
 sky130_fd_sc_hd__a41o_4 c139 (.A1(net17),
    .A2(net994),
    .A3(net1005),
    .A4(net16),
    .B1(net979),
    .X(net20));
 sky130_fd_sc_hd__a41o_4 c140 (.A1(net1132),
    .A2(net1011),
    .A3(net977),
    .A4(net998),
    .B1(net18),
    .X(net21));
 sky130_fd_sc_hd__a41o_4 c141 (.A1(net979),
    .A2(net1003),
    .A3(net1132),
    .A4(net1010),
    .B1(net972),
    .X(net22));
 sky130_fd_sc_hd__mux4_2 c142 (.A0(net22),
    .A1(net753),
    .A2(net993),
    .A3(net977),
    .S0(net17),
    .S1(net972),
    .X(net23));
 sky130_fd_sc_hd__a41o_4 c143 (.A1(net971),
    .A2(net753),
    .A3(net18),
    .A4(net977),
    .B1(net972),
    .X(net24));
 sky130_fd_sc_hd__mux4_2 c144 (.A0(net971),
    .A1(net24),
    .A2(net1132),
    .A3(net977),
    .S0(net1010),
    .S1(net972),
    .X(net25));
 sky130_fd_sc_hd__mux4_2 c145 (.A0(net977),
    .A1(net1135),
    .A2(net25),
    .A3(net1132),
    .S0(net1133),
    .S1(net1134),
    .X(net26));
 sky130_fd_sc_hd__a41o_4 c146 (.A1(net26),
    .A2(net18),
    .A3(net993),
    .A4(net1121),
    .B1(net25),
    .X(net27));
 sky130_fd_sc_hd__mux4_2 c147 (.A0(net17),
    .A1(net1134),
    .A2(net24),
    .A3(net980),
    .S0(net1010),
    .S1(net972),
    .X(net28));
 sky130_fd_sc_hd__a41o_1 c148 (.A1(net970),
    .A2(net971),
    .A3(net25),
    .A4(net22),
    .B1(net972),
    .X(net857));
 sky130_fd_sc_hd__a41o_2 c149 (.A1(net1132),
    .A2(net22),
    .A3(net973),
    .A4(net967),
    .B1(net971),
    .X(net29));
 sky130_fd_sc_hd__mux4_2 c150 (.A0(net966),
    .A1(net753),
    .A2(net756),
    .A3(net980),
    .S0(net971),
    .S1(net967),
    .X(net30));
 sky130_fd_sc_hd__a41o_4 c151 (.A1(net1148),
    .A2(net970),
    .A3(net26),
    .A4(net965),
    .B1(net1121),
    .X(net866));
 sky130_fd_sc_hd__mux4_2 c152 (.A0(net994),
    .A1(net963),
    .A2(net962),
    .A3(net1121),
    .S0(net980),
    .S1(net965),
    .X(net31));
 sky130_fd_sc_hd__mux4_2 c153 (.A0(net958),
    .A1(net25),
    .A2(net962),
    .A3(net22),
    .S0(net18),
    .S1(net970),
    .X(net32));
 sky130_fd_sc_hd__a41o_2 c154 (.A1(net778),
    .A2(net1016),
    .A3(net1017),
    .A4(net996),
    .B1(net1117),
    .X(net33));
 sky130_fd_sc_hd__mux4_2 c155 (.A0(net1134),
    .A1(net33),
    .A2(net779),
    .A3(net1019),
    .S0(net1017),
    .S1(net778),
    .X(net34));
 sky130_fd_sc_hd__a41o_4 c156 (.A1(net967),
    .A2(net994),
    .A3(net34),
    .A4(net18),
    .B1(net979),
    .X(net35));
 sky130_fd_sc_hd__mux4_2 c157 (.A0(net980),
    .A1(net771),
    .A2(net772),
    .A3(net1019),
    .S0(net773),
    .S1(net1017),
    .X(net36));
 sky130_fd_sc_hd__a41o_1 c158 (.A1(net33),
    .A2(net22),
    .A3(net964),
    .A4(net967),
    .B1(net784),
    .X(net37));
 sky130_fd_sc_hd__a41o_2 c159 (.A1(net779),
    .A2(net1135),
    .A3(net960),
    .A4(net994),
    .B1(net36),
    .X(net38));
 sky130_fd_sc_hd__a41o_4 c160 (.A1(net960),
    .A2(net994),
    .A3(net36),
    .A4(net1024),
    .B1(net964),
    .X(net898));
 sky130_fd_sc_hd__a41o_2 c161 (.A1(net957),
    .A2(net38),
    .A3(net33),
    .A4(net960),
    .B1(net964),
    .X(net39));
 sky130_fd_sc_hd__a41o_2 c162 (.A1(net1001),
    .A2(net779),
    .A3(net999),
    .A4(net36),
    .B1(net33),
    .X(net911));
 sky130_fd_sc_hd__mux4_2 c163 (.A0(net756),
    .A1(net957),
    .A2(net1008),
    .A3(net772),
    .S0(net960),
    .S1(net964),
    .X(net40));
 sky130_fd_sc_hd__mux4_2 c164 (.A0(net953),
    .A1(net784),
    .A2(net1019),
    .A3(net965),
    .S0(net1021),
    .S1(net778),
    .X(net41));
 sky130_fd_sc_hd__mux4_2 c165 (.A0(net954),
    .A1(net911),
    .A2(net953),
    .A3(net753),
    .S0(net966),
    .S1(net1003),
    .X(net42));
 sky130_fd_sc_hd__a41o_4 c166 (.A1(net42),
    .A2(net756),
    .A3(net788),
    .A4(net992),
    .B1(net954),
    .X(net43));
 sky130_fd_sc_hd__a41o_4 c167 (.A1(net943),
    .A2(net771),
    .A3(net957),
    .A4(net960),
    .B1(net34),
    .X(net44));
 sky130_fd_sc_hd__mux4_2 c168 (.A0(net999),
    .A1(net18),
    .A2(net953),
    .A3(net948),
    .S0(net911),
    .S1(net44),
    .X(net45));
 sky130_fd_sc_hd__mux4_2 c169 (.A0(net960),
    .A1(net45),
    .A2(net911),
    .A3(net33),
    .S0(net772),
    .S1(net999),
    .X(net862));
 sky130_fd_sc_hd__mux4_2 c170 (.A0(net44),
    .A1(net1024),
    .A2(net779),
    .A3(net766),
    .S0(net786),
    .S1(net771),
    .X(net46));
 sky130_fd_sc_hd__mux4_2 c171 (.A0(net948),
    .A1(net780),
    .A2(net957),
    .A3(net46),
    .S0(net960),
    .S1(net953),
    .X(net47));
 sky130_fd_sc_hd__mux4_2 c172 (.A0(net38),
    .A1(net44),
    .A2(net34),
    .A3(net954),
    .S0(net45),
    .S1(net46),
    .X(net48));
 sky130_fd_sc_hd__mux4_2 c173 (.A0(net772),
    .A1(net1006),
    .A2(net48),
    .A3(net15),
    .S0(net957),
    .S1(net47),
    .X(net49));
 sky130_fd_sc_hd__mux4_2 c174 (.A0(net48),
    .A1(net47),
    .A2(net44),
    .A3(net38),
    .S0(net46),
    .S1(net1019),
    .X(net50));
 sky130_fd_sc_hd__mux4_2 c175 (.A0(net46),
    .A1(net1024),
    .A2(net935),
    .A3(net48),
    .S0(net958),
    .S1(net44),
    .X(net51));
 sky130_fd_sc_hd__mux4_2 c176 (.A0(net811),
    .A1(net806),
    .A2(net800),
    .A3(net18),
    .S0(net998),
    .S1(net1021),
    .X(net52));
 sky130_fd_sc_hd__mux4_2 c177 (.A0(net18),
    .A1(net780),
    .A2(net911),
    .A3(net1017),
    .S0(net962),
    .S1(net935),
    .X(net53));
 sky130_fd_sc_hd__mux4_2 c178 (.A0(net802),
    .A1(net794),
    .A2(net1008),
    .A3(net791),
    .S0(net809),
    .S1(net803),
    .X(net54));
 sky130_fd_sc_hd__mux4_2 c179 (.A0(net1006),
    .A1(net800),
    .A2(net963),
    .A3(net808),
    .S0(net52),
    .S1(net998),
    .X(net55));
 sky130_fd_sc_hd__a41o_1 c180 (.A1(net1019),
    .A2(net812),
    .A3(net790),
    .A4(net809),
    .B1(net1133),
    .X(net56));
 sky130_fd_sc_hd__a41o_4 c181 (.A1(net784),
    .A2(net56),
    .A3(net781),
    .A4(net53),
    .B1(net962),
    .X(net57));
 sky130_fd_sc_hd__a41o_2 c182 (.A1(net1016),
    .A2(net808),
    .A3(net813),
    .A4(net793),
    .B1(net998),
    .X(net58));
 sky130_fd_sc_hd__mux4_2 c183 (.A0(net1021),
    .A1(net811),
    .A2(net812),
    .A3(net800),
    .S0(net794),
    .S1(net802),
    .X(net869));
 sky130_fd_sc_hd__mux4_1 c184 (.A0(net771),
    .A1(net57),
    .A2(net1114),
    .A3(net55),
    .S0(net56),
    .S1(net36),
    .X(net59));
 sky130_fd_sc_hd__a41o_2 c185 (.A1(net56),
    .A2(net54),
    .A3(net53),
    .A4(net1008),
    .B1(net649),
    .X(net60));
 sky130_fd_sc_hd__mux4_2 c186 (.A0(net793),
    .A1(net1112),
    .A2(net55),
    .A3(net772),
    .S0(net52),
    .S1(net969),
    .X(net61));
 sky130_fd_sc_hd__mux4_2 c187 (.A0(net772),
    .A1(net55),
    .A2(net54),
    .A3(net798),
    .S0(net1025),
    .S1(net1112),
    .X(net62));
 sky130_fd_sc_hd__mux4_2 c188 (.A0(net44),
    .A1(net802),
    .A2(net62),
    .A3(net55),
    .S0(net784),
    .S1(net649),
    .X(net63));
 sky130_fd_sc_hd__mux4_1 c189 (.A0(net60),
    .A1(net792),
    .A2(net54),
    .A3(net998),
    .S0(net62),
    .S1(net650),
    .X(net64));
 sky130_fd_sc_hd__mux4_2 c190 (.A0(net58),
    .A1(net63),
    .A2(net54),
    .A3(net1133),
    .S0(net886),
    .S1(net649),
    .X(net65));
 sky130_fd_sc_hd__mux4_2 c191 (.A0(net65),
    .A1(net869),
    .A2(net1009),
    .A3(net802),
    .S0(net943),
    .S1(net1053),
    .X(net66));
 sky130_fd_sc_hd__mux4_2 c192 (.A0(net62),
    .A1(net63),
    .A2(net1113),
    .A3(net1032),
    .S0(net66),
    .S1(net802),
    .X(net67));
 sky130_fd_sc_hd__mux4_2 c193 (.A0(net63),
    .A1(net809),
    .A2(net66),
    .A3(net67),
    .S0(net808),
    .S1(net813),
    .X(net68));
 sky130_fd_sc_hd__mux4_1 c194 (.A0(net68),
    .A1(net793),
    .A2(net784),
    .A3(net1136),
    .S0(net67),
    .X(net69));
 sky130_fd_sc_hd__mux4_1 c195 (.A0(net67),
    .A1(net1113),
    .A2(net791),
    .A3(net58),
    .S0(net68),
    .S1(net886),
    .X(net70));
 sky130_fd_sc_hd__mux4_1 c196 (.A0(net68),
    .A1(net810),
    .A2(net53),
    .A3(net886),
    .S0(net650),
    .S1(net651),
    .X(net71));
 sky130_fd_sc_hd__a41o_1 c197 (.A1(net65),
    .A2(net63),
    .A3(net780),
    .A4(net1024),
    .B1(net886),
    .X(net72));
 sky130_fd_sc_hd__mux4_1 c198 (.A0(net1136),
    .A1(net816),
    .A2(net1009),
    .A3(net948),
    .S0(net60),
    .S1(net1015),
    .X(net73));
 sky130_fd_sc_hd__mux4_2 c199 (.A0(net1003),
    .A1(net817),
    .A2(net1085),
    .A3(net958),
    .S0(net935),
    .S1(net650),
    .X(net74));
 sky130_fd_sc_hd__mux4_2 c200 (.A0(net1081),
    .A1(net1114),
    .A2(net53),
    .A3(net1062),
    .S0(net836),
    .S1(net886),
    .X(net75));
 sky130_fd_sc_hd__mux4_2 c201 (.A0(net806),
    .A1(net819),
    .A2(net1053),
    .A3(net1081),
    .S0(net50),
    .S1(net986),
    .X(net76));
 sky130_fd_sc_hd__mux4_2 c202 (.A0(net1063),
    .A1(net799),
    .A2(net66),
    .A3(net1112),
    .S0(net806),
    .S1(net986),
    .X(net77));
 sky130_fd_sc_hd__mux4_2 c203 (.A0(net1022),
    .A1(net58),
    .A2(net824),
    .A3(net1021),
    .S0(net1006),
    .S1(net988),
    .X(net78));
 sky130_fd_sc_hd__mux4_2 c204 (.A0(net826),
    .A1(net814),
    .A2(net76),
    .A3(net767),
    .S0(net799),
    .S1(net987),
    .X(net79));
 sky130_fd_sc_hd__mux4_2 c205 (.A0(net823),
    .A1(net935),
    .A2(net78),
    .A3(net1008),
    .S0(net961),
    .S1(net987),
    .X(net80));
 sky130_fd_sc_hd__mux4_2 c206 (.A0(net816),
    .A1(net78),
    .A2(net80),
    .A3(net1009),
    .S0(net826),
    .S1(net986),
    .X(net81));
 sky130_fd_sc_hd__mux4_1 c207 (.A0(net79),
    .A1(net75),
    .A2(net66),
    .A3(net78),
    .S0(net76),
    .S1(net987),
    .X(net82));
 sky130_fd_sc_hd__mux4_2 c208 (.A0(net771),
    .A1(net80),
    .A2(net820),
    .A3(net1015),
    .S0(net986),
    .S1(net654),
    .X(net83));
 sky130_fd_sc_hd__mux4_1 c209 (.A0(net81),
    .A1(net55),
    .A2(net1133),
    .A3(net886),
    .S0(net986),
    .S1(net1128),
    .X(net84));
 sky130_fd_sc_hd__mux4_1 c210 (.A0(net76),
    .A1(net821),
    .A2(net72),
    .A3(net55),
    .S0(net81),
    .S1(net79),
    .X(net85));
 sky130_fd_sc_hd__mux4_1 c211 (.A0(net819),
    .A1(net1104),
    .A2(net60),
    .A3(net789),
    .S0(net886),
    .S1(net986),
    .X(net86));
 sky130_fd_sc_hd__mux4_1 c212 (.A0(net81),
    .A1(net792),
    .A2(net837),
    .A3(net1081),
    .S0(net582),
    .S1(net985),
    .X(net87));
 sky130_fd_sc_hd__mux4_1 c213 (.A0(net827),
    .A1(net34),
    .A2(net76),
    .A3(net77),
    .S0(net798),
    .S1(net1124),
    .X(net88));
 sky130_fd_sc_hd__mux4_1 c214 (.A0(net810),
    .A1(net773),
    .A2(net80),
    .A3(net75),
    .S0(net880),
    .S1(net985),
    .X(net89));
 sky130_fd_sc_hd__mux4_2 c215 (.A0(net836),
    .A1(net72),
    .A2(net54),
    .A3(net827),
    .S0(net559),
    .S1(net985),
    .X(net884));
 sky130_fd_sc_hd__mux4_2 c216 (.A0(net813),
    .A1(net72),
    .A2(net767),
    .A3(net583),
    .S0(net986),
    .S1(net654),
    .X(net90));
 sky130_fd_sc_hd__mux4_1 c217 (.A0(net83),
    .A1(net90),
    .A2(net1162),
    .A3(net767),
    .S0(net559),
    .S1(net985),
    .X(net91));
 sky130_fd_sc_hd__mux4_2 c218 (.A0(net54),
    .A1(net90),
    .A2(net583),
    .A3(net986),
    .S0(net654),
    .S1(net985),
    .X(net92));
 sky130_fd_sc_hd__mux4_1 c219 (.A0(net933),
    .A1(net819),
    .A2(net15),
    .A3(net90),
    .S0(net1105),
    .S1(net986),
    .X(net93));
 sky130_fd_sc_hd__mux4_1 c220 (.A0(net1014),
    .A1(net57),
    .A2(net825),
    .A3(net67),
    .S0(net582),
    .S1(net987),
    .X(net94));
 sky130_fd_sc_hd__mux4_2 c221 (.A0(net1054),
    .A1(net991),
    .A2(net3),
    .A3(net935),
    .S0(net814),
    .S1(net1025),
    .X(net95));
 sky130_fd_sc_hd__mux4_2 c222 (.A0(net815),
    .A1(net838),
    .A2(net1105),
    .A3(net905),
    .S0(net843),
    .S1(net582),
    .X(net918));
 sky130_fd_sc_hd__mux4_1 c223 (.A0(net81),
    .A1(net0),
    .A2(net1001),
    .A3(net843),
    .S0(net1024),
    .S1(net1104),
    .X(net96));
 sky130_fd_sc_hd__mux4_2 c224 (.A0(net956),
    .A1(net962),
    .A2(net817),
    .A3(net948),
    .S0(net1024),
    .S1(net589),
    .X(net97));
 sky130_fd_sc_hd__mux4_2 c225 (.A0(net767),
    .A1(net764),
    .A2(net97),
    .A3(net814),
    .S0(net925),
    .S1(net810),
    .X(net98));
 sky130_fd_sc_hd__mux4_2 c226 (.A0(net61),
    .A1(net890),
    .A2(net1136),
    .A3(net956),
    .S0(net776),
    .S1(net988),
    .X(net99));
 sky130_fd_sc_hd__mux4_1 c227 (.A0(net838),
    .A1(net978),
    .A2(net95),
    .A3(net1114),
    .S0(net1006),
    .S1(net805),
    .X(net100));
 sky130_fd_sc_hd__mux4_1 c228 (.A0(net834),
    .A1(net869),
    .A2(net95),
    .A3(net1020),
    .S0(net905),
    .S1(net969),
    .X(net908));
 sky130_fd_sc_hd__mux4_1 c229 (.A0(net95),
    .A1(net100),
    .A2(net1008),
    .A3(net834),
    .S0(net1115),
    .S1(net589),
    .X(net101));
 sky130_fd_sc_hd__mux4_1 c230 (.A0(net805),
    .A1(net1115),
    .A2(net933),
    .A3(net61),
    .S0(net589),
    .S1(clknet_1_0__leaf_net656),
    .X(net102));
 sky130_fd_sc_hd__mux4_1 c231 (.A0(net814),
    .A1(net100),
    .A2(net764),
    .A3(net79),
    .S0(net933),
    .S1(net659),
    .X(net103));
 sky130_fd_sc_hd__mux4_1 c232 (.A0(net98),
    .A1(net57),
    .A2(net52),
    .A3(net1014),
    .S0(clknet_1_0__leaf_net657),
    .S1(clknet_1_1__leaf_net658),
    .X(net104));
 sky130_fd_sc_hd__mux4_1 c233 (.A0(net1024),
    .A1(net925),
    .A2(net98),
    .A3(clknet_1_0__leaf_net657),
    .S0(clknet_1_0__leaf_net658),
    .S1(net870),
    .X(net105));
 sky130_fd_sc_hd__mux4_1 c234 (.A0(net100),
    .A1(clknet_1_0__leaf_net105),
    .A2(net0),
    .A3(net825),
    .S0(net1014),
    .S1(net987),
    .X(net106));
 sky130_fd_sc_hd__mux4_1 c235 (.A0(net822),
    .A1(clknet_1_1__leaf_net105),
    .A2(net577),
    .A3(net589),
    .S0(clknet_1_0__leaf_net658),
    .S1(net659),
    .X(net107));
 sky130_fd_sc_hd__mux4_1 c236 (.A0(net98),
    .A1(net53),
    .A2(net821),
    .A3(net903),
    .S0(net902),
    .S1(net987),
    .X(net108));
 sky130_fd_sc_hd__mux4_1 c237 (.A0(net90),
    .A1(net62),
    .A2(net956),
    .A3(net1020),
    .S0(clknet_1_0__leaf_net107),
    .S1(net870),
    .X(net109));
 sky130_fd_sc_hd__mux4_1 c238 (.A0(net822),
    .A1(net53),
    .A2(clknet_1_0__leaf_net105),
    .A3(net969),
    .S0(net583),
    .S1(net660),
    .X(net921));
 sky130_fd_sc_hd__mux4_1 c239 (.A0(clknet_1_0__leaf_net109),
    .A1(net79),
    .A2(clknet_1_0__leaf_net921),
    .A3(net850),
    .S0(net761),
    .S1(net651),
    .X(net110));
 sky130_fd_sc_hd__mux4_1 c240 (.A0(net108),
    .A1(clknet_1_0__leaf_net109),
    .A2(net98),
    .A3(net825),
    .S0(net1017),
    .S1(net589),
    .X(net111));
 sky130_fd_sc_hd__mux4_1 c241 (.A0(net5),
    .A1(net108),
    .A2(clknet_1_1__leaf_net921),
    .A3(net908),
    .S0(net910),
    .S1(net589),
    .X(net112));
 sky130_fd_sc_hd__mux4_1 c256 (.A0(net7),
    .A1(net100),
    .A2(net926),
    .A3(net998),
    .S0(net905),
    .S1(net776),
    .X(net113));
 sky130_fd_sc_hd__mux4_1 c257 (.A0(net825),
    .A1(net11),
    .A2(net7),
    .A3(clknet_1_0__leaf_net921),
    .S0(net901),
    .S1(net817),
    .X(net114));
 sky130_fd_sc_hd__mux4_1 c258 (.A0(net108),
    .A1(net905),
    .A2(net850),
    .A3(net919),
    .S0(net659),
    .S1(net662),
    .X(net115));
 sky130_fd_sc_hd__mux4_1 c259 (.A0(net11),
    .A1(net918),
    .A2(net909),
    .A3(clknet_1_1__leaf_net921),
    .S0(net1102),
    .S1(net661),
    .X(net116));
 sky130_fd_sc_hd__mux4_1 c260 (.A0(net776),
    .A1(net825),
    .A2(net845),
    .A3(net925),
    .S0(net589),
    .S1(net661),
    .X(net906));
 sky130_fd_sc_hd__mux4_1 c261 (.A0(net809),
    .A1(net926),
    .A2(net886),
    .A3(net920),
    .S0(net870),
    .S1(net662),
    .X(net900));
 sky130_fd_sc_hd__mux4_1 c262 (.A0(net52),
    .A1(net900),
    .A2(net844),
    .A3(net920),
    .S0(clknet_1_1__leaf_net658),
    .S1(net662),
    .X(net907));
 sky130_fd_sc_hd__mux4_1 c263 (.A0(net14),
    .A1(net850),
    .A2(net900),
    .A3(net52),
    .S0(net786),
    .S1(clknet_1_0__leaf_net907),
    .X(net931));
 sky130_fd_sc_hd__a41o_4 c264 (.A1(net994),
    .A2(net24),
    .A3(net979),
    .A4(net1148),
    .B1(net25),
    .X(net117));
 sky130_fd_sc_hd__a41o_2 c265 (.A1(net1005),
    .A2(net15),
    .A3(net991),
    .A4(net1015),
    .B1(net963),
    .X(net888));
 sky130_fd_sc_hd__a41o_1 c266 (.A1(net1016),
    .A2(net888),
    .A3(net1020),
    .A4(net971),
    .B1(net1121),
    .X(net118));
 sky130_fd_sc_hd__a41o_4 c267 (.A1(net1007),
    .A2(net26),
    .A3(net949),
    .A4(net1021),
    .B1(net117),
    .X(net119));
 sky130_fd_sc_hd__a41o_4 c268 (.A1(net993),
    .A2(net117),
    .A3(net1022),
    .A4(net949),
    .B1(net963),
    .X(net120));
 sky130_fd_sc_hd__a41o_1 c269 (.A1(net117),
    .A2(net1081),
    .A3(net888),
    .A4(net949),
    .B1(net993),
    .X(net121));
 sky130_fd_sc_hd__a41o_2 c270 (.A1(net120),
    .A2(net950),
    .A3(net26),
    .A4(net117),
    .B1(net999),
    .X(net122));
 sky130_fd_sc_hd__a41o_4 c271 (.A1(net955),
    .A2(net117),
    .A3(net980),
    .A4(net1052),
    .B1(net949),
    .X(net123));
 sky130_fd_sc_hd__a41o_4 c272 (.A1(net944),
    .A2(net121),
    .A3(net1003),
    .A4(net22),
    .B1(net949),
    .X(net124));
 sky130_fd_sc_hd__a41o_1 c273 (.A1(net124),
    .A2(net119),
    .A3(net951),
    .A4(net945),
    .B1(net967),
    .X(net125));
 sky130_fd_sc_hd__mux4_2 c274 (.A0(net1021),
    .A1(net122),
    .A2(net973),
    .A3(net1020),
    .S0(net944),
    .S1(net949),
    .X(net126));
 sky130_fd_sc_hd__a41o_2 c275 (.A1(net125),
    .A2(net756),
    .A3(net1119),
    .A4(net122),
    .B1(net949),
    .X(net127));
 sky130_fd_sc_hd__mux4_2 c276 (.A0(net1025),
    .A1(net124),
    .A2(net122),
    .A3(net1003),
    .S0(net944),
    .S1(net949),
    .X(net128));
 sky130_fd_sc_hd__a41o_1 c277 (.A1(net888),
    .A2(net121),
    .A3(net1119),
    .A4(net950),
    .B1(net942),
    .X(net129));
 sky130_fd_sc_hd__a41o_4 c278 (.A1(net128),
    .A2(net944),
    .A3(net994),
    .A4(net125),
    .B1(net949),
    .X(net130));
 sky130_fd_sc_hd__a41o_2 c279 (.A1(net1022),
    .A2(net127),
    .A3(net950),
    .A4(net15),
    .B1(net1119),
    .X(net131));
 sky130_fd_sc_hd__a41o_1 c280 (.A1(net753),
    .A2(net944),
    .A3(net942),
    .A4(net122),
    .B1(net949),
    .X(net132));
 sky130_fd_sc_hd__mux4_2 c281 (.A0(net121),
    .A1(net129),
    .A2(net130),
    .A3(net945),
    .S0(net937),
    .S1(net1117),
    .X(net133));
 sky130_fd_sc_hd__mux4_2 c282 (.A0(net936),
    .A1(net125),
    .A2(net937),
    .A3(net1100),
    .S0(net1119),
    .S1(net950),
    .X(net134));
 sky130_fd_sc_hd__mux4_2 c283 (.A0(net130),
    .A1(net121),
    .A2(net936),
    .A3(net124),
    .S0(net937),
    .S1(net1119),
    .X(net135));
 sky130_fd_sc_hd__mux4_2 c284 (.A0(net122),
    .A1(net128),
    .A2(net945),
    .A3(net937),
    .S0(net936),
    .S1(net942),
    .X(net136));
 sky130_fd_sc_hd__mux4_2 c285 (.A0(net134),
    .A1(net128),
    .A2(net937),
    .A3(net130),
    .S0(net135),
    .S1(net753),
    .X(net137));
 sky130_fd_sc_hd__mux4_2 c286 (.A0(net48),
    .A1(net1006),
    .A2(net948),
    .A3(net1007),
    .S0(net1085),
    .S1(net1135),
    .X(net138));
 sky130_fd_sc_hd__a41o_4 c287 (.A1(net789),
    .A2(net939),
    .A3(net131),
    .A4(net948),
    .B1(net1036),
    .X(net139));
 sky130_fd_sc_hd__a41o_4 c288 (.A1(net33),
    .A2(net945),
    .A3(net966),
    .A4(net943),
    .B1(net955),
    .X(net140));
 sky130_fd_sc_hd__a41o_1 c289 (.A1(net766),
    .A2(net140),
    .A3(net1089),
    .A4(net778),
    .B1(net936),
    .X(net141));
 sky130_fd_sc_hd__mux4_2 c290 (.A0(net1008),
    .A1(net1134),
    .A2(net1117),
    .A3(net776),
    .S0(net766),
    .S1(net955),
    .X(net142));
 sky130_fd_sc_hd__a41o_2 c291 (.A1(net773),
    .A2(net130),
    .A3(net51),
    .A4(net119),
    .B1(net1098),
    .X(net143));
 sky130_fd_sc_hd__mux4_1 c292 (.A0(net143),
    .A1(net1037),
    .A2(net787),
    .A3(net140),
    .S0(net1134),
    .S1(net117),
    .X(net144));
 sky130_fd_sc_hd__a41o_1 c293 (.A1(net24),
    .A2(net1134),
    .A3(net964),
    .A4(net1003),
    .B1(net1017),
    .X(net145));
 sky130_fd_sc_hd__mux4_2 c294 (.A0(net145),
    .A1(net142),
    .A2(net936),
    .A3(net946),
    .S0(net943),
    .S1(net117),
    .X(net146));
 sky130_fd_sc_hd__mux4_1 c295 (.A0(net129),
    .A1(net1008),
    .A2(net139),
    .A3(net143),
    .S0(net973),
    .X(net147));
 sky130_fd_sc_hd__sdfbbn_2 c296 (.CLK_N(clknet_4_2_0_clk),
    .D(net22),
    .RESET_B(net960),
    .SCD(net143),
    .SCE(net766),
    .SET_B(net1117),
    .Q(net149),
    .Q_N(net148));
 sky130_fd_sc_hd__mux4_2 c297 (.A0(net965),
    .A1(net145),
    .A2(net36),
    .A3(net766),
    .S0(net911),
    .S1(net953),
    .X(net150));
 sky130_fd_sc_hd__mux4_2 c298 (.A0(net150),
    .A1(net51),
    .A2(net778),
    .A3(net141),
    .S0(net148),
    .S1(net973),
    .X(net151));
 sky130_fd_sc_hd__mux4_1 c299 (.A0(net131),
    .A1(net129),
    .A2(net150),
    .A3(net148),
    .S0(net151),
    .S1(net581),
    .X(net152));
 sky130_fd_sc_hd__mux4_2 c300 (.A0(net141),
    .A1(net149),
    .A2(net150),
    .A3(net51),
    .S0(net1120),
    .S1(net146),
    .X(net153));
 sky130_fd_sc_hd__mux4_2 c301 (.A0(net34),
    .A1(net1112),
    .A2(net149),
    .A3(net1090),
    .S0(net1089),
    .S1(net967),
    .X(net154));
 sky130_fd_sc_hd__mux4_1 c302 (.A0(net151),
    .A1(net141),
    .A2(net148),
    .A3(net756),
    .S0(net939),
    .S1(net1120),
    .X(net155));
 sky130_fd_sc_hd__a41o_1 c303 (.A1(net36),
    .A2(net153),
    .A3(net1039),
    .A4(net148),
    .B1(net139),
    .X(net156));
 sky130_fd_sc_hd__mux4_2 c304 (.A0(net146),
    .A1(net50),
    .A2(net45),
    .A3(net1114),
    .S0(net138),
    .S1(net989),
    .X(net157));
 sky130_fd_sc_hd__mux4_2 c305 (.A0(net51),
    .A1(net149),
    .A2(net154),
    .A3(net1021),
    .S0(net581),
    .S1(net663),
    .X(net158));
 sky130_fd_sc_hd__mux4_1 c306 (.A0(net157),
    .A1(net942),
    .A2(net158),
    .A3(net51),
    .S0(net138),
    .S1(net989),
    .X(net159));
 sky130_fd_sc_hd__a41o_1 c307 (.A1(net121),
    .A2(net149),
    .A3(net131),
    .A4(net154),
    .B1(net608),
    .X(net160));
 sky130_fd_sc_hd__mux4_2 c308 (.A0(net808),
    .A1(net42),
    .A2(net911),
    .A3(net936),
    .S0(net1011),
    .S1(net581),
    .X(net161));
 sky130_fd_sc_hd__mux4_2 c309 (.A0(net141),
    .A1(net1135),
    .A2(net1009),
    .A3(net120),
    .S0(net1091),
    .S1(net581),
    .X(net162));
 sky130_fd_sc_hd__a41o_4 c310 (.A1(net797),
    .A2(net954),
    .A3(net1135),
    .A4(net946),
    .B1(net989),
    .X(net163));
 sky130_fd_sc_hd__a41o_1 c311 (.A1(net150),
    .A2(net808),
    .A3(net797),
    .A4(net161),
    .B1(net581),
    .X(net164));
 sky130_fd_sc_hd__mux4_2 c312 (.A0(net145),
    .A1(net790),
    .A2(net1006),
    .A3(net794),
    .S0(net1085),
    .S1(net797),
    .X(net165));
 sky130_fd_sc_hd__mux4_2 c313 (.A0(net1074),
    .A1(net165),
    .A2(net781),
    .A3(net42),
    .S0(net798),
    .S1(net581),
    .X(net885));
 sky130_fd_sc_hd__mux4_1 c314 (.A0(net119),
    .A1(net799),
    .A2(net951),
    .A3(net869),
    .S0(net1108),
    .S1(net161),
    .X(net166));
 sky130_fd_sc_hd__mux4_2 c315 (.A0(net166),
    .A1(net50),
    .A2(net979),
    .A3(net805),
    .S0(net165),
    .S1(net989),
    .X(net167));
 sky130_fd_sc_hd__mux4_2 c316 (.A0(net780),
    .A1(net163),
    .A2(net790),
    .A3(net161),
    .S0(net142),
    .S1(net1028),
    .X(net168));
 sky130_fd_sc_hd__a41o_1 c317 (.A1(net161),
    .A2(net885),
    .A3(net162),
    .A4(net954),
    .B1(net62),
    .X(net169));
 sky130_fd_sc_hd__mux4_1 c318 (.A0(net63),
    .A1(net1021),
    .A2(net162),
    .A3(net1093),
    .S0(net165),
    .S1(net891),
    .X(net170));
 sky130_fd_sc_hd__mux4_1 c319 (.A0(net781),
    .A1(net167),
    .A2(net1092),
    .A3(net1086),
    .S0(net780),
    .S1(net891),
    .X(net171));
 sky130_fd_sc_hd__mux4_2 c320 (.A0(net56),
    .A1(net164),
    .A2(net163),
    .A3(net122),
    .S0(net891),
    .S1(net983),
    .X(net172));
 sky130_fd_sc_hd__mux4_1 c321 (.A0(net167),
    .A1(net790),
    .A2(net165),
    .A3(net954),
    .S0(net172),
    .S1(net990),
    .X(net173));
 sky130_fd_sc_hd__mux4_2 c322 (.A0(net129),
    .A1(net161),
    .A2(net808),
    .A3(net581),
    .S0(net983),
    .S1(net665),
    .X(net174));
 sky130_fd_sc_hd__mux4_1 c323 (.A0(net862),
    .A1(net773),
    .A2(net161),
    .A3(net162),
    .S0(net989),
    .S1(net983),
    .X(net175));
 sky130_fd_sc_hd__mux4_1 c324 (.A0(net165),
    .A1(net174),
    .A2(net948),
    .A3(net172),
    .S0(net647),
    .S1(net1123),
    .X(net176));
 sky130_fd_sc_hd__mux4_2 c325 (.A0(net130),
    .A1(net163),
    .A2(net990),
    .A3(net891),
    .S0(net983),
    .S1(net665),
    .X(net879));
 sky130_fd_sc_hd__a41o_2 c326 (.A1(net879),
    .A2(net61),
    .A3(net888),
    .A4(net647),
    .B1(net665),
    .X(net177));
 sky130_fd_sc_hd__mux4_2 c327 (.A0(net163),
    .A1(net129),
    .A2(net177),
    .A3(net166),
    .S0(net1025),
    .S1(net990),
    .X(net896));
 sky130_fd_sc_hd__mux4_1 c328 (.A0(net177),
    .A1(net1006),
    .A2(net879),
    .A3(net948),
    .S0(net990),
    .S1(net983),
    .X(net178));
 sky130_fd_sc_hd__mux4_2 c329 (.A0(net178),
    .A1(net142),
    .A2(net885),
    .A3(net177),
    .S0(net990),
    .S1(net983),
    .X(net179));
 sky130_fd_sc_hd__mux4_1 c330 (.A0(net991),
    .A1(net799),
    .A2(net943),
    .A3(net1001),
    .S0(net773),
    .S1(net583),
    .X(net180));
 sky130_fd_sc_hd__mux4_1 c331 (.A0(net824),
    .A1(net15),
    .A2(net148),
    .A3(net969),
    .S0(net76),
    .S1(net647),
    .X(net181));
 sky130_fd_sc_hd__mux4_2 c332 (.A0(net149),
    .A1(net951),
    .A2(net65),
    .A3(net754),
    .S0(net776),
    .S1(net647),
    .X(net182));
 sky130_fd_sc_hd__mux4_1 c333 (.A0(net885),
    .A1(net174),
    .A2(net812),
    .A3(net180),
    .S0(net566),
    .S1(net650),
    .X(net183));
 sky130_fd_sc_hd__mux4_1 c334 (.A0(net180),
    .A1(net167),
    .A2(net1105),
    .A3(net140),
    .S0(net791),
    .S1(net985),
    .X(net184));
 sky130_fd_sc_hd__mux4_1 c335 (.A0(net80),
    .A1(net885),
    .A2(net764),
    .A3(net158),
    .S0(net884),
    .S1(net896),
    .X(net185));
 sky130_fd_sc_hd__mux4_1 c336 (.A0(net182),
    .A1(net948),
    .A2(net933),
    .A3(net986),
    .S0(net654),
    .S1(net983),
    .X(net186));
 sky130_fd_sc_hd__mux4_1 c337 (.A0(net72),
    .A1(net183),
    .A2(net933),
    .A3(net83),
    .S0(net831),
    .S1(net61),
    .X(net187));
 sky130_fd_sc_hd__mux4_2 c338 (.A0(net991),
    .A1(net879),
    .A2(net165),
    .A3(net989),
    .S0(net666),
    .S1(net667),
    .X(net188));
 sky130_fd_sc_hd__mux4_2 c339 (.A0(net820),
    .A1(net888),
    .A2(net803),
    .A3(net581),
    .S0(net666),
    .S1(net667),
    .X(net189));
 sky130_fd_sc_hd__mux4_2 c340 (.A0(net122),
    .A1(net182),
    .A2(net74),
    .A3(net966),
    .S0(net189),
    .S1(net831),
    .X(net190));
 sky130_fd_sc_hd__mux4_2 c341 (.A0(net55),
    .A1(net174),
    .A2(net1027),
    .A3(net61),
    .S0(net1017),
    .S1(net587),
    .X(net191));
 sky130_fd_sc_hd__mux4_2 c342 (.A0(net831),
    .A1(net821),
    .A2(net800),
    .A3(net182),
    .S0(net989),
    .S1(net985),
    .X(net873));
 sky130_fd_sc_hd__mux4_1 c343 (.A0(net158),
    .A1(net1005),
    .A2(net1086),
    .A3(net188),
    .S0(net990),
    .S1(net988),
    .X(net192));
 sky130_fd_sc_hd__mux4_2 c344 (.A0(net74),
    .A1(net188),
    .A2(net792),
    .A3(net960),
    .S0(net804),
    .S1(net668),
    .X(net193));
 sky130_fd_sc_hd__mux4_2 c345 (.A0(net180),
    .A1(net190),
    .A2(net995),
    .A3(net193),
    .S0(net581),
    .X(net635));
 sky130_fd_sc_hd__mux4_1 c346 (.A0(net965),
    .A1(net177),
    .A2(net191),
    .A3(net1115),
    .S0(net636),
    .S1(net666),
    .X(net195));
 sky130_fd_sc_hd__mux4_2 c347 (.A0(net990),
    .A1(net636),
    .A2(net988),
    .A3(net983),
    .S0(net666),
    .S1(net889),
    .X(net196));
 sky130_fd_sc_hd__mux4_2 c348 (.A0(net837),
    .A1(net196),
    .A2(net165),
    .A3(net873),
    .S0(net636),
    .S1(net669),
    .X(net197));
 sky130_fd_sc_hd__mux4_1 c349 (.A0(net168),
    .A1(net191),
    .A2(net1099),
    .A3(net55),
    .S0(net559),
    .S1(net666),
    .X(net198));
 sky130_fd_sc_hd__a41o_1 c350 (.A1(net1099),
    .A2(net884),
    .A3(net191),
    .B1(net636),
    .X(net199));
 sky130_fd_sc_hd__mux4_1 c351 (.A0(net183),
    .A1(net196),
    .A2(net197),
    .A3(net988),
    .S0(net668),
    .S1(net670),
    .X(net200));
 sky130_fd_sc_hd__mux4_1 c352 (.A0(net1075),
    .A1(net845),
    .A2(net960),
    .A3(net174),
    .S0(net1001),
    .S1(net789),
    .X(net201));
 sky130_fd_sc_hd__mux4_1 c353 (.A0(net947),
    .A1(net179),
    .A2(net143),
    .A3(net933),
    .S0(net62),
    .S1(net845),
    .X(net202));
 sky130_fd_sc_hd__mux4_1 c354 (.A0(net1104),
    .A1(net823),
    .A2(net873),
    .A3(net99),
    .S0(clknet_1_1__leaf_net644),
    .S1(net647),
    .X(net203));
 sky130_fd_sc_hd__mux4_1 c355 (.A0(net799),
    .A1(net3),
    .A2(net66),
    .A3(net98),
    .S0(net143),
    .S1(net823),
    .X(net204));
 sky130_fd_sc_hd__a41o_1 c356 (.A1(net4),
    .A2(net817),
    .A3(net849),
    .A4(net867),
    .B1(clknet_1_1__leaf_net644),
    .X(net887));
 sky130_fd_sc_hd__mux4_1 c357 (.A0(net0),
    .A1(net165),
    .A2(clknet_1_0__leaf_net107),
    .A3(net885),
    .S0(net812),
    .S1(net647),
    .X(net205));
 sky130_fd_sc_hd__mux4_1 c358 (.A0(net918),
    .A1(clknet_1_0__leaf_net205),
    .A2(net1009),
    .A3(net821),
    .S0(net880),
    .S1(clknet_1_0__leaf_net644),
    .X(net206));
 sky130_fd_sc_hd__mux4_1 c359 (.A0(net201),
    .A1(net1035),
    .A2(net905),
    .A3(net842),
    .S0(net933),
    .S1(net639),
    .X(net207));
 sky130_fd_sc_hd__mux4_1 c360 (.A0(clknet_1_0__leaf_net205),
    .A1(net182),
    .A2(net821),
    .A3(net3),
    .S0(net165),
    .S1(net895),
    .X(net208));
 sky130_fd_sc_hd__mux4_1 c361 (.A0(net812),
    .A1(net787),
    .A2(net77),
    .A3(net1087),
    .S0(net844),
    .S1(net817),
    .X(net209));
 sky130_fd_sc_hd__mux4_1 c362 (.A0(net849),
    .A1(clknet_1_1__leaf_net109),
    .A2(net97),
    .A3(net52),
    .S0(net845),
    .S1(net878),
    .X(net210));
 sky130_fd_sc_hd__mux4_1 c363 (.A0(net821),
    .A1(clknet_1_1__leaf_net205),
    .A2(net99),
    .A3(clknet_1_0__leaf_net912),
    .S0(clknet_1_0__leaf_net656),
    .S1(net889),
    .X(net211));
 sky130_fd_sc_hd__mux4_1 c364 (.A0(net95),
    .A1(net174),
    .A2(net947),
    .A3(net1061),
    .S0(net622),
    .S1(net895),
    .X(net212));
 sky130_fd_sc_hd__mux4_1 c365 (.A0(net1075),
    .A1(net799),
    .A2(net764),
    .A3(net916),
    .S0(clknet_1_0__leaf_net912),
    .S1(net639),
    .X(net213));
 sky130_fd_sc_hd__mux4_1 c366 (.A0(net165),
    .A1(net97),
    .A2(clknet_1_0__leaf_net203),
    .A3(net1025),
    .S0(net920),
    .S1(net666),
    .X(net214));
 sky130_fd_sc_hd__mux4_1 c367 (.A0(net212),
    .A1(net62),
    .A2(net77),
    .A3(net191),
    .S0(net916),
    .S1(net1125),
    .X(net215));
 sky130_fd_sc_hd__mux4_1 c368 (.A0(net3),
    .A1(net182),
    .A2(net95),
    .A3(net849),
    .S0(clknet_1_0__leaf_net644),
    .S1(net891),
    .X(net216));
 sky130_fd_sc_hd__mux4_1 c369 (.A0(net810),
    .A1(net97),
    .A2(net212),
    .A3(clknet_1_1__leaf_net216),
    .S0(net902),
    .S1(net982),
    .X(net217));
 sky130_fd_sc_hd__mux4_1 c370 (.A0(net213),
    .A1(net143),
    .A2(net212),
    .A3(clknet_1_0__leaf_net216),
    .S0(net78),
    .S1(net982),
    .X(net218));
 sky130_fd_sc_hd__mux4_1 c371 (.A0(net66),
    .A1(net76),
    .A2(clknet_1_0__leaf_net216),
    .A3(net68),
    .S0(net933),
    .S1(net982),
    .X(net219));
 sky130_fd_sc_hd__mux4_1 c372 (.A0(net57),
    .A1(net1104),
    .A2(clknet_1_0__leaf_net216),
    .A3(net622),
    .S0(clknet_1_1__leaf_net644),
    .S1(net666),
    .X(net220));
 sky130_fd_sc_hd__a41o_1 c373 (.A1(clknet_1_0__leaf_net216),
    .A2(clknet_1_1__leaf_net912),
    .A3(net622),
    .B1(net672),
    .X(net221));
 sky130_fd_sc_hd__a41o_2 c396 (.A1(net124),
    .A2(net1022),
    .A3(net973),
    .A4(net967),
    .B1(net993),
    .X(net222));
 sky130_fd_sc_hd__a41o_2 c397 (.A1(net963),
    .A2(net1003),
    .A3(net1007),
    .A4(net937),
    .B1(net974),
    .X(net223));
 sky130_fd_sc_hd__a41o_1 c398 (.A1(net941),
    .A2(net958),
    .A3(net130),
    .A4(net1066),
    .B1(net1134),
    .X(net224));
 sky130_fd_sc_hd__a41o_4 c399 (.A1(net980),
    .A2(net1095),
    .A3(net993),
    .A4(net937),
    .B1(net1071),
    .X(net225));
 sky130_fd_sc_hd__a41o_2 c400 (.A1(net941),
    .A2(net937),
    .A3(net934),
    .A4(net1051),
    .B1(net762),
    .X(net226));
 sky130_fd_sc_hd__a41o_2 c401 (.A1(net967),
    .A2(net1100),
    .A3(net1070),
    .A4(net934),
    .B1(net1005),
    .X(net227));
 sky130_fd_sc_hd__sdfbbn_1 c402 (.CLK_N(clknet_4_0_0_clk),
    .D(net227),
    .RESET_B(net888),
    .SCD(net224),
    .SCE(net1120),
    .SET_B(net1094),
    .Q(net229),
    .Q_N(net228));
 sky130_fd_sc_hd__mux4_2 c403 (.A0(net1070),
    .A1(net229),
    .A2(net753),
    .A3(net223),
    .S0(net224),
    .S1(net934),
    .X(net230));
 sky130_fd_sc_hd__a41o_2 c404 (.A1(net225),
    .A2(net127),
    .A3(net993),
    .A4(net119),
    .B1(net941),
    .X(net231));
 sky130_fd_sc_hd__sdfbbp_1 c405 (.CLK(clknet_4_0_0_clk),
    .D(net226),
    .RESET_B(net1022),
    .SCD(net223),
    .SCE(net1005),
    .SET_B(net993),
    .Q(net233),
    .Q_N(net232));
 sky130_fd_sc_hd__sdfbbn_2 c406 (.CLK_N(clknet_4_0_0_clk),
    .D(net227),
    .RESET_B(net1039),
    .SCD(net229),
    .SCE(net1105),
    .SET_B(net934),
    .Q(net235),
    .Q_N(net234));
 sky130_fd_sc_hd__sdfbbn_2 c407 (.CLK_N(clknet_4_0_0_clk),
    .D(net1100),
    .RESET_B(net233),
    .SCD(net231),
    .SCE(net226),
    .SET_B(net230),
    .Q(net237),
    .Q_N(net236));
 sky130_fd_sc_hd__sdfbbp_1 c408 (.CLK(clknet_4_4_0_clk),
    .D(net229),
    .RESET_B(net230),
    .SCD(net236),
    .SCE(net938),
    .SET_B(net1012),
    .Q(net239),
    .Q_N(net238));
 sky130_fd_sc_hd__sdfbbn_2 c409 (.CLK_N(clknet_4_4_0_clk),
    .D(net231),
    .RESET_B(net233),
    .SCD(net968),
    .SCE(net941),
    .SET_B(net234),
    .Q(net241),
    .Q_N(net240));
 sky130_fd_sc_hd__mux4_1 c410 (.A0(net224),
    .A1(net239),
    .A2(net1006),
    .A3(net945),
    .S0(net950),
    .S1(net226),
    .X(net242));
 sky130_fd_sc_hd__a41o_1 c411 (.A1(net237),
    .A2(net980),
    .A3(net238),
    .A4(net228),
    .B1(net231),
    .X(net243));
 sky130_fd_sc_hd__mux4_1 c412 (.A0(net756),
    .A1(net227),
    .A2(net232),
    .A3(net937),
    .S0(net228),
    .S1(clknet_1_0__leaf_net673),
    .X(net244));
 sky130_fd_sc_hd__mux4_1 c413 (.A0(net124),
    .A1(net223),
    .A2(net236),
    .A3(net230),
    .S0(net1135),
    .S1(clknet_1_0__leaf_net673),
    .X(net245));
 sky130_fd_sc_hd__mux4_1 c414 (.A0(net980),
    .A1(net238),
    .A2(net934),
    .A3(net575),
    .S0(clknet_1_0__leaf_net673),
    .S1(clknet_1_0__leaf_net674),
    .X(net246));
 sky130_fd_sc_hd__sdfbbn_2 c415 (.CLK_N(clknet_4_1_0_clk),
    .D(clknet_1_0__leaf_net246),
    .RESET_B(net233),
    .SCD(net575),
    .SCE(clknet_1_0__leaf_net673),
    .SET_B(clknet_1_0__leaf_net675),
    .Q(net248),
    .Q_N(net247));
 sky130_fd_sc_hd__mux4_1 c416 (.A0(net1155),
    .A1(net235),
    .A2(net232),
    .A3(net240),
    .S0(net247),
    .S1(clknet_1_0__leaf_net246),
    .X(net249));
 sky130_fd_sc_hd__mux4_1 c417 (.A0(net240),
    .A1(net941),
    .A2(net247),
    .A3(net576),
    .S0(clknet_1_1__leaf_net673),
    .S1(clknet_1_0__leaf_net675),
    .X(net250));
 sky130_fd_sc_hd__mux4_1 c418 (.A0(net753),
    .A1(net160),
    .A2(net41),
    .A3(net34),
    .S0(net942),
    .S1(net1025),
    .X(net251));
 sky130_fd_sc_hd__mux4_2 c419 (.A0(net762),
    .A1(net142),
    .A2(net1085),
    .A3(net34),
    .S0(net1068),
    .S1(net1120),
    .X(net252));
 sky130_fd_sc_hd__mux4_1 c420 (.A0(net776),
    .A1(net227),
    .A2(net252),
    .A3(net787),
    .S0(net942),
    .S1(net576),
    .X(net253));
 sky130_fd_sc_hd__mux4_2 c421 (.A0(net142),
    .A1(net1100),
    .A2(net150),
    .A3(net1019),
    .S0(net575),
    .S1(net679),
    .X(net254));
 sky130_fd_sc_hd__a41o_2 c422 (.A1(net51),
    .A2(net252),
    .A3(net234),
    .A4(net247),
    .B1(net787),
    .X(net255));
 sky130_fd_sc_hd__mux4_2 c423 (.A0(net1007),
    .A1(net937),
    .A2(net139),
    .A3(net789),
    .S0(net786),
    .S1(net679),
    .X(net256));
 sky130_fd_sc_hd__a41o_4 c424 (.A1(net252),
    .A2(net256),
    .A3(net778),
    .A4(net236),
    .B1(net678),
    .X(net257));
 sky130_fd_sc_hd__mux4_1 c425 (.A0(net117),
    .A1(net160),
    .A2(net932),
    .A3(net840),
    .S0(net256),
    .S1(net786),
    .X(net258));
 sky130_fd_sc_hd__mux4_1 c426 (.A0(net255),
    .A1(net227),
    .A2(net51),
    .A3(net252),
    .S0(net787),
    .S1(net576),
    .X(net259));
 sky130_fd_sc_hd__a41o_1 c427 (.A1(net256),
    .A2(net160),
    .A3(net1155),
    .A4(net840),
    .B1(net677),
    .X(net260));
 sky130_fd_sc_hd__a41o_1 c428 (.A1(net1009),
    .A2(net16),
    .A3(net252),
    .A4(net1039),
    .B1(net606),
    .X(net261));
 sky130_fd_sc_hd__mux4_1 c429 (.A0(net781),
    .A1(net38),
    .A2(net255),
    .A3(net225),
    .S0(net573),
    .S1(net608),
    .X(net262));
 sky130_fd_sc_hd__sdfbbp_1 c430 (.CLK(clknet_4_2_0_clk),
    .D(net1161),
    .RESET_B(net932),
    .SCD(net1017),
    .SCE(net576),
    .SET_B(net682),
    .Q(net264),
    .Q_N(net263));
 sky130_fd_sc_hd__mux4_1 c431 (.A0(net254),
    .A1(net35),
    .A2(net932),
    .A3(net263),
    .S0(net676),
    .S1(net678),
    .X(net265));
 sky130_fd_sc_hd__mux4_1 c432 (.A0(net1111),
    .A1(net254),
    .A2(net223),
    .A3(net261),
    .S0(clknet_1_0__leaf_net675),
    .S1(net681),
    .X(net266));
 sky130_fd_sc_hd__mux4_2 c433 (.A0(net263),
    .A1(net961),
    .A2(net1012),
    .A3(net573),
    .S0(net606),
    .S1(net683),
    .X(net267));
 sky130_fd_sc_hd__mux4_2 c434 (.A0(net840),
    .A1(net267),
    .A2(net254),
    .A3(net36),
    .S0(net680),
    .S1(net682),
    .X(net861));
 sky130_fd_sc_hd__a41o_2 c435 (.A1(net940),
    .A2(net951),
    .A3(net263),
    .A4(net247),
    .B1(net608),
    .X(net268));
 sky130_fd_sc_hd__mux4_1 c436 (.A0(net261),
    .A1(net940),
    .A2(net862),
    .A3(net932),
    .S0(net573),
    .S1(net680),
    .X(net269));
 sky130_fd_sc_hd__mux4_1 c437 (.A0(net268),
    .A1(net1133),
    .A2(net954),
    .A3(net940),
    .S0(net681),
    .S1(net684),
    .X(net270));
 sky130_fd_sc_hd__mux4_1 c438 (.A0(net254),
    .A1(net264),
    .A2(net268),
    .A3(net932),
    .S0(net940),
    .S1(net683),
    .X(net271));
 sky130_fd_sc_hd__mux4_1 c439 (.A0(net255),
    .A1(net268),
    .A2(net160),
    .A3(net573),
    .S0(net607),
    .S1(net684),
    .X(net272));
 sky130_fd_sc_hd__mux4_1 c440 (.A0(net1009),
    .A1(net162),
    .A2(net57),
    .A3(net268),
    .S0(net763),
    .S1(net153),
    .X(net273));
 sky130_fd_sc_hd__mux4_2 c441 (.A0(net130),
    .A1(net940),
    .A2(net966),
    .A3(net150),
    .S0(net886),
    .S1(net685),
    .X(net274));
 sky130_fd_sc_hd__mux4_2 c442 (.A0(net1065),
    .A1(net163),
    .A2(net789),
    .A3(net967),
    .S0(net840),
    .S1(net934),
    .X(net275));
 sky130_fd_sc_hd__mux4_1 c443 (.A0(net178),
    .A1(net241),
    .A2(net268),
    .A3(net274),
    .S0(net238),
    .S1(net983),
    .X(net276));
 sky130_fd_sc_hd__mux4_1 c444 (.A0(net1005),
    .A1(net794),
    .A2(net1086),
    .A3(net274),
    .S0(net275),
    .S1(net685),
    .X(net277));
 sky130_fd_sc_hd__mux4_2 c445 (.A0(net790),
    .A1(net798),
    .A2(net810),
    .A3(net177),
    .S0(net1085),
    .S1(net686),
    .X(net278));
 sky130_fd_sc_hd__mux4_1 c446 (.A0(net154),
    .A1(net275),
    .A2(net999),
    .A3(net1104),
    .S0(net607),
    .S1(net686),
    .X(net279));
 sky130_fd_sc_hd__mux4_1 c447 (.A0(net276),
    .A1(net162),
    .A2(net788),
    .A3(net254),
    .S0(net685),
    .S1(net686),
    .X(net280));
 sky130_fd_sc_hd__mux4_1 c448 (.A0(net162),
    .A1(net255),
    .A2(net1033),
    .A3(net172),
    .S0(net605),
    .S1(net683),
    .X(net281));
 sky130_fd_sc_hd__mux4_1 c449 (.A0(net1135),
    .A1(net951),
    .A2(net792),
    .A3(net942),
    .S0(net663),
    .S1(net893),
    .X(net282));
 sky130_fd_sc_hd__mux4_1 c450 (.A0(net61),
    .A1(net1050),
    .A2(net227),
    .A3(net282),
    .S0(net1008),
    .S1(net663),
    .X(net283));
 sky130_fd_sc_hd__mux4_2 c451 (.A0(net939),
    .A1(net786),
    .A2(net274),
    .A3(net23),
    .S0(net684),
    .S1(net688),
    .X(net284));
 sky130_fd_sc_hd__mux4_1 c452 (.A0(net278),
    .A1(net1033),
    .A2(net275),
    .A3(net57),
    .S0(net1113),
    .S1(net162),
    .X(net285));
 sky130_fd_sc_hd__mux4_1 c453 (.A0(net268),
    .A1(net172),
    .A2(net936),
    .A3(net637),
    .S0(net676),
    .S1(net690),
    .X(net286));
 sky130_fd_sc_hd__mux4_2 c454 (.A0(net139),
    .A1(net1055),
    .A2(net284),
    .A3(net235),
    .S0(net605),
    .S1(net690),
    .X(net897));
 sky130_fd_sc_hd__mux4_1 c455 (.A0(net164),
    .A1(net276),
    .A2(net241),
    .A3(net687),
    .S0(net690),
    .S1(net1127),
    .X(net287));
 sky130_fd_sc_hd__mux4_2 c456 (.A0(net282),
    .A1(net274),
    .A2(net284),
    .A3(net897),
    .S0(net637),
    .S1(net691),
    .X(net288));
 sky130_fd_sc_hd__mux4_1 c457 (.A0(net897),
    .A1(net288),
    .A2(net267),
    .A3(net605),
    .S0(net637),
    .S1(net1127),
    .X(net289));
 sky130_fd_sc_hd__mux4_1 c458 (.A0(net288),
    .A1(net792),
    .A2(net781),
    .A3(net961),
    .S0(net36),
    .S1(net981),
    .X(net290));
 sky130_fd_sc_hd__mux4_1 c459 (.A0(net275),
    .A1(net248),
    .A2(net68),
    .A3(net590),
    .S0(net607),
    .S1(net1129),
    .X(net291));
 sky130_fd_sc_hd__mux4_1 c460 (.A0(net167),
    .A1(net162),
    .A2(net261),
    .A3(net1069),
    .S0(net610),
    .S1(net637),
    .X(net292));
 sky130_fd_sc_hd__mux4_1 c461 (.A0(net162),
    .A1(net590),
    .A3(net984),
    .S0(net684),
    .S1(net692),
    .X(net293));
 sky130_fd_sc_hd__mux4_1 c462 (.A0(net792),
    .A1(net196),
    .A2(net237),
    .A3(net284),
    .S0(net1029),
    .S1(net961),
    .X(net294));
 sky130_fd_sc_hd__mux4_2 c463 (.A0(net823),
    .A1(net237),
    .A2(net958),
    .A3(net635),
    .S0(net668),
    .S1(net687),
    .X(net295));
 sky130_fd_sc_hd__mux4_1 c464 (.A0(net136),
    .A1(net294),
    .A2(net181),
    .A3(net654),
    .S0(net895),
    .S1(net893),
    .X(net296));
 sky130_fd_sc_hd__mux4_2 c465 (.A0(net168),
    .A1(net965),
    .A2(net997),
    .A3(net610),
    .S0(net667),
    .S1(net688),
    .X(net297));
 sky130_fd_sc_hd__mux4_1 c466 (.A0(net75),
    .A1(net248),
    .A2(net297),
    .A3(net1101),
    .S0(net663),
    .S1(net689),
    .X(net298));
 sky130_fd_sc_hd__mux4_1 c467 (.A0(net294),
    .A1(net1001),
    .A2(net248),
    .A3(net167),
    .S0(net933),
    .S1(net65),
    .X(net299));
 sky130_fd_sc_hd__mux4_1 c468 (.A0(net1076),
    .A1(net167),
    .A2(net247),
    .A3(net932),
    .S0(net754),
    .S1(clknet_1_0__leaf_net693),
    .X(net300));
 sky130_fd_sc_hd__mux4_1 c469 (.A0(net179),
    .A1(net227),
    .A2(net792),
    .A3(net663),
    .S0(clknet_1_1__leaf_net693),
    .S1(clknet_1_0__leaf_net694),
    .X(net301));
 sky130_fd_sc_hd__mux4_1 c470 (.A0(net177),
    .A1(net998),
    .A2(net568),
    .A3(clknet_1_0__leaf_net882),
    .S0(net669),
    .S1(clknet_1_1__leaf_net694),
    .X(net302));
 sky130_fd_sc_hd__mux4_1 c471 (.A0(net154),
    .A1(net824),
    .A2(net197),
    .A3(net765),
    .S0(net651),
    .S1(clknet_1_0__leaf_net693),
    .X(net303));
 sky130_fd_sc_hd__mux4_2 c472 (.A0(net15),
    .A1(net823),
    .A2(net884),
    .A3(net41),
    .S0(net225),
    .S1(net988),
    .X(net858));
 sky130_fd_sc_hd__mux4_2 c473 (.A0(net177),
    .A1(net941),
    .A2(net1001),
    .A3(net568),
    .S0(net616),
    .S1(net692),
    .X(net854));
 sky130_fd_sc_hd__mux4_1 c474 (.A0(net792),
    .A1(net53),
    .A2(net587),
    .A3(net679),
    .S0(clknet_1_1__leaf_net693),
    .S1(clknet_1_0__leaf_net694),
    .X(net868));
 sky130_fd_sc_hd__mux4_1 c475 (.A0(net196),
    .A1(net1046),
    .A2(net284),
    .A3(net52),
    .S0(net803),
    .S1(net568),
    .X(net304));
 sky130_fd_sc_hd__mux4_1 c476 (.A0(net1058),
    .A1(net136),
    .A2(net823),
    .A3(net1076),
    .S0(net1103),
    .S1(clknet_1_0__leaf_net693),
    .X(net305));
 sky130_fd_sc_hd__mux4_1 c477 (.A0(net58),
    .A1(clknet_1_0__leaf_net868),
    .A2(net1047),
    .A3(net304),
    .S0(clknet_1_0__leaf_net882),
    .S1(net637),
    .X(net306));
 sky130_fd_sc_hd__mux4_1 c478 (.A0(net896),
    .A1(net873),
    .A2(net858),
    .A3(clknet_1_0__leaf_net302),
    .S0(net568),
    .S1(net628),
    .X(net307));
 sky130_fd_sc_hd__mux4_1 c479 (.A0(clknet_1_0__leaf_net302),
    .A1(net77),
    .A2(net854),
    .A3(net83),
    .S0(net75),
    .S1(net883),
    .X(net308));
 sky130_fd_sc_hd__mux4_1 c480 (.A0(net197),
    .A1(net1048),
    .A2(net140),
    .A3(net297),
    .S0(net689),
    .S1(net697),
    .X(net309));
 sky130_fd_sc_hd__mux4_1 c481 (.A0(net1148),
    .A1(net120),
    .A2(net35),
    .A3(net904),
    .S0(clknet_1_0__leaf_net695),
    .S1(net696),
    .X(net310));
 sky130_fd_sc_hd__mux4_1 c482 (.A0(net941),
    .A1(clknet_1_0__leaf_net310),
    .A2(clknet_1_0__leaf_net868),
    .A3(clknet_1_0__leaf_net694),
    .S0(clknet_1_0__leaf_net695),
    .S1(net697),
    .X(net311));
 sky130_fd_sc_hd__mux4_1 c483 (.A0(net304),
    .A1(net858),
    .A2(clknet_1_0__leaf_net310),
    .A3(clknet_1_1__leaf_net302),
    .S0(net1001),
    .S1(net699),
    .X(net312));
 sky130_fd_sc_hd__mux4_2 c484 (.A0(net1015),
    .A1(net78),
    .A2(net845),
    .A3(net890),
    .S0(net566),
    .S1(net577),
    .X(net313));
 sky130_fd_sc_hd__mux4_1 c485 (.A0(net97),
    .A1(net842),
    .A2(clknet_1_1__leaf_net216),
    .A3(net823),
    .S0(clknet_1_1__leaf_net656),
    .S1(net678),
    .X(net314));
 sky130_fd_sc_hd__mux4_1 c486 (.A0(net98),
    .A1(net191),
    .A2(net754),
    .A3(net916),
    .S0(clknet_1_0__leaf_net657),
    .S1(net672),
    .X(net315));
 sky130_fd_sc_hd__mux4_1 c487 (.A0(net787),
    .A1(net803),
    .A2(net997),
    .A3(net76),
    .S0(clknet_1_1__leaf_net656),
    .S1(net982),
    .X(net316));
 sky130_fd_sc_hd__mux4_1 c488 (.A0(clknet_1_1__leaf_net105),
    .A1(net313),
    .A2(net897),
    .A3(net628),
    .S0(clknet_1_1__leaf_net657),
    .S1(net982),
    .X(net317));
 sky130_fd_sc_hd__mux4_1 c489 (.A0(clknet_1_1__leaf_net107),
    .A1(net76),
    .A2(net1007),
    .A3(net659),
    .S0(net672),
    .S1(net698),
    .X(net318));
 sky130_fd_sc_hd__mux4_1 c490 (.A0(net174),
    .A1(net98),
    .A2(net1001),
    .A3(clknet_1_0__leaf_net887),
    .S0(net146),
    .S1(net27),
    .X(net319));
 sky130_fd_sc_hd__mux4_1 c491 (.A0(net255),
    .A1(clknet_1_0__leaf_net310),
    .A2(clknet_1_0__leaf_net318),
    .A3(net934),
    .S0(net313),
    .S1(net699),
    .X(net320));
 sky130_fd_sc_hd__mux4_1 c492 (.A0(net843),
    .A1(net947),
    .A2(net235),
    .A3(clknet_1_1__leaf_net107),
    .S0(clknet_1_0__leaf_net319),
    .S1(net628),
    .X(net321));
 sky130_fd_sc_hd__mux4_1 c493 (.A0(clknet_1_1__leaf_net216),
    .A1(net862),
    .A2(net99),
    .A3(net783),
    .S0(net146),
    .S1(net607),
    .X(net322));
 sky130_fd_sc_hd__mux4_1 c494 (.A0(net933),
    .A1(clknet_1_0__leaf_net319),
    .A2(net154),
    .A3(net862),
    .S0(net616),
    .S1(clknet_1_1__leaf_net657),
    .X(net323));
 sky130_fd_sc_hd__mux4_1 c495 (.A0(net317),
    .A1(net956),
    .A2(net842),
    .A3(clknet_1_1__leaf_net107),
    .S0(net920),
    .S1(net690),
    .X(net324));
 sky130_fd_sc_hd__mux4_1 c496 (.A0(net154),
    .A1(net252),
    .A2(clknet_1_0__leaf_net887),
    .A3(net902),
    .S0(net982),
    .S1(net700),
    .X(net325));
 sky130_fd_sc_hd__mux4_1 c497 (.A0(clknet_1_1__leaf_net318),
    .A1(net67),
    .A2(net92),
    .A3(net862),
    .S0(net284),
    .S1(net982),
    .X(net326));
 sky130_fd_sc_hd__mux4_1 c498 (.A0(clknet_1_0__leaf_net203),
    .A1(clknet_1_0__leaf_net868),
    .A2(net832),
    .A3(net920),
    .S0(net679),
    .S1(clknet_1_1__leaf_net695),
    .X(net327));
 sky130_fd_sc_hd__mux4_1 c499 (.A0(net325),
    .A1(net903),
    .A2(net50),
    .A3(net1108),
    .S0(net805),
    .S1(net702),
    .X(net328));
 sky130_fd_sc_hd__mux4_1 c500 (.A0(net139),
    .A1(net823),
    .A2(clknet_1_1__leaf_net216),
    .A3(net1161),
    .S0(clknet_1_1__leaf_net882),
    .S1(net702),
    .X(net329));
 sky130_fd_sc_hd__mux4_2 c501 (.A0(net823),
    .A1(net146),
    .A2(net842),
    .A3(net902),
    .S0(net988),
    .S1(net702),
    .X(net892));
 sky130_fd_sc_hd__mux4_1 c502 (.A0(net78),
    .A1(net819),
    .A2(net892),
    .A3(net99),
    .S0(net999),
    .S1(net765),
    .X(net330));
 sky130_fd_sc_hd__mux4_2 c503 (.A0(net27),
    .A1(net892),
    .A2(net843),
    .A3(net660),
    .S0(net692),
    .S1(net701),
    .X(net331));
 sky130_fd_sc_hd__mux4_1 c504 (.A0(net191),
    .A1(net237),
    .A2(net120),
    .A3(net892),
    .S0(net672),
    .S1(net701),
    .X(net332));
 sky130_fd_sc_hd__mux4_1 c505 (.A0(net52),
    .A1(net330),
    .A2(net892),
    .A3(net606),
    .S0(net902),
    .S1(net1122),
    .X(net333));
 sky130_fd_sc_hd__sdfbbn_2 c528 (.CLK_N(clknet_4_4_0_clk),
    .D(net1086),
    .RESET_B(net230),
    .SCD(net965),
    .SCE(net1012),
    .SET_B(clknet_1_0__leaf_net674),
    .Q(net335),
    .Q_N(net334));
 sky130_fd_sc_hd__a41o_1 c529 (.A1(net125),
    .A2(net223),
    .A3(net962),
    .A4(net1161),
    .B1(net951),
    .X(net336));
 sky130_fd_sc_hd__a41o_1 c530 (.A1(net131),
    .A2(net952),
    .A3(net999),
    .A4(net226),
    .B1(net938),
    .X(net337));
 sky130_fd_sc_hd__mux4_1 c531 (.A0(net231),
    .A1(net241),
    .A2(net996),
    .A3(net234),
    .S0(net1012),
    .S1(clknet_1_0__leaf_net675),
    .X(net338));
 sky130_fd_sc_hd__sdfbbn_1 c532 (.CLK_N(clknet_4_1_0_clk),
    .D(net119),
    .RESET_B(net1052),
    .SCD(net955),
    .SCE(net226),
    .SET_B(net979),
    .Q(net340),
    .Q_N(net339));
 sky130_fd_sc_hd__a41o_2 c533 (.A1(net1133),
    .A2(net336),
    .A3(net1095),
    .A4(net938),
    .B1(net974),
    .X(net874));
 sky130_fd_sc_hd__a41o_1 c534 (.A1(net968),
    .A2(net336),
    .A3(net339),
    .A4(net228),
    .B1(clknet_1_0__leaf_net673),
    .X(net341));
 sky130_fd_sc_hd__a41o_1 c535 (.A1(net232),
    .A2(net1003),
    .A3(net1012),
    .A4(net561),
    .B1(clknet_1_1__leaf_net674),
    .X(net342));
 sky130_fd_sc_hd__mux4_1 c536 (.A0(net224),
    .A1(net874),
    .A2(clknet_1_0__leaf_net342),
    .A3(net339),
    .S0(net1098),
    .S1(net1012),
    .X(net343));
 sky130_fd_sc_hd__mux4_1 c537 (.A0(net759),
    .A1(clknet_1_0__leaf_net342),
    .A2(clknet_1_0__leaf_net343),
    .A3(net1098),
    .S0(net1012),
    .S1(clknet_1_0__leaf_net675),
    .X(net344));
 sky130_fd_sc_hd__sdfbbp_1 c538 (.CLK(clknet_4_4_0_clk),
    .D(net336),
    .RESET_B(clknet_1_0__leaf_net342),
    .SCD(clknet_1_1__leaf_net246),
    .SCE(net999),
    .SET_B(net334),
    .Q(net346),
    .Q_N(net345));
 sky130_fd_sc_hd__a41o_1 c539 (.A1(clknet_1_0__leaf_net342),
    .A2(net952),
    .A3(net965),
    .A4(net1007),
    .B1(net345),
    .X(net347));
 sky130_fd_sc_hd__mux4_1 c540 (.A0(net335),
    .A1(net340),
    .A2(net1004),
    .A3(net1005),
    .S0(net974),
    .S1(clknet_1_1__leaf_net674),
    .X(net348));
 sky130_fd_sc_hd__mux4_1 c541 (.A0(net1052),
    .A1(net125),
    .A2(clknet_1_0__leaf_net250),
    .A3(net1022),
    .S0(clknet_1_0__leaf_net341),
    .S1(net705),
    .X(net349));
 sky130_fd_sc_hd__sdfbbn_1 c542 (.CLK_N(clknet_4_4_0_clk),
    .D(net1020),
    .RESET_B(clknet_1_0__leaf_net348),
    .SCD(clknet_1_0__leaf_net246),
    .SCE(net962),
    .SET_B(net231),
    .Q(net351),
    .Q_N(net350));
 sky130_fd_sc_hd__mux4_1 c543 (.A0(net346),
    .A1(net335),
    .A2(net970),
    .A3(net1118),
    .S0(net350),
    .S1(clknet_1_1__leaf_net674),
    .X(net352));
 sky130_fd_sc_hd__a41o_1 c544 (.A1(net136),
    .A2(clknet_1_0__leaf_net341),
    .A3(clknet_1_0__leaf_net348),
    .A4(clknet_1_1__leaf_net347),
    .B1(clknet_1_0__leaf_net352),
    .X(net353));
 sky130_fd_sc_hd__mux4_1 c545 (.A0(net226),
    .A1(net999),
    .A2(net339),
    .A3(net231),
    .S0(clknet_1_0__leaf_net352),
    .S1(clknet_1_1__leaf_net353),
    .X(net354));
 sky130_fd_sc_hd__sdfbbn_1 c546 (.CLK_N(clknet_4_4_0_clk),
    .D(net127),
    .RESET_B(net351),
    .SCD(clknet_1_0__leaf_net353),
    .SCE(clknet_1_0__leaf_net352),
    .SET_B(clknet_1_0__leaf_net349),
    .Q(net356),
    .Q_N(net355));
 sky130_fd_sc_hd__a41o_1 c547 (.A1(net1155),
    .A2(net1133),
    .A3(clknet_1_0__leaf_net347),
    .A4(net355),
    .B1(clknet_1_0__leaf_net352),
    .X(net357));
 sky130_fd_sc_hd__mux4_1 c548 (.A0(net229),
    .A1(net356),
    .A2(clknet_1_0__leaf_net347),
    .A3(clknet_1_0__leaf_net352),
    .S0(net1016),
    .S1(net706),
    .X(net358));
 sky130_fd_sc_hd__mux4_1 c549 (.A0(net230),
    .A1(clknet_1_0__leaf_net353),
    .A2(net355),
    .A3(net340),
    .S0(net946),
    .S1(net562),
    .X(net359));
 sky130_fd_sc_hd__mux4_1 c550 (.A0(net160),
    .A1(clknet_1_0__leaf_net341),
    .A2(net1020),
    .A3(net240),
    .S0(net932),
    .S1(net1019),
    .X(net360));
 sky130_fd_sc_hd__mux4_1 c551 (.A0(net138),
    .A1(net223),
    .A2(net932),
    .A3(net934),
    .S0(clknet_1_0__leaf_net352),
    .S1(net855),
    .X(net361));
 sky130_fd_sc_hd__mux4_1 c552 (.A0(net139),
    .A1(net160),
    .A2(net979),
    .A3(net225),
    .S0(clknet_1_0__leaf_net352),
    .S1(net955),
    .X(net362));
 sky130_fd_sc_hd__mux4_1 c553 (.A0(net1039),
    .A1(net36),
    .A2(net131),
    .A3(net1012),
    .S0(net605),
    .S1(net706),
    .X(net363));
 sky130_fd_sc_hd__mux4_1 c554 (.A0(net38),
    .A1(net150),
    .A2(net225),
    .A3(net248),
    .S0(net254),
    .S1(net709),
    .X(net364));
 sky130_fd_sc_hd__mux4_1 c555 (.A0(net351),
    .A1(net140),
    .A2(net932),
    .A3(net241),
    .S0(net237),
    .S1(net709),
    .X(net365));
 sky130_fd_sc_hd__mux4_1 c556 (.A0(net157),
    .A1(net1072),
    .A2(net270),
    .A3(clknet_1_0__leaf_net348),
    .S0(net350),
    .S1(net139),
    .X(net366));
 sky130_fd_sc_hd__mux4_1 c557 (.A0(net778),
    .A1(net38),
    .A2(net120),
    .A3(net786),
    .S0(clknet_1_0__leaf_net341),
    .S1(net709),
    .X(net367));
 sky130_fd_sc_hd__mux4_1 c558 (.A0(clknet_1_1__leaf_net367),
    .A1(net1041),
    .A2(net778),
    .A3(net119),
    .S0(net1022),
    .S1(clknet_1_0__leaf_net366),
    .X(net368));
 sky130_fd_sc_hd__mux4_1 c559 (.A0(clknet_1_0__leaf_net367),
    .A1(clknet_1_0__leaf_net341),
    .A2(net862),
    .A3(clknet_1_0__leaf_net343),
    .S0(net138),
    .S1(net364),
    .X(net369));
 sky130_fd_sc_hd__mux4_1 c560 (.A0(clknet_1_1__leaf_net347),
    .A1(clknet_1_0__leaf_net348),
    .A2(net1005),
    .A3(net605),
    .S0(net709),
    .S1(net712),
    .X(net370));
 sky130_fd_sc_hd__mux4_1 c561 (.A0(net954),
    .A1(net150),
    .A2(net1022),
    .A3(net240),
    .S0(clknet_1_0__leaf_net349),
    .S1(net712),
    .X(net371));
 sky130_fd_sc_hd__mux4_1 c562 (.A0(net334),
    .A1(net363),
    .A2(net157),
    .A3(clknet_1_0__leaf_net370),
    .S0(net561),
    .S1(clknet_1_1__leaf_net713),
    .X(net372));
 sky130_fd_sc_hd__mux4_1 c563 (.A0(clknet_1_1__leaf_net353),
    .A1(net1068),
    .A2(net585),
    .A3(net855),
    .S0(net712),
    .S1(clknet_1_0__leaf_net713),
    .X(net373));
 sky130_fd_sc_hd__mux4_1 c564 (.A0(clknet_1_0__leaf_net366),
    .A1(net157),
    .A2(clknet_1_1__leaf_net367),
    .A3(net707),
    .S0(clknet_1_0__leaf_net713),
    .S1(clknet_1_0__leaf_net714),
    .X(net374));
 sky130_fd_sc_hd__mux4_1 c565 (.A0(net970),
    .A1(net706),
    .A2(net855),
    .A3(clknet_1_1__leaf_net713),
    .S0(clknet_1_0__leaf_net714),
    .S1(clknet_1_0__leaf_net715),
    .X(net375));
 sky130_fd_sc_hd__mux4_1 c566 (.A0(clknet_1_0__leaf_net357),
    .A1(net940),
    .A2(net936),
    .A3(clknet_1_1__leaf_net372),
    .S0(clknet_1_0__leaf_net714),
    .S1(clknet_1_1__leaf_net715),
    .X(net376));
 sky130_fd_sc_hd__mux4_1 c567 (.A0(clknet_1_0__leaf_net375),
    .A1(net1080),
    .A2(net940),
    .A3(net683),
    .S0(net712),
    .S1(clknet_1_1__leaf_net715),
    .X(net377));
 sky130_fd_sc_hd__mux4_1 c568 (.A0(net223),
    .A1(net264),
    .A2(clknet_1_1__leaf_net349),
    .A3(net855),
    .S0(net712),
    .S1(net716),
    .X(net378));
 sky130_fd_sc_hd__mux4_1 c569 (.A0(net119),
    .A1(clknet_1_1__leaf_net349),
    .A2(clknet_1_1__leaf_net366),
    .A3(net151),
    .S0(net585),
    .S1(net718),
    .X(net379));
 sky130_fd_sc_hd__mux4_1 c570 (.A0(clknet_1_1__leaf_net375),
    .A1(clknet_1_0__leaf_net377),
    .A2(net712),
    .A3(clknet_1_0__leaf_net715),
    .S0(net719),
    .S1(net721),
    .X(net380));
 sky130_fd_sc_hd__mux4_1 c571 (.A0(clknet_1_0__leaf_net380),
    .A1(net940),
    .A2(clknet_1_0__leaf_net349),
    .A3(clknet_1_0__leaf_net366),
    .S0(net706),
    .S1(net720),
    .X(net381));
 sky130_fd_sc_hd__mux4_1 c572 (.A0(clknet_1_0__leaf_net372),
    .A1(net874),
    .A2(net150),
    .A3(net1086),
    .S0(net794),
    .S1(net663),
    .X(net382));
 sky130_fd_sc_hd__mux4_1 c573 (.A0(net172),
    .A1(net1069),
    .A2(net150),
    .A3(net939),
    .S0(net810),
    .S1(net996),
    .X(net383));
 sky130_fd_sc_hd__mux4_1 c574 (.A0(clknet_1_0__leaf_net367),
    .A1(clknet_1_1__leaf_net348),
    .A2(net1001),
    .A3(net651),
    .S0(net686),
    .S1(net705),
    .X(net384));
 sky130_fd_sc_hd__mux4_2 c575 (.A0(net794),
    .A1(net961),
    .A2(net278),
    .A3(net604),
    .S0(net981),
    .S1(net718),
    .X(net385));
 sky130_fd_sc_hd__mux4_1 c576 (.A0(net1013),
    .A1(net789),
    .A2(net604),
    .A3(net648),
    .S0(net984),
    .S1(net690),
    .X(net386));
 sky130_fd_sc_hd__mux4_1 c577 (.A0(net363),
    .A1(net288),
    .A2(net805),
    .A3(net648),
    .S0(net705),
    .S1(net708),
    .X(net387));
 sky130_fd_sc_hd__mux4_2 c578 (.A0(net1068),
    .A1(net954),
    .A2(net1040),
    .A3(net810),
    .S0(net942),
    .S1(net719),
    .X(net388));
 sky130_fd_sc_hd__mux4_2 c579 (.A0(net264),
    .A1(net1007),
    .A2(net1098),
    .A3(net386),
    .S0(net236),
    .S1(net705),
    .X(net389));
 sky130_fd_sc_hd__mux4_1 c580 (.A0(net267),
    .A1(net998),
    .A2(clknet_1_0__leaf_net377),
    .A3(net172),
    .S0(net706),
    .S1(net712),
    .X(net390));
 sky130_fd_sc_hd__mux4_1 c581 (.A0(net241),
    .A1(net942),
    .A2(net996),
    .A3(net637),
    .S0(net648),
    .S1(net720),
    .X(net391));
 sky130_fd_sc_hd__mux4_1 c582 (.A0(net391),
    .A1(net388),
    .A2(net21),
    .A3(net172),
    .S0(clknet_1_1__leaf_net348),
    .S1(net648),
    .X(net392));
 sky130_fd_sc_hd__mux4_1 c583 (.A0(clknet_1_1__leaf_net343),
    .A1(net278),
    .A2(net385),
    .A3(net1007),
    .S0(net62),
    .S1(net723),
    .X(net393));
 sky130_fd_sc_hd__mux4_1 c584 (.A0(clknet_1_1__leaf_net348),
    .A1(net21),
    .A2(net241),
    .A3(net288),
    .S0(net648),
    .S1(net716),
    .X(net394));
 sky130_fd_sc_hd__mux4_1 c585 (.A0(net364),
    .A1(net783),
    .A2(net810),
    .A3(net163),
    .S0(net869),
    .S1(net1002),
    .X(net395));
 sky130_fd_sc_hd__mux4_2 c586 (.A0(net236),
    .A1(net225),
    .A2(net706),
    .A3(net722),
    .S0(net723),
    .S1(net724),
    .X(net872));
 sky130_fd_sc_hd__mux4_2 c587 (.A0(net388),
    .A1(net955),
    .A2(net267),
    .A3(net254),
    .S0(net140),
    .S1(net627),
    .X(net396));
 sky130_fd_sc_hd__mux4_1 c588 (.A0(clknet_1_1__leaf_net349),
    .A1(clknet_1_1__leaf_net342),
    .A2(net248),
    .A3(net1108),
    .S0(net710),
    .S1(net724),
    .X(net397));
 sky130_fd_sc_hd__mux4_1 c589 (.A0(clknet_1_1__leaf_net380),
    .A1(net36),
    .A2(net284),
    .A3(net872),
    .S0(net865),
    .S1(net648),
    .X(net398));
 sky130_fd_sc_hd__mux4_1 c590 (.A0(net1073),
    .A1(net389),
    .A2(clknet_1_1__leaf_net348),
    .A3(net872),
    .S0(net968),
    .S1(net723),
    .X(net399));
 sky130_fd_sc_hd__mux4_1 c591 (.A0(clknet_1_1__leaf_net377),
    .A1(clknet_1_1__leaf_net367),
    .A2(net385),
    .A3(net590),
    .S0(net692),
    .S1(net723),
    .X(net400));
 sky130_fd_sc_hd__mux4_2 c592 (.A0(net386),
    .A1(net278),
    .A2(net240),
    .A3(net391),
    .S0(net590),
    .S1(net729),
    .X(net401));
 sky130_fd_sc_hd__mux4_1 c593 (.A0(net396),
    .A1(net872),
    .A2(net401),
    .A3(net783),
    .S0(net725),
    .S1(net729),
    .X(net402));
 sky130_fd_sc_hd__mux4_1 c594 (.A0(clknet_1_1__leaf_net370),
    .A1(net874),
    .A2(net389),
    .A3(net1042),
    .S0(net962),
    .S1(net650),
    .X(net403));
 sky130_fd_sc_hd__mux4_1 c595 (.A0(net248),
    .A1(net53),
    .A2(net832),
    .A3(net962),
    .S0(clknet_1_0__leaf_net868),
    .S1(net627),
    .X(net404));
 sky130_fd_sc_hd__mux4_1 c596 (.A0(net274),
    .A1(net268),
    .A2(net1098),
    .A3(net297),
    .S0(net652),
    .S1(clknet_1_1__leaf_net694),
    .X(net405));
 sky130_fd_sc_hd__mux4_2 c597 (.A0(net177),
    .A1(net948),
    .A2(net873),
    .A3(net800),
    .S0(net904),
    .S1(net722),
    .X(net406));
 sky130_fd_sc_hd__mux4_1 c598 (.A0(clknet_1_1__leaf_net342),
    .A1(net873),
    .A2(net1017),
    .A3(net805),
    .S0(net632),
    .S1(clknet_1_1__leaf_net714),
    .X(net407));
 sky130_fd_sc_hd__mux4_1 c599 (.A0(clknet_1_1__leaf_net407),
    .A1(net763),
    .A2(net941),
    .A3(net235),
    .S0(clknet_1_1__leaf_net694),
    .S1(net711),
    .X(net408));
 sky130_fd_sc_hd__mux4_1 c600 (.A0(net35),
    .A1(net873),
    .A2(net832),
    .A3(net406),
    .S0(net257),
    .S1(clknet_1_1__leaf_net695),
    .X(net409));
 sky130_fd_sc_hd__mux4_1 c601 (.A0(net969),
    .A1(net1002),
    .A2(net140),
    .A3(net824),
    .S0(net627),
    .S1(net628),
    .X(net410));
 sky130_fd_sc_hd__mux4_1 c602 (.A0(net941),
    .A1(net401),
    .A2(net873),
    .A3(clknet_1_1__leaf_net352),
    .S0(net824),
    .S1(net638),
    .X(net411));
 sky130_fd_sc_hd__mux4_1 c603 (.A0(net75),
    .A1(clknet_1_0__leaf_net407),
    .A2(net35),
    .A3(net649),
    .S0(net692),
    .S1(net875),
    .X(net412));
 sky130_fd_sc_hd__mux4_1 c604 (.A0(net832),
    .A1(net998),
    .A2(net904),
    .A3(net615),
    .S0(net616),
    .S1(net875),
    .X(net413));
 sky130_fd_sc_hd__mux4_1 c605 (.A0(net261),
    .A1(net932),
    .A2(net941),
    .A3(net75),
    .S0(net385),
    .S1(net1130),
    .X(net414));
 sky130_fd_sc_hd__mux4_1 c606 (.A0(net140),
    .A1(net60),
    .A2(net1057),
    .A3(net120),
    .S0(net1004),
    .S1(net894),
    .X(net415));
 sky130_fd_sc_hd__mux4_1 c607 (.A0(net976),
    .A1(clknet_1_1__leaf_net352),
    .A2(net616),
    .A3(net628),
    .S0(net629),
    .S1(net725),
    .X(net877));
 sky130_fd_sc_hd__mux4_1 c608 (.A0(net136),
    .A1(clknet_1_1__leaf_net342),
    .A2(clknet_1_0__leaf_net403),
    .A3(net684),
    .S0(clknet_1_1__leaf_net714),
    .S1(net730),
    .X(net416));
 sky130_fd_sc_hd__mux4_1 c609 (.A0(net413),
    .A1(net783),
    .A2(net406),
    .A3(clknet_1_0__leaf_net877),
    .S0(net615),
    .S1(net722),
    .X(net417));
 sky130_fd_sc_hd__mux4_1 c610 (.A0(net57),
    .A1(clknet_1_0__leaf_net877),
    .A2(net959),
    .A3(clknet_1_1__leaf_net407),
    .S0(net605),
    .S1(net670),
    .X(net418));
 sky130_fd_sc_hd__mux4_1 c611 (.A0(net940),
    .A1(clknet_1_0__leaf_net877),
    .A2(net406),
    .A3(net832),
    .S0(net642),
    .S1(net981),
    .X(net419));
 sky130_fd_sc_hd__mux4_1 c612 (.A0(net413),
    .A1(net789),
    .A2(net222),
    .A3(net604),
    .S0(net634),
    .S1(net730),
    .X(net420));
 sky130_fd_sc_hd__mux4_1 c613 (.A0(net1057),
    .A1(clknet_1_0__leaf_net407),
    .A2(net1017),
    .A3(net634),
    .S0(clknet_1_0__leaf_net643),
    .S1(net730),
    .X(net421));
 sky130_fd_sc_hd__mux4_1 c614 (.A0(net410),
    .A1(clknet_1_1__leaf_net352),
    .A2(net139),
    .A3(clknet_1_0__leaf_net877),
    .S0(net863),
    .S1(clknet_1_1__leaf_net693),
    .X(net422));
 sky130_fd_sc_hd__mux4_1 c615 (.A0(net422),
    .A1(net765),
    .A2(net406),
    .A3(net631),
    .S0(clknet_1_0__leaf_net643),
    .S1(net985),
    .X(net423));
 sky130_fd_sc_hd__mux4_2 c616 (.A0(net237),
    .A1(net903),
    .A2(net1005),
    .A3(net832),
    .S0(net629),
    .S1(net982),
    .X(net864));
 sky130_fd_sc_hd__mux4_1 c617 (.A0(net1050),
    .A1(net254),
    .A2(net800),
    .A3(net787),
    .S0(net864),
    .S1(net855),
    .X(net876));
 sky130_fd_sc_hd__mux4_1 c618 (.A0(net331),
    .A1(net57),
    .A2(net139),
    .A3(net844),
    .S0(net810),
    .S1(net652),
    .X(net424));
 sky130_fd_sc_hd__mux4_1 c619 (.A0(net41),
    .A1(clknet_1_0__leaf_net316),
    .A2(net961),
    .A3(net916),
    .S0(net717),
    .S1(net731),
    .X(net425));
 sky130_fd_sc_hd__mux4_2 c620 (.A0(net783),
    .A1(net803),
    .A2(net1018),
    .A3(net1043),
    .S0(net663),
    .S1(net703),
    .X(net859));
 sky130_fd_sc_hd__mux4_1 c621 (.A0(net866),
    .A1(clknet_1_0__leaf_net877),
    .A2(net331),
    .A3(net916),
    .S0(net614),
    .S1(net881),
    .X(net426));
 sky130_fd_sc_hd__mux4_1 c622 (.A0(clknet_1_1__leaf_net319),
    .A1(net68),
    .A2(net805),
    .A3(net1009),
    .S0(net652),
    .S1(clknet_1_1__leaf_net695),
    .X(net427));
 sky130_fd_sc_hd__mux4_1 c623 (.A0(net1045),
    .A1(net873),
    .A2(net881),
    .A3(net639),
    .S0(net703),
    .S1(net726),
    .X(net428));
 sky130_fd_sc_hd__mux4_1 c624 (.A0(net120),
    .A1(net810),
    .A2(net146),
    .A3(net873),
    .S0(net682),
    .S1(clknet_1_0__leaf_net732),
    .X(net429));
 sky130_fd_sc_hd__mux4_1 c625 (.A0(net800),
    .A1(net864),
    .A2(net77),
    .A3(net726),
    .S0(clknet_1_0__leaf_net732),
    .S1(clknet_1_0__leaf_net733),
    .X(net430));
 sky130_fd_sc_hd__mux4_1 c626 (.A0(net956),
    .A1(net1008),
    .A2(net1000),
    .A3(net997),
    .S0(net637),
    .S1(net670),
    .X(net431));
 sky130_fd_sc_hd__mux4_1 c627 (.A0(net146),
    .A1(clknet_1_0__leaf_net429),
    .A2(net401),
    .A3(net616),
    .S0(net646),
    .S1(net852),
    .X(net432));
 sky130_fd_sc_hd__mux4_1 c628 (.A0(net389),
    .A1(net1018),
    .A2(net859),
    .A3(net872),
    .S0(net639),
    .S1(net902),
    .X(net433));
 sky130_fd_sc_hd__mux4_1 c629 (.A0(net961),
    .A1(net866),
    .A2(clknet_1_0__leaf_net316),
    .A3(net637),
    .S0(net652),
    .S1(net982),
    .X(net434));
 sky130_fd_sc_hd__mux4_1 c630 (.A0(net832),
    .A1(net431),
    .A2(net428),
    .A3(net631),
    .S0(net856),
    .S1(net731),
    .X(net435));
 sky130_fd_sc_hd__mux4_1 c631 (.A0(net330),
    .A1(net765),
    .A2(net284),
    .A3(net940),
    .S0(net1008),
    .S1(clknet_1_1__leaf_net734),
    .X(net436));
 sky130_fd_sc_hd__mux4_1 c632 (.A0(net99),
    .A1(net428),
    .A2(clknet_1_1__leaf_net203),
    .A3(net663),
    .S0(net671),
    .S1(clknet_1_0__leaf_net734),
    .X(net437));
 sky130_fd_sc_hd__mux4_1 c633 (.A0(net431),
    .A1(clknet_1_1__leaf_net319),
    .A2(net428),
    .A3(net856),
    .S0(net670),
    .S1(clknet_1_0__leaf_net734),
    .X(net438));
 sky130_fd_sc_hd__mux4_1 c634 (.A0(net401),
    .A1(net1107),
    .A2(net869),
    .A3(net431),
    .S0(net663),
    .S1(clknet_1_0__leaf_net733),
    .X(net439));
 sky130_fd_sc_hd__mux4_1 c635 (.A0(clknet_1_1__leaf_net316),
    .A1(net858),
    .A2(net254),
    .A3(net1000),
    .S0(net630),
    .S1(net703),
    .X(net440));
 sky130_fd_sc_hd__mux4_1 c636 (.A0(net789),
    .A1(net934),
    .A2(net331),
    .A3(net853),
    .S0(net630),
    .S1(net639),
    .X(net441));
 sky130_fd_sc_hd__a41o_1 c637 (.A1(clknet_1_1__leaf_net203),
    .A2(net77),
    .A3(net853),
    .A4(net717),
    .B1(net735),
    .X(net442));
 sky130_fd_sc_hd__a41o_1 c660 (.A1(clknet_1_1__leaf_net250),
    .A2(net1022),
    .A3(clknet_1_1__leaf_net341),
    .A4(net979),
    .B1(net938),
    .X(net443));
 sky130_fd_sc_hd__mux4_1 c661 (.A0(net356),
    .A1(net938),
    .A2(net1133),
    .A3(clknet_1_0__leaf_net342),
    .S0(net946),
    .S1(net1016),
    .X(net444));
 sky130_fd_sc_hd__mux4_1 c662 (.A0(net233),
    .A1(net1022),
    .A2(net1096),
    .A3(clknet_1_0__leaf_net443),
    .S0(net127),
    .S1(net968),
    .X(net445));
 sky130_fd_sc_hd__a41o_1 c663 (.A1(net336),
    .A2(net335),
    .A3(clknet_1_0__leaf_net250),
    .A4(net996),
    .B1(net234),
    .X(net446));
 sky130_fd_sc_hd__a41o_1 c664 (.A1(net996),
    .A2(clknet_1_0__leaf_net444),
    .A3(clknet_1_0__leaf_net446),
    .A4(net938),
    .B1(net707),
    .X(net447));
 sky130_fd_sc_hd__a41o_1 c665 (.A1(net934),
    .A2(net1118),
    .A3(net1082),
    .A4(net232),
    .B1(net562),
    .X(net448));
 sky130_fd_sc_hd__sdfbbp_1 c666 (.CLK(clknet_4_5_0_clk),
    .D(net448),
    .RESET_B(net1097),
    .SCD(net938),
    .SCE(net976),
    .SET_B(net738),
    .Q(net450),
    .Q_N(net449));
 sky130_fd_sc_hd__a41o_1 c667 (.A1(net127),
    .A2(clknet_1_0__leaf_net352),
    .A3(net1020),
    .A4(net449),
    .B1(clknet_1_0__leaf_net675),
    .X(net451));
 sky130_fd_sc_hd__mux4_1 c668 (.A0(net938),
    .A1(net996),
    .A2(net959),
    .A3(net448),
    .S0(clknet_1_0__leaf_net451),
    .S1(net738),
    .X(net452));
 sky130_fd_sc_hd__sdfbbn_1 c669 (.CLK_N(clknet_4_4_0_clk),
    .D(clknet_1_1__leaf_net246),
    .RESET_B(net235),
    .SCD(net334),
    .SCE(net562),
    .SET_B(net739),
    .Q(net454),
    .Q_N(net453));
 sky130_fd_sc_hd__mux4_1 c670 (.A0(net450),
    .A1(net959),
    .A2(net1005),
    .A3(clknet_1_0__leaf_net451),
    .S0(net127),
    .S1(net938),
    .X(net455));
 sky130_fd_sc_hd__mux4_1 c671 (.A0(clknet_1_0__leaf_net444),
    .A1(net1016),
    .A2(net1012),
    .A3(net453),
    .S0(clknet_1_1__leaf_net250),
    .S1(clknet_1_1__leaf_net673),
    .X(net456));
 sky130_fd_sc_hd__a41o_1 c672 (.A1(clknet_1_0__leaf_net455),
    .A2(clknet_1_0__leaf_net456),
    .A3(net127),
    .A4(net1016),
    .B1(net740),
    .X(net457));
 sky130_fd_sc_hd__a41o_1 c673 (.A1(net340),
    .A2(clknet_1_0__leaf_net455),
    .A3(clknet_1_0__leaf_net457),
    .A4(clknet_1_0__leaf_net446),
    .B1(net739),
    .X(net458));
 sky130_fd_sc_hd__sdfbbn_1 c674 (.CLK_N(clknet_4_5_0_clk),
    .D(clknet_1_0__leaf_net458),
    .RESET_B(clknet_1_0__leaf_net457),
    .SCD(net975),
    .SCE(net939),
    .SET_B(net1002),
    .Q(net460),
    .Q_N(net459));
 sky130_fd_sc_hd__mux4_1 c675 (.A0(net448),
    .A1(net959),
    .A2(clknet_1_0__leaf_net457),
    .A3(net450),
    .S0(net460),
    .S1(net1020),
    .X(net461));
 sky130_fd_sc_hd__mux4_1 c676 (.A0(net346),
    .A1(clknet_1_0__leaf_net458),
    .A2(clknet_1_0__leaf_net455),
    .A3(clknet_1_0__leaf_net352),
    .S0(clknet_1_0__leaf_net443),
    .S1(net1007),
    .X(net462));
 sky130_fd_sc_hd__mux4_1 c677 (.A0(clknet_1_1__leaf_net456),
    .A1(net460),
    .A2(clknet_1_0__leaf_net457),
    .A3(net952),
    .S0(net740),
    .S1(net742),
    .X(net463));
 sky130_fd_sc_hd__sdfbbp_1 c678 (.CLK(clknet_4_5_0_clk),
    .D(clknet_1_1__leaf_net443),
    .RESET_B(clknet_1_1__leaf_net463),
    .SCD(net459),
    .SCE(net936),
    .SET_B(net739),
    .Q(net465),
    .Q_N(net464));
 sky130_fd_sc_hd__mux4_1 c679 (.A0(net946),
    .A1(clknet_1_1__leaf_net444),
    .A2(clknet_1_0__leaf_net463),
    .A3(net464),
    .S0(net459),
    .S1(net449),
    .X(net466));
 sky130_fd_sc_hd__mux4_1 c680 (.A0(clknet_1_0__leaf_net463),
    .A1(clknet_1_1__leaf_net458),
    .A2(net464),
    .A3(net459),
    .S0(net562),
    .X(net467));
 sky130_fd_sc_hd__mux4_1 c681 (.A0(clknet_1_0__leaf_net455),
    .A1(clknet_1_1__leaf_net463),
    .A2(net465),
    .A3(clknet_1_0__leaf_net457),
    .S0(net459),
    .S1(net737),
    .X(net468));
 sky130_fd_sc_hd__mux4_1 c682 (.A0(clknet_1_1__leaf_net451),
    .A1(clknet_1_0__leaf_net358),
    .A2(net225),
    .A3(net1133),
    .S0(net1025),
    .S1(net739),
    .X(net469));
 sky130_fd_sc_hd__mux4_1 c683 (.A0(net1038),
    .A1(net777),
    .A2(net1077),
    .A3(net234),
    .S0(net954),
    .S1(net709),
    .X(net470));
 sky130_fd_sc_hd__mux4_1 c684 (.A0(net151),
    .A1(net1118),
    .A2(net979),
    .A3(net573),
    .S0(clknet_1_0__leaf_net714),
    .S1(net741),
    .X(net471));
 sky130_fd_sc_hd__mux4_1 c685 (.A0(clknet_1_1__leaf_net341),
    .A1(net465),
    .A2(net460),
    .A3(net1079),
    .S0(net1031),
    .S1(net709),
    .X(net472));
 sky130_fd_sc_hd__mux4_1 c686 (.A0(net1016),
    .A1(net1019),
    .A2(net1116),
    .A3(clknet_1_0__leaf_net469),
    .S0(net238),
    .S1(net684),
    .X(net473));
 sky130_fd_sc_hd__mux4_1 c687 (.A0(net460),
    .A1(net465),
    .A2(net683),
    .A3(net711),
    .S0(net720),
    .S1(net743),
    .X(net474));
 sky130_fd_sc_hd__mux4_1 c688 (.A0(net1002),
    .A1(net1020),
    .A2(net777),
    .A3(net151),
    .S0(net464),
    .S1(net757),
    .X(net475));
 sky130_fd_sc_hd__mux4_1 c689 (.A0(net465),
    .A1(net1019),
    .A2(net459),
    .A3(net1009),
    .S0(net711),
    .S1(net740),
    .X(net476));
 sky130_fd_sc_hd__mux4_1 c690 (.A0(net952),
    .A1(net938),
    .A2(net1110),
    .A3(net965),
    .S0(net476),
    .S1(net742),
    .X(net477));
 sky130_fd_sc_hd__mux4_1 c691 (.A0(net1016),
    .A1(net1000),
    .A2(net561),
    .A3(net573),
    .S0(net707),
    .S1(net745),
    .X(net478));
 sky130_fd_sc_hd__mux4_1 c692 (.A0(net39),
    .A1(net752),
    .A2(clknet_1_0__leaf_net447),
    .A3(net334),
    .S0(net684),
    .S1(net741),
    .X(net479));
 sky130_fd_sc_hd__mux4_1 c693 (.A0(net345),
    .A1(net234),
    .A2(net1020),
    .A3(net711),
    .S0(net742),
    .S1(net746),
    .X(net480));
 sky130_fd_sc_hd__mux4_1 c694 (.A0(clknet_1_1__leaf_net446),
    .A1(net476),
    .A2(net996),
    .A3(net1012),
    .S0(net1018),
    .S1(net745),
    .X(net481));
 sky130_fd_sc_hd__mux4_1 c695 (.A0(net477),
    .A1(clknet_1_1__leaf_net366),
    .A2(net1025),
    .A3(net740),
    .S0(net745),
    .S1(net746),
    .X(net482));
 sky130_fd_sc_hd__mux4_1 c696 (.A0(net478),
    .A1(net777),
    .A2(net683),
    .A3(net710),
    .S0(net741),
    .S1(net746),
    .X(net483));
 sky130_fd_sc_hd__mux4_1 c697 (.A0(net480),
    .A1(clknet_1_0__leaf_net357),
    .A2(net1025),
    .A3(net1118),
    .S0(net741),
    .S1(net747),
    .X(net484));
 sky130_fd_sc_hd__mux4_1 c698 (.A0(net483),
    .A1(clknet_1_0__leaf_net469),
    .A2(clknet_1_0__leaf_net457),
    .A3(net464),
    .S0(net708),
    .S1(net746),
    .X(net485));
 sky130_fd_sc_hd__mux4_1 c699 (.A0(net270),
    .A1(net484),
    .A2(clknet_1_1__leaf_net366),
    .A3(net153),
    .S0(net1162),
    .S1(clknet_1_1__leaf_net675),
    .X(net486));
 sky130_fd_sc_hd__mux4_1 c700 (.A0(net151),
    .A1(net1034),
    .A2(net225),
    .A3(net744),
    .S0(net745),
    .S1(net747),
    .X(net487));
 sky130_fd_sc_hd__mux4_1 c701 (.A0(clknet_1_0__leaf_net455),
    .A1(net465),
    .A2(net480),
    .A3(net474),
    .S0(net620),
    .S1(net740),
    .X(net488));
 sky130_fd_sc_hd__mux4_1 c702 (.A0(net488),
    .A1(net460),
    .A2(net335),
    .A3(net785),
    .S0(net1009),
    .S1(net620),
    .X(net489));
 sky130_fd_sc_hd__mux4_1 c703 (.A0(net470),
    .A1(net153),
    .A2(net1019),
    .A3(net584),
    .S0(net709),
    .S1(net744),
    .X(net490));
 sky130_fd_sc_hd__mux4_1 c704 (.A0(net472),
    .A1(net1133),
    .A2(net238),
    .A3(net1116),
    .S0(net385),
    .S1(net708),
    .X(net491));
 sky130_fd_sc_hd__mux4_1 c705 (.A0(clknet_1_0__leaf_net358),
    .A1(net39),
    .A2(net454),
    .A3(net721),
    .S0(net723),
    .S1(net729),
    .X(net492));
 sky130_fd_sc_hd__mux4_1 c706 (.A0(net1018),
    .A1(net1056),
    .A2(net803),
    .A3(net768),
    .S0(net791),
    .S1(net580),
    .X(net493));
 sky130_fd_sc_hd__mux4_1 c707 (.A0(net788),
    .A1(net385),
    .A2(net163),
    .A3(net584),
    .S0(net984),
    .S1(net981),
    .X(net494));
 sky130_fd_sc_hd__mux4_1 c708 (.A0(net284),
    .A1(clknet_1_1__leaf_net675),
    .A2(net723),
    .A3(net724),
    .S0(net748),
    .S1(net750),
    .X(net495));
 sky130_fd_sc_hd__mux4_1 c709 (.A0(clknet_1_1__leaf_net457),
    .A1(net777),
    .A2(net788),
    .A3(clknet_1_0__leaf_net495),
    .S0(net580),
    .S1(net746),
    .X(net496));
 sky130_fd_sc_hd__mux4_1 c710 (.A0(clknet_1_1__leaf_net447),
    .A1(net288),
    .A2(net786),
    .A3(net984),
    .S0(clknet_1_1__leaf_net675),
    .S1(clknet_1_0__leaf_net714),
    .X(net497));
 sky130_fd_sc_hd__mux4_1 c711 (.A0(net788),
    .A1(net34),
    .A2(net976),
    .A3(net68),
    .S0(net723),
    .S1(net748),
    .X(net498));
 sky130_fd_sc_hd__a41o_1 c712 (.A1(clknet_1_1__leaf_net455),
    .A2(net284),
    .A3(net39),
    .A4(net580),
    .B1(net686),
    .X(net499));
 sky130_fd_sc_hd__mux4_1 c713 (.A0(net968),
    .A1(net396),
    .A2(clknet_1_0__leaf_net499),
    .A3(net561),
    .S0(net709),
    .S1(net728),
    .X(net500));
 sky130_fd_sc_hd__mux4_1 c714 (.A0(net153),
    .A1(net335),
    .A2(net791),
    .A3(clknet_1_1__leaf_net457),
    .S0(net257),
    .S1(net942),
    .X(net501));
 sky130_fd_sc_hd__mux4_1 c715 (.A0(net454),
    .A1(net194),
    .A2(clknet_1_0__leaf_net499),
    .A3(net723),
    .S0(net726),
    .S1(net748),
    .X(net502));
 sky130_fd_sc_hd__mux4_1 c716 (.A0(net1083),
    .A1(net788),
    .A2(net334),
    .A3(net453),
    .S0(net855),
    .S1(net860),
    .X(net503));
 sky130_fd_sc_hd__mux4_1 c717 (.A0(net979),
    .A1(net803),
    .A2(clknet_1_1__leaf_net495),
    .A3(net677),
    .S0(net682),
    .S1(net691),
    .X(net504));
 sky130_fd_sc_hd__mux4_1 c718 (.A0(clknet_1_1__leaf_net502),
    .A1(clknet_1_1__leaf_net455),
    .A2(clknet_1_0__leaf_net714),
    .A3(net728),
    .S0(net743),
    .S1(net748),
    .X(net505));
 sky130_fd_sc_hd__mux4_1 c719 (.A0(clknet_1_1__leaf_net443),
    .A1(clknet_1_0__leaf_net502),
    .A2(net1116),
    .A3(net757),
    .S0(net683),
    .S1(net723),
    .X(net506));
 sky130_fd_sc_hd__mux4_1 c720 (.A0(net496),
    .A1(clknet_1_0__leaf_net502),
    .A2(net975),
    .A3(net624),
    .S0(net727),
    .S1(net860),
    .X(net507));
 sky130_fd_sc_hd__mux4_1 c721 (.A0(net763),
    .A1(clknet_1_1__leaf_net358),
    .A2(clknet_1_0__leaf_net495),
    .A3(net760),
    .S0(net1000),
    .S1(net620),
    .X(net508));
 sky130_fd_sc_hd__mux4_1 c722 (.A0(net474),
    .A1(clknet_1_0__leaf_net492),
    .A2(net1109),
    .A3(net760),
    .S0(net624),
    .S1(net690),
    .X(net509));
 sky130_fd_sc_hd__mux4_1 c723 (.A0(clknet_1_0__leaf_net492),
    .A1(clknet_1_1__leaf_net502),
    .A2(clknet_1_1__leaf_net457),
    .A3(net1101),
    .S0(net677),
    .S1(net749),
    .X(net510));
 sky130_fd_sc_hd__mux4_1 c724 (.A0(net503),
    .A1(net388),
    .A2(net1084),
    .A3(clknet_1_0__leaf_net492),
    .S0(clknet_1_0__leaf_net499),
    .S1(net750),
    .X(net511));
 sky130_fd_sc_hd__mux4_1 c725 (.A0(net511),
    .A1(net163),
    .A2(clknet_1_0__leaf_net499),
    .A3(net665),
    .S0(net711),
    .S1(net750),
    .X(net512));
 sky130_fd_sc_hd__mux4_1 c726 (.A0(net504),
    .A1(net832),
    .A2(net959),
    .A3(clknet_1_1__leaf_net675),
    .S0(net981),
    .S1(net721),
    .X(net513));
 sky130_fd_sc_hd__mux4_1 c727 (.A0(net189),
    .A1(net786),
    .A2(clknet_1_1__leaf_net352),
    .A3(net670),
    .S0(net744),
    .S1(net751),
    .X(net514));
 sky130_fd_sc_hd__mux4_1 c728 (.A0(net959),
    .A1(net952),
    .A2(net239),
    .A3(net385),
    .S0(net665),
    .S1(net710),
    .X(net515));
 sky130_fd_sc_hd__mux4_2 c729 (.A0(net396),
    .A1(net508),
    .A2(clknet_1_0__leaf_net481),
    .A3(net235),
    .S0(net947),
    .S1(net1004),
    .X(net516));
 sky130_fd_sc_hd__mux4_1 c730 (.A0(clknet_1_1__leaf_net352),
    .A1(net1060),
    .A2(net791),
    .A3(net297),
    .S0(net239),
    .S1(clknet_1_0__leaf_net509),
    .X(net517));
 sky130_fd_sc_hd__mux4_1 c731 (.A0(net77),
    .A1(clknet_1_1__leaf_net492),
    .A2(net824),
    .A3(clknet_1_1__leaf_net499),
    .S0(net65),
    .S1(net610),
    .X(net518));
 sky130_fd_sc_hd__mux4_1 c732 (.A0(clknet_1_1__leaf_net492),
    .A1(net854),
    .A2(net297),
    .A3(net642),
    .S0(net670),
    .S1(net684),
    .X(net519));
 sky130_fd_sc_hd__mux4_1 c733 (.A0(net194),
    .A1(net181),
    .A2(net824),
    .A3(net420),
    .S0(net786),
    .S1(net1030),
    .X(net520));
 sky130_fd_sc_hd__mux4_1 c734 (.A0(net777),
    .A1(net1056),
    .A2(clknet_1_1__leaf_net509),
    .A3(net976),
    .S0(clknet_1_1__leaf_net499),
    .S1(clknet_1_1__leaf_net913),
    .X(net521));
 sky130_fd_sc_hd__mux4_1 c735 (.A0(clknet_1_1__leaf_net489),
    .A1(net62),
    .A2(clknet_1_1__leaf_net469),
    .A3(clknet_1_0__leaf_net913),
    .S0(net721),
    .S1(net751),
    .X(net522));
 sky130_fd_sc_hd__mux4_1 c736 (.A0(net1018),
    .A1(net824),
    .A2(clknet_1_1__leaf_net352),
    .A3(net570),
    .S0(net645),
    .S1(net747),
    .X(net523));
 sky130_fd_sc_hd__mux4_1 c737 (.A0(net50),
    .A1(net1077),
    .A2(net570),
    .A3(net640),
    .S0(net710),
    .S1(net751),
    .X(net524));
 sky130_fd_sc_hd__mux4_1 c738 (.A0(net385),
    .A1(net83),
    .A2(net225),
    .A3(net295),
    .S0(net1131),
    .S1(net1126),
    .X(net525));
 sky130_fd_sc_hd__mux4_1 c739 (.A0(net1078),
    .A1(clknet_1_1__leaf_net403),
    .A2(net478),
    .A3(net1060),
    .S0(net239),
    .S1(net640),
    .X(net526));
 sky130_fd_sc_hd__mux4_1 c740 (.A0(clknet_1_1__leaf_net877),
    .A1(clknet_1_1__leaf_net310),
    .A2(net194),
    .A3(net863),
    .S0(net642),
    .S1(net645),
    .X(net527));
 sky130_fd_sc_hd__mux4_1 c741 (.A0(net194),
    .A1(net1087),
    .A2(net965),
    .A3(net627),
    .S0(clknet_1_1__leaf_net643),
    .S1(net670),
    .X(net528));
 sky130_fd_sc_hd__mux4_1 c742 (.A0(clknet_1_0__leaf_net528),
    .A1(clknet_1_1__leaf_net495),
    .A2(clknet_1_1__leaf_net527),
    .A3(net824),
    .S0(net665),
    .S1(net743),
    .X(net529));
 sky130_fd_sc_hd__mux4_1 c743 (.A0(clknet_1_1__leaf_net481),
    .A1(net65),
    .A2(net858),
    .A3(clknet_1_0__leaf_net527),
    .S0(clknet_1_0__leaf_net528),
    .S1(net952),
    .X(net530));
 sky130_fd_sc_hd__mux4_1 c744 (.A0(clknet_1_0__leaf_net509),
    .A1(clknet_1_0__leaf_net523),
    .A2(clknet_1_1__leaf_net528),
    .A3(clknet_1_1__leaf_net499),
    .S0(net570),
    .S1(net855),
    .X(net531));
 sky130_fd_sc_hd__mux4_1 c745 (.A0(net531),
    .A1(net1033),
    .A2(clknet_1_1__leaf_net528),
    .A3(clknet_1_1__leaf_net352),
    .S0(net385),
    .S1(net751),
    .X(net532));
 sky130_fd_sc_hd__mux4_2 c746 (.A0(net295),
    .A1(net420),
    .A2(clknet_1_1__leaf_net523),
    .A3(clknet_1_1__leaf_net528),
    .S0(net641),
    .S1(net856),
    .X(net533));
 sky130_fd_sc_hd__mux4_1 c747 (.A0(clknet_1_1__leaf_net499),
    .A1(clknet_1_0__leaf_net489),
    .A2(net1049),
    .A3(net936),
    .S0(net1101),
    .S1(net610),
    .X(net534));
 sky130_fd_sc_hd__mux4_1 c748 (.A0(net782),
    .A1(net514),
    .A2(net53),
    .A3(net704),
    .S0(net855),
    .S1(clknet_1_1__leaf_net733),
    .X(net535));
 sky130_fd_sc_hd__mux4_2 c749 (.A0(net1000),
    .A1(net533),
    .A2(net997),
    .A3(net844),
    .S0(net623),
    .S1(net704),
    .X(net536));
 sky130_fd_sc_hd__mux4_1 c750 (.A0(clknet_1_1__leaf_net357),
    .A1(net1108),
    .A2(net68),
    .A3(net524),
    .S0(net976),
    .S1(net622),
    .X(net537));
 sky130_fd_sc_hd__mux4_1 c751 (.A0(net225),
    .A1(net791),
    .A2(net785),
    .A3(net1004),
    .S0(net984),
    .S1(net717),
    .X(net538));
 sky130_fd_sc_hd__mux4_1 c752 (.A0(net493),
    .A1(net1088),
    .A2(net947),
    .A3(net614),
    .S0(net646),
    .S1(net736),
    .X(net539));
 sky130_fd_sc_hd__mux4_1 c753 (.A0(net1060),
    .A1(clknet_1_1__leaf_net357),
    .A2(net803),
    .A3(net622),
    .S0(net633),
    .S1(clknet_1_1__leaf_net714),
    .X(net540));
 sky130_fd_sc_hd__mux4_1 c754 (.A0(net257),
    .A1(net976),
    .A2(clknet_1_1__leaf_net429),
    .A3(clknet_1_1__leaf_net521),
    .S0(net524),
    .S1(net749),
    .X(net541));
 sky130_fd_sc_hd__mux4_1 c755 (.A0(net19),
    .A1(net284),
    .A2(clknet_1_1__leaf_net469),
    .A3(net774),
    .S0(net760),
    .S1(net692),
    .X(net542));
 sky130_fd_sc_hd__mux4_1 c756 (.A0(net53),
    .A1(clknet_1_0__leaf_net521),
    .A2(net760),
    .A3(net844),
    .S0(net670),
    .S1(net852),
    .X(net543));
 sky130_fd_sc_hd__mux4_1 c757 (.A0(net1029),
    .A1(net775),
    .A2(net623),
    .A3(net640),
    .S0(net985),
    .S1(net749),
    .X(net544));
 sky130_fd_sc_hd__mux4_1 c758 (.A0(net297),
    .A1(net786),
    .A2(net1041),
    .A3(net29),
    .S0(net627),
    .S1(net638),
    .X(net545));
 sky130_fd_sc_hd__mux4_1 c759 (.A0(net791),
    .A1(net406),
    .A2(net540),
    .A3(net757),
    .S0(net665),
    .S1(net731),
    .X(net546));
 sky130_fd_sc_hd__mux4_1 c760 (.A0(net757),
    .A1(net29),
    .A2(net626),
    .A3(net863),
    .S0(net984),
    .S1(net731),
    .X(net547));
 sky130_fd_sc_hd__mux4_1 c761 (.A0(net235),
    .A1(net1002),
    .A2(net547),
    .A3(net544),
    .S0(net19),
    .S1(net625),
    .X(net548));
 sky130_fd_sc_hd__mux4_1 c762 (.A0(net1004),
    .A1(net539),
    .A2(net1108),
    .A3(net638),
    .S0(net655),
    .S1(net725),
    .X(net549));
 sky130_fd_sc_hd__mux4_1 c763 (.A0(clknet_1_1__leaf_net310),
    .A1(net62),
    .A2(net548),
    .A3(net997),
    .S0(net690),
    .S1(net704),
    .X(net550));
 sky130_fd_sc_hd__mux4_1 c764 (.A0(clknet_1_1__leaf_net342),
    .A1(net796),
    .A2(net406),
    .A3(net665),
    .S0(net692),
    .S1(net743),
    .X(net551));
 sky130_fd_sc_hd__mux4_1 c765 (.A0(net239),
    .A1(net77),
    .A2(net610),
    .A3(net633),
    .S0(net640),
    .S1(net747),
    .X(net552));
 sky130_fd_sc_hd__mux4_1 c766 (.A0(net549),
    .A1(net832),
    .A2(net535),
    .A3(net550),
    .S0(net68),
    .S1(net625),
    .X(net553));
 sky130_fd_sc_hd__mux4_1 c767 (.A0(clknet_1_1__leaf_net203),
    .A1(net538),
    .A2(net626),
    .A3(net638),
    .S0(net642),
    .S1(net747),
    .X(net554));
 sky130_fd_sc_hd__a41o_1 c768 (.A1(net785),
    .A2(net529),
    .A3(net641),
    .A4(clknet_1_1__leaf_net643),
    .B1(clknet_1_1__leaf_net732),
    .X(net555));
 sky130_fd_sc_hd__a41o_1 c769 (.A1(net50),
    .A2(net34),
    .A3(net627),
    .A4(clknet_1_0__leaf_net913),
    .B1(net682));
 sky130_fd_sc_hd__xnor2_1 merge790 (.A(net425),
    .B(net432),
    .Y(net556));
 sky130_fd_sc_hd__xnor2_1 merge791 (.A(net482),
    .B(net486),
    .Y(net557));
 sky130_fd_sc_hd__xnor2_1 merge792 (.A(net200),
    .B(net184),
    .Y(net558));
 sky130_fd_sc_hd__dfrbp_2 merge793 (.CLK(clknet_4_8_0_clk),
    .D(net86),
    .RESET_B(net88),
    .Q(net880),
    .Q_N(net559));
 sky130_fd_sc_hd__xnor2_1 merge794 (.A(net513),
    .B(net515),
    .Y(net560));
 sky130_fd_sc_hd__dfrbp_2 merge795 (.CLK(clknet_4_4_0_clk),
    .D(net337),
    .RESET_B(net338),
    .Q(net562),
    .Q_N(net561));
 sky130_fd_sc_hd__xnor2_1 merge796 (.A(net381),
    .B(net362),
    .Y(net563));
 sky130_fd_sc_hd__xnor2_1 merge797 (.A(net315),
    .B(net320),
    .Y(net564));
 sky130_fd_sc_hd__xnor2_1 merge798 (.A(net404),
    .B(net405),
    .Y(net565));
 sky130_fd_sc_hd__dfrtn_1 merge799 (.CLK_N(clknet_4_8_0_clk),
    .D(net171),
    .RESET_B(net176),
    .Q(net566));
 sky130_fd_sc_hd__xnor2_1 merge800 (.A(net152),
    .B(net159),
    .Y(net567));
 sky130_fd_sc_hd__dfrtp_1 merge801 (.CLK(clknet_4_9_0_clk),
    .D(net296),
    .RESET_B(net300),
    .Q(net568));
 sky130_fd_sc_hd__xnor2_1 merge802 (.A(net208),
    .B(net209),
    .Y(net569));
 sky130_fd_sc_hd__dfrtp_1 merge803 (.CLK(clknet_4_5_0_clk),
    .D(net466),
    .Q(net467));
 sky130_fd_sc_hd__xnor2_1 merge804 (.A(net71),
    .B(net64),
    .Y(net571));
 sky130_fd_sc_hd__xnor2_1 merge805 (.A(net113),
    .B(net115),
    .Y(net572));
 sky130_fd_sc_hd__dfrtp_4 merge806 (.CLK(clknet_4_0_0_clk),
    .D(net259),
    .RESET_B(net266),
    .Q(net573));
 sky130_fd_sc_hd__xnor2_1 merge807 (.A(net494),
    .B(net497),
    .Y(net574));
 sky130_fd_sc_hd__dfsbp_2 merge808 (.CLK(clknet_4_1_0_clk),
    .D(net249),
    .SET_B(net243),
    .Q(net576),
    .Q_N(net575));
 sky130_fd_sc_hd__dfsbp_1 merge809 (.CLK(clknet_4_10_0_clk),
    .D(net104),
    .SET_B(net111),
    .Q(net577),
    .Q_N(net910));
 sky130_fd_sc_hd__xnor2_2 merge810 (.A(net536),
    .B(net537),
    .Y(net578));
 sky130_fd_sc_hd__xnor2_1 merge811 (.A(net279),
    .B(net283),
    .Y(net579));
 sky130_fd_sc_hd__dfstp_1 merge812 (.CLK(clknet_4_6_0_clk),
    .D(net402),
    .SET_B(net383),
    .Q(net865));
 sky130_fd_sc_hd__dfstp_1 merge813 (.CLK(clknet_4_5_0_clk),
    .D(net485),
    .SET_B(net468),
    .Q(net580));
 sky130_fd_sc_hd__dfstp_1 merge814 (.CLK(clknet_4_0_0_clk),
    .D(net144),
    .Q(net147));
 sky130_fd_sc_hd__dlrbn_1 merge815 (.D(net89),
    .GATE_N(clknet_4_8_0_clk),
    .RESET_B(net84),
    .Q(net583),
    .Q_N(net582));
 sky130_fd_sc_hd__dlrbn_1 merge816 (.D(net368),
    .GATE_N(clknet_4_5_0_clk),
    .RESET_B(net557),
    .Q(net585),
    .Q_N(net584));
 sky130_fd_sc_hd__xnor2_1 merge817 (.A(net219),
    .B(net217),
    .Y(net586));
 sky130_fd_sc_hd__dlrbp_2 merge818 (.GATE(clknet_4_9_0_clk),
    .RESET_B(net558),
    .Q(net904),
    .Q_N(net199));
 sky130_fd_sc_hd__xnor2_1 merge819 (.A(net408),
    .B(net442),
    .Y(net588));
 sky130_fd_sc_hd__dlrbp_1 merge820 (.D(net112),
    .GATE(clknet_4_11_0_clk),
    .RESET_B(net572),
    .Q(net867),
    .Q_N(net930));
 sky130_fd_sc_hd__dlrtn_2 merge821 (.D(net94),
    .GATE_N(clknet_4_10_0_clk),
    .RESET_B(net106),
    .Q(net916));
 sky130_fd_sc_hd__dlrtn_2 merge822 (.D(net110),
    .GATE_N(clknet_4_10_0_clk),
    .RESET_B(net87),
    .Q(net589));
 sky130_fd_sc_hd__dlrtn_1 merge823 (.D(net398),
    .GATE_N(clknet_4_6_0_clk),
    .RESET_B(net289),
    .Q(net590));
 sky130_fd_sc_hd__dlrtp_1 merge824 (.GATE(clknet_4_8_0_clk),
    .RESET_B(net571),
    .Q(net69));
 sky130_fd_sc_hd__xnor2_1 merge825 (.A(net322),
    .B(net332),
    .Y(net591));
 sky130_fd_sc_hd__xnor2_1 merge826 (.A(net586),
    .B(net211),
    .Y(net592));
 sky130_fd_sc_hd__xnor2_1 merge827 (.A(net323),
    .B(net326),
    .Y(net593));
 sky130_fd_sc_hd__xnor2_1 merge828 (.A(net416),
    .B(net534),
    .Y(net594));
 sky130_fd_sc_hd__xnor2_1 merge829 (.A(net505),
    .B(net555),
    .Y(net595));
 sky130_fd_sc_hd__xnor2_1 merge830 (.A(net210),
    .B(net564),
    .Y(net596));
 sky130_fd_sc_hd__xnor2_1 merge831 (.A(net517),
    .B(net554),
    .Y(net597));
 sky130_fd_sc_hd__xnor2_1 merge832 (.A(net433),
    .B(net553),
    .Y(net598));
 sky130_fd_sc_hd__xnor2_1 merge833 (.A(net434),
    .B(net421),
    .Y(net599));
 sky130_fd_sc_hd__xnor2_1 merge834 (.A(net530),
    .B(net411),
    .Y(net600));
 sky130_fd_sc_hd__xnor2_1 merge835 (.A(net512),
    .B(net507),
    .Y(net601));
 sky130_fd_sc_hd__xnor2_1 merge836 (.A(net520),
    .B(net498),
    .Y(net602));
 sky130_fd_sc_hd__xnor2_1 merge837 (.A(net506),
    .B(net500),
    .Y(net603));
 sky130_fd_sc_hd__dlrtp_1 merge838 (.D(net414),
    .GATE(clknet_4_6_0_clk),
    .RESET_B(net291),
    .Q(net604));
 sky130_fd_sc_hd__dlrtp_2 merge839 (.D(net272),
    .GATE(clknet_4_1_0_clk),
    .RESET_B(net563),
    .Q(net605));
 sky130_fd_sc_hd__edfxbp_1 merge840 (.CLK(clknet_4_3_0_clk),
    .D(net271),
    .DE(net260),
    .Q(net607),
    .Q_N(net606));
 sky130_fd_sc_hd__edfxtp_1 merge841 (.CLK(clknet_4_2_0_clk),
    .D(net156),
    .DE(net567),
    .Q(net608));
 sky130_fd_sc_hd__xnor2_1 merge842 (.A(net436),
    .B(net437),
    .Y(net609));
 sky130_fd_sc_hd__sdlclkp_1 merge843 (.CLK(clknet_4_14_0_clk),
    .GATE(net593),
    .SCE(net301),
    .GCLK(net882));
 sky130_fd_sc_hd__sdlclkp_2 merge844 (.CLK(clknet_4_11_0_clk),
    .GATE(net207),
    .SCE(net218),
    .GCLK(net912));
 sky130_fd_sc_hd__sdlclkp_4 merge845 (.CLK(clknet_4_3_0_clk),
    .GATE(net290),
    .GCLK(net293));
 sky130_fd_sc_hd__xnor2_1 merge846 (.A(net518),
    .B(net552),
    .Y(net611));
 sky130_fd_sc_hd__dfrbp_2 merge847 (.CLK(clknet_4_12_0_clk),
    .D(net309),
    .RESET_B(net305),
    .Q(net894),
    .Q_N(net883));
 sky130_fd_sc_hd__xnor2_1 merge848 (.A(net532),
    .B(net551),
    .Y(net612));
 sky130_fd_sc_hd__xnor2_1 merge849 (.A(net440),
    .B(net438),
    .Y(net613));
 sky130_fd_sc_hd__dfrbp_1 merge850 (.CLK(clknet_4_13_0_clk),
    .D(net409),
    .RESET_B(net594),
    .Q(net615),
    .Q_N(net614));
 sky130_fd_sc_hd__dfrtn_1 merge851 (.CLK_N(clknet_4_14_0_clk),
    .D(net591),
    .RESET_B(net333),
    .Q(net881));
 sky130_fd_sc_hd__dfrtp_4 merge852 (.CLK(clknet_4_14_0_clk),
    .D(net303),
    .RESET_B(net312),
    .Q(net616));
 sky130_fd_sc_hd__xnor2_1 merge853 (.A(net569),
    .B(net321),
    .Y(net617));
 sky130_fd_sc_hd__xnor2_1 merge854 (.A(net542),
    .B(net546),
    .Y(net618));
 sky130_fd_sc_hd__xnor2_1 merge855 (.A(net545),
    .B(net541),
    .Y(net619));
 sky130_fd_sc_hd__dfrtp_4 merge856 (.CLK(clknet_4_7_0_clk),
    .D(net487),
    .RESET_B(net601),
    .Q(net620));
 sky130_fd_sc_hd__xnor2_1 merge857 (.A(net595),
    .B(net619),
    .Y(net621));
 sky130_fd_sc_hd__dfrtp_4 merge858 (.CLK(clknet_4_11_0_clk),
    .D(net592),
    .RESET_B(net215),
    .Q(net622));
 sky130_fd_sc_hd__dfsbp_1 merge859 (.CLK(clknet_4_7_0_clk),
    .D(net603),
    .SET_B(net574),
    .Q(net624),
    .Q_N(net623));
 sky130_fd_sc_hd__dfsbp_1 merge860 (.CLK(clknet_4_13_0_clk),
    .D(net618),
    .SET_B(net525),
    .Q(net626),
    .Q_N(net625));
 sky130_fd_sc_hd__dfstp_1 merge861 (.CLK(clknet_4_15_0_clk),
    .D(net613),
    .SET_B(net609),
    .Q(net853));
 sky130_fd_sc_hd__dfstp_2 merge862 (.CLK(clknet_4_6_0_clk),
    .D(net394),
    .SET_B(net621),
    .Q(net627));
 sky130_fd_sc_hd__dfstp_1 merge863 (.CLK(clknet_4_14_0_clk),
    .D(net314),
    .SET_B(net306),
    .Q(net628));
 sky130_fd_sc_hd__dlrbn_1 merge864 (.D(net439),
    .GATE_N(clknet_4_14_0_clk),
    .RESET_B(net412),
    .Q(net630),
    .Q_N(net629));
 sky130_fd_sc_hd__dlrbn_1 merge865 (.D(net565),
    .GATE_N(clknet_4_12_0_clk),
    .RESET_B(net599),
    .Q(net632),
    .Q_N(net631));
 sky130_fd_sc_hd__dlrbp_1 merge866 (.D(net417),
    .GATE(clknet_4_13_0_clk),
    .RESET_B(net578),
    .Q(net634),
    .Q_N(net633));
 sky130_fd_sc_hd__dlrbp_1 merge867 (.GATE(clknet_4_9_0_clk),
    .RESET_B(net192),
    .Q(net636),
    .Q_N(net635));
 sky130_fd_sc_hd__dlrtn_4 merge868 (.D(net579),
    .GATE_N(clknet_4_9_0_clk),
    .RESET_B(net287),
    .Q(net637));
 sky130_fd_sc_hd__dlrtn_1 merge869 (.D(net588),
    .GATE_N(clknet_4_15_0_clk),
    .RESET_B(net611),
    .Q(net638));
 sky130_fd_sc_hd__dlrtn_2 merge870 (.D(net116),
    .GATE_N(clknet_4_11_0_clk),
    .RESET_B(net596),
    .Q(net920));
 sky130_fd_sc_hd__dlrtp_1 merge871 (.GATE(clknet_4_11_0_clk),
    .RESET_B(net206),
    .Q(net221));
 sky130_fd_sc_hd__dlrtp_2 merge872 (.D(net418),
    .GATE(clknet_4_13_0_clk),
    .RESET_B(net602),
    .Q(net863));
 sky130_fd_sc_hd__dlrtp_1 merge873 (.D(net516),
    .GATE(clknet_4_7_0_clk),
    .RESET_B(net543),
    .Q(net640));
 sky130_fd_sc_hd__edfxbp_1 merge874 (.CLK(clknet_4_13_0_clk),
    .D(net612),
    .DE(net598),
    .Q(net641),
    .Q_N(net923));
 sky130_fd_sc_hd__edfxtp_1 merge875 (.CLK(clknet_4_13_0_clk),
    .D(net423),
    .DE(net600),
    .Q(net642));
 sky130_fd_sc_hd__sdlclkp_1 merge876 (.CLK(clknet_4_13_0_clk),
    .GATE(net597),
    .SCE(net419),
    .GCLK(net643));
 sky130_fd_sc_hd__sdlclkp_2 merge877 (.CLK(clknet_4_7_0_clk),
    .GATE(net560),
    .SCE(net519),
    .GCLK(net913));
 sky130_fd_sc_hd__sdlclkp_4 merge878 (.CLK(clknet_4_11_0_clk),
    .GATE(net204),
    .SCE(net202),
    .GCLK(net644));
 sky130_fd_sc_hd__dfrbp_1 merge879 (.CLK(clknet_4_15_0_clk),
    .D(net430),
    .RESET_B(net522),
    .Q(net646),
    .Q_N(net645));
 sky130_fd_sc_hd__dfrbp_2 merge880 (.CLK(clknet_4_8_0_clk),
    .D(net175),
    .RESET_B(net169),
    .Q(net647),
    .Q_N(net891));
 sky130_fd_sc_hd__dfrtn_1 merge881 (.CLK_N(clknet_4_15_0_clk),
    .D(net556),
    .RESET_B(net526),
    .Q(net856));
 sky130_fd_sc_hd__dfrtp_4 merge882 (.CLK(clknet_4_8_0_clk),
    .D(net91),
    .RESET_B(net617),
    .Q(net902));
 sky130_fd_sc_hd__dfrtp_4 merge883 (.CLK(clknet_4_6_0_clk),
    .D(net390),
    .RESET_B(net382),
    .Q(net648));
 sky130_fd_sc_hd__dfxbp_2 s884 (.CLK(clknet_4_2_0_clk),
    .D(net59),
    .Q(net650),
    .Q_N(net649));
 sky130_fd_sc_hd__dfxbp_2 s885 (.CLK(clknet_4_12_0_clk),
    .D(net70),
    .Q(net652),
    .Q_N(net651));
 sky130_fd_sc_hd__dfxtp_1 s886 (.CLK(clknet_4_8_0_clk),
    .D(net73),
    .Q(net653));
 sky130_fd_sc_hd__dfxtp_2 s887 (.CLK(clknet_4_10_0_clk),
    .D(net82),
    .Q(net654));
 sky130_fd_sc_hd__dfxtp_2 s888 (.CLK(clknet_4_10_0_clk),
    .D(net85),
    .Q(net655));
 sky130_fd_sc_hd__dlclkp_1 s889 (.CLK(clknet_4_8_0_clk),
    .GATE(net93),
    .GCLK(net656));
 sky130_fd_sc_hd__dlclkp_2 s890 (.CLK(clknet_4_10_0_clk),
    .GATE(net96),
    .GCLK(net657));
 sky130_fd_sc_hd__dlclkp_4 s891 (.CLK(clknet_4_10_0_clk),
    .GATE(net101),
    .GCLK(net658));
 sky130_fd_sc_hd__dlxbn_2 s892 (.D(net102),
    .GATE_N(clknet_4_11_0_clk),
    .Q(net870),
    .Q_N(net659));
 sky130_fd_sc_hd__dlxbn_1 s893 (.D(net103),
    .GATE_N(clknet_4_11_0_clk),
    .Q(net878),
    .Q_N(net660));
 sky130_fd_sc_hd__dlxbp_1 s894 (.D(net114),
    .GATE(clknet_4_10_0_clk),
    .Q(net662),
    .Q_N(net661));
 sky130_fd_sc_hd__dlxtn_4 s895 (.D(net155),
    .GATE_N(clknet_4_2_0_clk),
    .Q(net663));
 sky130_fd_sc_hd__dlxtn_1 s896 (.D(net170),
    .GATE_N(clknet_4_2_0_clk),
    .Q(net664));
 sky130_fd_sc_hd__dlxtn_4 s897 (.D(net173),
    .GATE_N(clknet_4_2_0_clk),
    .Q(net665));
 sky130_fd_sc_hd__dlxtp_1 s898 (.D(net185),
    .GATE(clknet_4_9_0_clk),
    .Q(net666));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s899 (.D(net186),
    .SLEEP_B(clknet_4_8_0_clk),
    .Q(net895));
 sky130_fd_sc_hd__dfxbp_1 s900 (.CLK(clknet_4_8_0_clk),
    .D(net187),
    .Q(net668),
    .Q_N(net667));
 sky130_fd_sc_hd__dfxbp_1 s901 (.CLK(clknet_4_9_0_clk),
    .D(net195),
    .Q(net889),
    .Q_N(net669));
 sky130_fd_sc_hd__dfxtp_4 s902 (.CLK(clknet_4_9_0_clk),
    .D(net198),
    .Q(net670));
 sky130_fd_sc_hd__dfxtp_1 s903 (.CLK(clknet_4_11_0_clk),
    .D(net214),
    .Q(net671));
 sky130_fd_sc_hd__dfxtp_1 s904 (.CLK(clknet_4_11_0_clk),
    .D(net220),
    .Q(net672));
 sky130_fd_sc_hd__dlclkp_1 s905 (.CLK(clknet_4_0_0_clk),
    .GATE(net242),
    .GCLK(net673));
 sky130_fd_sc_hd__dlclkp_2 s906 (.CLK(clknet_4_1_0_clk),
    .GATE(net244),
    .GCLK(net674));
 sky130_fd_sc_hd__dlclkp_4 s907 (.CLK(clknet_4_1_0_clk),
    .GATE(net245),
    .GCLK(net675));
 sky130_fd_sc_hd__dlxbn_1 s908 (.D(net251),
    .GATE_N(clknet_4_3_0_clk),
    .Q(net677),
    .Q_N(net676));
 sky130_fd_sc_hd__dlxbn_2 s909 (.D(net253),
    .GATE_N(clknet_4_0_0_clk),
    .Q(net679),
    .Q_N(net678));
 sky130_fd_sc_hd__dlxbp_1 s910 (.D(net258),
    .GATE(clknet_4_1_0_clk),
    .Q(net681),
    .Q_N(net680));
 sky130_fd_sc_hd__dlxtn_2 s911 (.D(net262),
    .GATE_N(clknet_4_2_0_clk),
    .Q(net682));
 sky130_fd_sc_hd__dlxtn_2 s912 (.D(net265),
    .GATE_N(clknet_4_3_0_clk),
    .Q(net683));
 sky130_fd_sc_hd__dlxtn_4 s913 (.D(net269),
    .GATE_N(clknet_4_1_0_clk),
    .Q(net684));
 sky130_fd_sc_hd__dlxtp_1 s914 (.D(net273),
    .GATE(clknet_4_3_0_clk),
    .Q(net685));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s915 (.D(net277),
    .SLEEP_B(clknet_4_3_0_clk),
    .Q(net686));
 sky130_fd_sc_hd__dfxbp_1 s916 (.CLK(clknet_4_9_0_clk),
    .D(net280),
    .Q(net893),
    .Q_N(net687));
 sky130_fd_sc_hd__dfxbp_1 s917 (.CLK(clknet_4_12_0_clk),
    .D(net281),
    .Q(net689),
    .Q_N(net688));
 sky130_fd_sc_hd__dfxtp_4 s918 (.CLK(clknet_4_3_0_clk),
    .D(net285),
    .Q(net690));
 sky130_fd_sc_hd__dfxtp_1 s919 (.CLK(clknet_4_3_0_clk),
    .D(net286),
    .Q(net691));
 sky130_fd_sc_hd__dfxtp_4 s920 (.CLK(clknet_4_3_0_clk),
    .D(net292),
    .Q(net692));
 sky130_fd_sc_hd__dlclkp_1 s921 (.CLK(clknet_4_12_0_clk),
    .GATE(net298),
    .GCLK(net693));
 sky130_fd_sc_hd__dlclkp_2 s922 (.CLK(clknet_4_12_0_clk),
    .GATE(net299),
    .GCLK(net694));
 sky130_fd_sc_hd__dlclkp_4 s923 (.CLK(clknet_4_12_0_clk),
    .GATE(net307),
    .GCLK(net695));
 sky130_fd_sc_hd__dlxbn_1 s924 (.D(net308),
    .GATE_N(clknet_4_12_0_clk),
    .Q(net697),
    .Q_N(net696));
 sky130_fd_sc_hd__dlxbn_1 s925 (.D(net311),
    .GATE_N(clknet_4_11_0_clk),
    .Q(net699),
    .Q_N(net698));
 sky130_fd_sc_hd__dlxbp_1 s926 (.D(net324),
    .GATE(clknet_4_14_0_clk),
    .Q(net701),
    .Q_N(net700));
 sky130_fd_sc_hd__dlxtn_1 s927 (.D(net327),
    .GATE_N(clknet_4_14_0_clk),
    .Q(net702));
 sky130_fd_sc_hd__dlxtn_1 s928 (.D(net328),
    .GATE_N(clknet_4_14_0_clk),
    .Q(net703));
 sky130_fd_sc_hd__dlxtn_1 s929 (.D(net329),
    .GATE_N(clknet_4_15_0_clk),
    .Q(net704));
 sky130_fd_sc_hd__dlxtp_1 s930 (.D(net344),
    .GATE(clknet_4_1_0_clk),
    .Q(net705));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s931 (.D(net354),
    .SLEEP_B(clknet_4_4_0_clk),
    .Q(net706));
 sky130_fd_sc_hd__dfxbp_1 s932 (.CLK(clknet_4_4_0_clk),
    .D(net359),
    .Q(net708),
    .Q_N(net707));
 sky130_fd_sc_hd__dfxbp_2 s933 (.CLK(clknet_4_1_0_clk),
    .D(net360),
    .Q(net855),
    .Q_N(net709));
 sky130_fd_sc_hd__dfxtp_1 s934 (.CLK(clknet_4_6_0_clk),
    .D(net361),
    .Q(net710));
 sky130_fd_sc_hd__dfxtp_2 s935 (.CLK(clknet_4_4_0_clk),
    .D(net365),
    .Q(net711));
 sky130_fd_sc_hd__dfxtp_2 s936 (.CLK(clknet_4_3_0_clk),
    .D(net369),
    .Q(net712));
 sky130_fd_sc_hd__dlclkp_1 s937 (.CLK(clknet_4_4_0_clk),
    .GATE(net371),
    .GCLK(net713));
 sky130_fd_sc_hd__dlclkp_2 s938 (.CLK(clknet_4_4_0_clk),
    .GATE(net373),
    .GCLK(net714));
 sky130_fd_sc_hd__dlclkp_4 s939 (.CLK(clknet_4_4_0_clk),
    .GATE(net374),
    .GCLK(net715));
 sky130_fd_sc_hd__dlxbn_1 s940 (.D(net376),
    .GATE_N(clknet_4_6_0_clk),
    .Q(net717),
    .Q_N(net716));
 sky130_fd_sc_hd__dlxbn_1 s941 (.D(net378),
    .GATE_N(clknet_4_6_0_clk),
    .Q(net719),
    .Q_N(net718));
 sky130_fd_sc_hd__dlxbp_1 s942 (.D(net379),
    .GATE(clknet_4_6_0_clk),
    .Q(net721),
    .Q_N(net720));
 sky130_fd_sc_hd__dlxtn_1 s943 (.D(net384),
    .GATE_N(clknet_4_3_0_clk),
    .Q(net722));
 sky130_fd_sc_hd__dlxtn_1 s944 (.D(net387),
    .GATE_N(clknet_4_6_0_clk),
    .Q(net875));
 sky130_fd_sc_hd__dlxtn_2 s945 (.D(net392),
    .GATE_N(clknet_4_6_0_clk),
    .Q(net723));
 sky130_fd_sc_hd__dlxtp_1 s946 (.D(net393),
    .GATE(clknet_4_6_0_clk),
    .Q(net724));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s947 (.D(net395),
    .SLEEP_B(clknet_4_6_0_clk),
    .Q(net852));
 sky130_fd_sc_hd__dfxbp_1 s948 (.CLK(clknet_4_6_0_clk),
    .D(net397),
    .Q(net726),
    .Q_N(net725));
 sky130_fd_sc_hd__dfxbp_1 s949 (.CLK(clknet_4_7_0_clk),
    .D(net399),
    .Q(net728),
    .Q_N(net727));
 sky130_fd_sc_hd__dfxtp_1 s950 (.CLK(clknet_4_6_0_clk),
    .D(net400),
    .Q(net729));
 sky130_fd_sc_hd__dfxtp_1 s951 (.CLK(clknet_4_12_0_clk),
    .D(net415),
    .Q(net730));
 sky130_fd_sc_hd__dfxtp_1 s952 (.CLK(clknet_4_14_0_clk),
    .D(net424),
    .Q(net731));
 sky130_fd_sc_hd__dlclkp_1 s953 (.CLK(clknet_4_15_0_clk),
    .GATE(net426),
    .GCLK(net732));
 sky130_fd_sc_hd__dlclkp_2 s954 (.CLK(clknet_4_14_0_clk),
    .GATE(net427),
    .GCLK(net733));
 sky130_fd_sc_hd__dlclkp_4 s955 (.CLK(clknet_4_15_0_clk),
    .GATE(net435),
    .GCLK(net734));
 sky130_fd_sc_hd__dlxbn_1 s956 (.D(net441),
    .GATE_N(clknet_4_15_0_clk),
    .Q(net736),
    .Q_N(net735));
 sky130_fd_sc_hd__dlxbn_1 s957 (.D(net445),
    .GATE_N(clknet_4_5_0_clk),
    .Q(net738),
    .Q_N(net737));
 sky130_fd_sc_hd__dlxbp_1 s958 (.D(net452),
    .GATE(clknet_4_5_0_clk),
    .Q(net740),
    .Q_N(net739));
 sky130_fd_sc_hd__dlxtn_1 s959 (.D(net461),
    .GATE_N(clknet_4_5_0_clk),
    .Q(net741));
 sky130_fd_sc_hd__dlxtn_1 s960 (.D(net462),
    .GATE_N(clknet_4_5_0_clk),
    .Q(net742));
 sky130_fd_sc_hd__dlxtn_2 s961 (.D(net471),
    .GATE_N(clknet_4_5_0_clk),
    .Q(net743));
 sky130_fd_sc_hd__dlxtp_1 s962 (.D(net473),
    .GATE(clknet_4_7_0_clk),
    .Q(net744));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s963 (.D(net475),
    .SLEEP_B(clknet_4_5_0_clk),
    .Q(net745));
 sky130_fd_sc_hd__dfxbp_2 s964 (.CLK(clknet_4_5_0_clk),
    .D(net479),
    .Q(net747),
    .Q_N(net746));
 sky130_fd_sc_hd__dfxbp_1 s965 (.CLK(clknet_4_7_0_clk),
    .D(net490),
    .Q(net749),
    .Q_N(net748));
 sky130_fd_sc_hd__dfxtp_1 s966 (.CLK(clknet_4_7_0_clk),
    .D(net491),
    .Q(net750));
 sky130_fd_sc_hd__dfxtp_1 s967 (.CLK(clknet_4_7_0_clk),
    .D(net501),
    .Q(net860));
 sky130_fd_sc_hd__dfxtp_1 s968 (.CLK(clknet_4_7_0_clk),
    .D(net510),
    .Q(net751));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Right_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Right_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Right_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Right_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Right_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Right_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Right_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Right_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Right_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Right_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Right_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Right_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Right_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Right_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Right_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Right_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Right_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Right_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Right_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Right_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Right_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_161 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_162 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_163 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_164 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_165 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_166 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_167 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_168 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_169 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_170 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_171 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_172 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_173 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_174 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_175 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_176 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_177 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_178 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_179 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_180 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_181 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_182 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Left_183 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Left_184 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Left_185 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Left_186 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Left_187 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Left_188 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Left_189 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Left_190 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Left_191 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Left_192 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Left_193 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Left_194 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Left_195 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Left_196 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Left_197 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Left_198 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Left_199 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Left_200 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Left_201 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Left_202 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Left_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1347 ();
 sky130_fd_sc_hd__clkbuf_4 input1 (.A(in0),
    .X(net194));
 sky130_fd_sc_hd__clkbuf_2 input2 (.A(in1),
    .X(net752));
 sky130_fd_sc_hd__buf_2 input3 (.A(in10),
    .X(net753));
 sky130_fd_sc_hd__buf_2 input4 (.A(in11),
    .X(net754));
 sky130_fd_sc_hd__clkbuf_2 input5 (.A(in12),
    .X(net755));
 sky130_fd_sc_hd__clkbuf_4 input6 (.A(in13),
    .X(net756));
 sky130_fd_sc_hd__buf_2 input7 (.A(in14),
    .X(net757));
 sky130_fd_sc_hd__clkbuf_2 input8 (.A(in15),
    .X(net758));
 sky130_fd_sc_hd__buf_1 input9 (.A(in16),
    .X(net759));
 sky130_fd_sc_hd__buf_2 input10 (.A(in17),
    .X(net760));
 sky130_fd_sc_hd__clkbuf_2 input11 (.A(in18),
    .X(net761));
 sky130_fd_sc_hd__clkbuf_2 input12 (.A(in19),
    .X(net762));
 sky130_fd_sc_hd__buf_2 input13 (.A(in2),
    .X(net763));
 sky130_fd_sc_hd__buf_2 input14 (.A(in20),
    .X(net764));
 sky130_fd_sc_hd__clkbuf_4 input15 (.A(in21),
    .X(net765));
 sky130_fd_sc_hd__buf_2 input16 (.A(in22),
    .X(net766));
 sky130_fd_sc_hd__clkbuf_2 input17 (.A(in23),
    .X(net767));
 sky130_fd_sc_hd__clkbuf_2 input18 (.A(in24),
    .X(net768));
 sky130_fd_sc_hd__clkbuf_2 input19 (.A(in25),
    .X(net769));
 sky130_fd_sc_hd__clkbuf_2 input20 (.A(in26),
    .X(net770));
 sky130_fd_sc_hd__clkbuf_2 input21 (.A(in27),
    .X(net771));
 sky130_fd_sc_hd__buf_2 input22 (.A(in28),
    .X(net772));
 sky130_fd_sc_hd__clkbuf_4 input23 (.A(in29),
    .X(net773));
 sky130_fd_sc_hd__buf_12 input24 (.A(in3),
    .X(net774));
 sky130_fd_sc_hd__clkbuf_2 input25 (.A(in30),
    .X(net775));
 sky130_fd_sc_hd__buf_4 input26 (.A(in31),
    .X(net776));
 sky130_fd_sc_hd__clkbuf_2 input27 (.A(in32),
    .X(net777));
 sky130_fd_sc_hd__clkbuf_4 input28 (.A(in33),
    .X(net778));
 sky130_fd_sc_hd__dlymetal6s2s_1 input29 (.A(in34),
    .X(net779));
 sky130_fd_sc_hd__clkbuf_2 input30 (.A(in35),
    .X(net780));
 sky130_fd_sc_hd__buf_2 input31 (.A(in36),
    .X(net781));
 sky130_fd_sc_hd__buf_2 input32 (.A(in37),
    .X(net782));
 sky130_fd_sc_hd__clkbuf_2 input33 (.A(in38),
    .X(net783));
 sky130_fd_sc_hd__buf_2 input34 (.A(in39),
    .X(net784));
 sky130_fd_sc_hd__clkbuf_4 input35 (.A(in4),
    .X(net785));
 sky130_fd_sc_hd__buf_6 input36 (.A(in40),
    .X(net786));
 sky130_fd_sc_hd__buf_4 input37 (.A(in41),
    .X(net787));
 sky130_fd_sc_hd__buf_2 input38 (.A(in42),
    .X(net788));
 sky130_fd_sc_hd__buf_4 input39 (.A(in43),
    .X(net789));
 sky130_fd_sc_hd__clkbuf_2 input40 (.A(in44),
    .X(net790));
 sky130_fd_sc_hd__buf_4 input41 (.A(in45),
    .X(net791));
 sky130_fd_sc_hd__clkbuf_4 input42 (.A(in46),
    .X(net792));
 sky130_fd_sc_hd__buf_1 input43 (.A(in47),
    .X(net793));
 sky130_fd_sc_hd__clkbuf_4 input44 (.A(in48),
    .X(net794));
 sky130_fd_sc_hd__dlymetal6s2s_1 input45 (.A(in49),
    .X(net795));
 sky130_fd_sc_hd__buf_2 input46 (.A(in5),
    .X(net796));
 sky130_fd_sc_hd__dlymetal6s2s_1 input47 (.A(in50),
    .X(net797));
 sky130_fd_sc_hd__buf_2 input48 (.A(in51),
    .X(net798));
 sky130_fd_sc_hd__clkbuf_4 input49 (.A(in52),
    .X(net799));
 sky130_fd_sc_hd__clkbuf_4 input50 (.A(in53),
    .X(net800));
 sky130_fd_sc_hd__clkbuf_2 input51 (.A(in54),
    .X(net801));
 sky130_fd_sc_hd__clkbuf_2 input52 (.A(in55),
    .X(net802));
 sky130_fd_sc_hd__buf_4 input53 (.A(in56),
    .X(net803));
 sky130_fd_sc_hd__buf_2 input54 (.A(in57),
    .X(net804));
 sky130_fd_sc_hd__buf_4 input55 (.A(in58),
    .X(net805));
 sky130_fd_sc_hd__buf_1 input56 (.A(in59),
    .X(net806));
 sky130_fd_sc_hd__clkbuf_2 input57 (.A(in6),
    .X(net807));
 sky130_fd_sc_hd__buf_2 input58 (.A(in60),
    .X(net808));
 sky130_fd_sc_hd__buf_2 input59 (.A(in61),
    .X(net809));
 sky130_fd_sc_hd__buf_4 input60 (.A(in62),
    .X(net810));
 sky130_fd_sc_hd__clkbuf_1 input61 (.A(in63),
    .X(net811));
 sky130_fd_sc_hd__clkbuf_2 input62 (.A(in64),
    .X(net812));
 sky130_fd_sc_hd__dlymetal6s2s_1 input63 (.A(in65),
    .X(net813));
 sky130_fd_sc_hd__dlymetal6s2s_1 input64 (.A(in66),
    .X(net814));
 sky130_fd_sc_hd__clkbuf_1 input65 (.A(in67),
    .X(net815));
 sky130_fd_sc_hd__clkbuf_1 input66 (.A(in68),
    .X(net816));
 sky130_fd_sc_hd__clkbuf_4 input67 (.A(in69),
    .X(net817));
 sky130_fd_sc_hd__clkbuf_2 input68 (.A(in7),
    .X(net818));
 sky130_fd_sc_hd__clkbuf_4 input69 (.A(in70),
    .X(net819));
 sky130_fd_sc_hd__buf_1 input70 (.A(in71),
    .X(net820));
 sky130_fd_sc_hd__buf_2 input71 (.A(in72),
    .X(net821));
 sky130_fd_sc_hd__dlymetal6s2s_1 input72 (.A(in73),
    .X(net822));
 sky130_fd_sc_hd__clkbuf_4 input73 (.A(in74),
    .X(net823));
 sky130_fd_sc_hd__clkbuf_4 input74 (.A(in75),
    .X(net824));
 sky130_fd_sc_hd__clkbuf_2 input75 (.A(in76),
    .X(net825));
 sky130_fd_sc_hd__buf_1 input76 (.A(in77),
    .X(net826));
 sky130_fd_sc_hd__clkbuf_1 input77 (.A(in78),
    .X(net827));
 sky130_fd_sc_hd__buf_1 input78 (.A(in79),
    .X(net828));
 sky130_fd_sc_hd__clkbuf_2 input79 (.A(in8),
    .X(net829));
 sky130_fd_sc_hd__buf_1 input80 (.A(in80),
    .X(net830));
 sky130_fd_sc_hd__dlymetal6s2s_1 input81 (.A(in81),
    .X(net831));
 sky130_fd_sc_hd__clkbuf_4 input82 (.A(in82),
    .X(net832));
 sky130_fd_sc_hd__buf_2 input83 (.A(in83),
    .X(net833));
 sky130_fd_sc_hd__buf_1 input84 (.A(in84),
    .X(net834));
 sky130_fd_sc_hd__clkbuf_1 input85 (.A(in85),
    .X(net835));
 sky130_fd_sc_hd__buf_1 input86 (.A(in86),
    .X(net836));
 sky130_fd_sc_hd__buf_1 input87 (.A(in87),
    .X(net837));
 sky130_fd_sc_hd__buf_1 input88 (.A(in88),
    .X(net838));
 sky130_fd_sc_hd__buf_1 input89 (.A(in89),
    .X(net839));
 sky130_fd_sc_hd__buf_4 input90 (.A(in9),
    .X(net840));
 sky130_fd_sc_hd__buf_1 input91 (.A(in90),
    .X(net841));
 sky130_fd_sc_hd__clkbuf_4 input92 (.A(in91),
    .X(net842));
 sky130_fd_sc_hd__clkbuf_4 input93 (.A(in92),
    .X(net843));
 sky130_fd_sc_hd__buf_4 input94 (.A(in93),
    .X(net844));
 sky130_fd_sc_hd__buf_2 input95 (.A(in94),
    .X(net845));
 sky130_fd_sc_hd__buf_1 input96 (.A(in95),
    .X(net846));
 sky130_fd_sc_hd__clkbuf_1 input97 (.A(in96),
    .X(net847));
 sky130_fd_sc_hd__buf_2 input98 (.A(in97),
    .X(net848));
 sky130_fd_sc_hd__clkbuf_2 input99 (.A(in98),
    .X(net849));
 sky130_fd_sc_hd__buf_1 input100 (.A(in99),
    .X(net850));
 sky130_fd_sc_hd__buf_2 output101 (.A(net1118),
    .X(out0));
 sky130_fd_sc_hd__buf_2 output102 (.A(net852),
    .X(out10));
 sky130_fd_sc_hd__clkbuf_4 output103 (.A(net853),
    .X(out11));
 sky130_fd_sc_hd__buf_2 output104 (.A(net854),
    .X(out12));
 sky130_fd_sc_hd__buf_2 output105 (.A(net855),
    .X(out13));
 sky130_fd_sc_hd__buf_2 output106 (.A(net856),
    .X(out14));
 sky130_fd_sc_hd__buf_2 output107 (.A(net967),
    .X(out15));
 sky130_fd_sc_hd__clkbuf_4 output108 (.A(net858),
    .X(out18));
 sky130_fd_sc_hd__clkbuf_4 output109 (.A(net859),
    .X(out19));
 sky130_fd_sc_hd__buf_2 output110 (.A(net860),
    .X(out2));
 sky130_fd_sc_hd__clkbuf_4 output111 (.A(net861),
    .X(out20));
 sky130_fd_sc_hd__buf_2 output112 (.A(net862),
    .X(out22));
 sky130_fd_sc_hd__buf_2 output113 (.A(net863),
    .X(out23));
 sky130_fd_sc_hd__clkbuf_4 output114 (.A(net864),
    .X(out24));
 sky130_fd_sc_hd__buf_2 output115 (.A(net865),
    .X(out25));
 sky130_fd_sc_hd__buf_2 output116 (.A(net962),
    .X(out26));
 sky130_fd_sc_hd__clkbuf_4 output117 (.A(net867),
    .X(out27));
 sky130_fd_sc_hd__clkbuf_1 output118 (.A(clknet_1_1__leaf_net868),
    .X(out28));
 sky130_fd_sc_hd__buf_2 output119 (.A(net869),
    .X(out29));
 sky130_fd_sc_hd__clkbuf_4 output120 (.A(net870),
    .X(out30));
 sky130_fd_sc_hd__clkbuf_4 output121 (.A(net871),
    .X(out31));
 sky130_fd_sc_hd__buf_2 output122 (.A(net872),
    .X(out32));
 sky130_fd_sc_hd__clkbuf_4 output123 (.A(net873),
    .X(out33));
 sky130_fd_sc_hd__buf_2 output124 (.A(net874),
    .X(out34));
 sky130_fd_sc_hd__buf_2 output125 (.A(net875),
    .X(out35));
 sky130_fd_sc_hd__clkbuf_4 output126 (.A(net876),
    .X(out36));
 sky130_fd_sc_hd__clkbuf_1 output127 (.A(clknet_1_1__leaf_net877),
    .X(out37));
 sky130_fd_sc_hd__clkbuf_4 output128 (.A(net878),
    .X(out38));
 sky130_fd_sc_hd__clkbuf_4 output129 (.A(net1044),
    .X(out39));
 sky130_fd_sc_hd__buf_2 output130 (.A(net880),
    .X(out42));
 sky130_fd_sc_hd__clkbuf_4 output131 (.A(net881),
    .X(out43));
 sky130_fd_sc_hd__clkbuf_1 output132 (.A(clknet_1_1__leaf_net882),
    .X(out45));
 sky130_fd_sc_hd__clkbuf_4 output133 (.A(net883),
    .X(out47));
 sky130_fd_sc_hd__buf_2 output134 (.A(net884),
    .X(out48));
 sky130_fd_sc_hd__buf_2 output135 (.A(net885),
    .X(out49));
 sky130_fd_sc_hd__buf_2 output136 (.A(net886),
    .X(out50));
 sky130_fd_sc_hd__clkbuf_1 output137 (.A(clknet_1_1__leaf_net887),
    .X(out52));
 sky130_fd_sc_hd__buf_2 output138 (.A(net888),
    .X(out53));
 sky130_fd_sc_hd__clkbuf_4 output139 (.A(net889),
    .X(out54));
 sky130_fd_sc_hd__clkbuf_4 output140 (.A(net890),
    .X(out55));
 sky130_fd_sc_hd__buf_2 output141 (.A(net891),
    .X(out57));
 sky130_fd_sc_hd__clkbuf_4 output142 (.A(net892),
    .X(out58));
 sky130_fd_sc_hd__buf_2 output143 (.A(net893),
    .X(out59));
 sky130_fd_sc_hd__buf_2 output144 (.A(net894),
    .X(out6));
 sky130_fd_sc_hd__clkbuf_4 output145 (.A(net895),
    .X(out60));
 sky130_fd_sc_hd__buf_2 output146 (.A(net896),
    .X(out62));
 sky130_fd_sc_hd__clkbuf_4 output147 (.A(net897),
    .X(out63));
 sky130_fd_sc_hd__buf_2 output148 (.A(net1114),
    .X(out64));
 sky130_fd_sc_hd__clkbuf_4 output149 (.A(net899),
    .X(out66));
 sky130_fd_sc_hd__clkbuf_4 output150 (.A(net900),
    .X(out67));
 sky130_fd_sc_hd__clkbuf_4 output151 (.A(net901),
    .X(out68));
 sky130_fd_sc_hd__clkbuf_4 output152 (.A(net902),
    .X(out69));
 sky130_fd_sc_hd__clkbuf_4 output153 (.A(net903),
    .X(out7));
 sky130_fd_sc_hd__clkbuf_4 output154 (.A(net904),
    .X(out70));
 sky130_fd_sc_hd__clkbuf_4 output155 (.A(net905),
    .X(out71));
 sky130_fd_sc_hd__clkbuf_4 output156 (.A(net906),
    .X(out73));
 sky130_fd_sc_hd__clkbuf_1 output157 (.A(clknet_1_1__leaf_net907),
    .X(out74));
 sky130_fd_sc_hd__clkbuf_4 output158 (.A(net908),
    .X(out75));
 sky130_fd_sc_hd__clkbuf_4 output159 (.A(net909),
    .X(out76));
 sky130_fd_sc_hd__clkbuf_4 output160 (.A(net910),
    .X(out77));
 sky130_fd_sc_hd__buf_2 output161 (.A(net911),
    .X(out78));
 sky130_fd_sc_hd__clkbuf_1 output162 (.A(clknet_1_1__leaf_net912),
    .X(out79));
 sky130_fd_sc_hd__clkbuf_1 output163 (.A(clknet_1_1__leaf_net913),
    .X(out8));
 sky130_fd_sc_hd__buf_2 output164 (.A(net914),
    .X(out80));
 sky130_fd_sc_hd__buf_2 output165 (.A(net915),
    .X(out81));
 sky130_fd_sc_hd__clkbuf_4 output166 (.A(net916),
    .X(out82));
 sky130_fd_sc_hd__buf_2 output167 (.A(net917),
    .X(out84));
 sky130_fd_sc_hd__clkbuf_4 output168 (.A(net918),
    .X(out85));
 sky130_fd_sc_hd__clkbuf_4 output169 (.A(net919),
    .X(out86));
 sky130_fd_sc_hd__clkbuf_4 output170 (.A(net920),
    .X(out87));
 sky130_fd_sc_hd__clkbuf_1 output171 (.A(clknet_1_1__leaf_net921),
    .X(out88));
 sky130_fd_sc_hd__clkbuf_4 output172 (.A(net1106),
    .X(out89));
 sky130_fd_sc_hd__buf_2 output173 (.A(net923),
    .X(out9));
 sky130_fd_sc_hd__buf_2 output174 (.A(net924),
    .X(out90));
 sky130_fd_sc_hd__clkbuf_4 output175 (.A(net925),
    .X(out91));
 sky130_fd_sc_hd__clkbuf_4 output176 (.A(net926),
    .X(out93));
 sky130_fd_sc_hd__clkbuf_4 output177 (.A(net927),
    .X(out94));
 sky130_fd_sc_hd__buf_2 output178 (.A(net928),
    .X(out95));
 sky130_fd_sc_hd__clkbuf_4 output179 (.A(net929),
    .X(out96));
 sky130_fd_sc_hd__clkbuf_4 output180 (.A(net930),
    .X(out97));
 sky130_fd_sc_hd__clkbuf_1 output181 (.A(net931),
    .X(out99));
 sky130_fd_sc_hd__clkbuf_4 fanout182 (.A(net257),
    .X(net932));
 sky130_fd_sc_hd__clkbuf_4 fanout183 (.A(net92),
    .X(net933));
 sky130_fd_sc_hd__buf_4 fanout184 (.A(net137),
    .X(net934));
 sky130_fd_sc_hd__buf_12 fanout185 (.A(net49),
    .X(net935));
 sky130_fd_sc_hd__buf_8 fanout186 (.A(net133),
    .X(net936));
 sky130_fd_sc_hd__buf_6 fanout187 (.A(net939),
    .X(net937));
 sky130_fd_sc_hd__buf_2 fanout188 (.A(net939),
    .X(net938));
 sky130_fd_sc_hd__buf_4 fanout189 (.A(net132),
    .X(net939));
 sky130_fd_sc_hd__clkbuf_4 fanout190 (.A(net861),
    .X(net940));
 sky130_fd_sc_hd__clkbuf_4 fanout191 (.A(net222),
    .X(net941));
 sky130_fd_sc_hd__buf_6 fanout192 (.A(net126),
    .X(net942));
 sky130_fd_sc_hd__buf_12 fanout193 (.A(net43),
    .X(net943));
 sky130_fd_sc_hd__buf_8 fanout194 (.A(net945),
    .X(net944));
 sky130_fd_sc_hd__buf_8 fanout195 (.A(net946),
    .X(net945));
 sky130_fd_sc_hd__buf_12 fanout196 (.A(net947),
    .X(net946));
 sky130_fd_sc_hd__buf_12 fanout197 (.A(net123),
    .X(net947));
 sky130_fd_sc_hd__buf_4 fanout198 (.A(net41),
    .X(net948));
 sky130_fd_sc_hd__clkbuf_4 fanout199 (.A(net950),
    .X(net949));
 sky130_fd_sc_hd__clkbuf_2 fanout200 (.A(net951),
    .X(net950));
 sky130_fd_sc_hd__buf_2 fanout201 (.A(net952),
    .X(net951));
 sky130_fd_sc_hd__clkbuf_4 fanout202 (.A(net118),
    .X(net952));
 sky130_fd_sc_hd__buf_8 fanout203 (.A(net40),
    .X(net953));
 sky130_fd_sc_hd__buf_4 fanout204 (.A(net39),
    .X(net954));
 sky130_fd_sc_hd__buf_8 fanout205 (.A(net32),
    .X(net955));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout206 (.A(net1059),
    .X(net956));
 sky130_fd_sc_hd__buf_8 fanout207 (.A(net898),
    .X(net957));
 sky130_fd_sc_hd__buf_12 fanout208 (.A(net31),
    .X(net958));
 sky130_fd_sc_hd__clkbuf_2 fanout209 (.A(net1064),
    .X(net959));
 sky130_fd_sc_hd__buf_8 fanout210 (.A(net961),
    .X(net960));
 sky130_fd_sc_hd__buf_8 fanout211 (.A(net37),
    .X(net961));
 sky130_fd_sc_hd__clkbuf_8 fanout212 (.A(net866),
    .X(net962));
 sky130_fd_sc_hd__buf_12 fanout213 (.A(net30),
    .X(net963));
 sky130_fd_sc_hd__buf_8 fanout214 (.A(net35),
    .X(net964));
 sky130_fd_sc_hd__buf_4 fanout215 (.A(net29),
    .X(net965));
 sky130_fd_sc_hd__buf_12 fanout216 (.A(net27),
    .X(net966));
 sky130_fd_sc_hd__buf_8 fanout217 (.A(net969),
    .X(net967));
 sky130_fd_sc_hd__buf_2 fanout218 (.A(net969),
    .X(net968));
 sky130_fd_sc_hd__buf_8 fanout219 (.A(net857),
    .X(net969));
 sky130_fd_sc_hd__buf_8 fanout220 (.A(net28),
    .X(net970));
 sky130_fd_sc_hd__buf_8 fanout221 (.A(net23),
    .X(net971));
 sky130_fd_sc_hd__buf_12 fanout222 (.A(net973),
    .X(net972));
 sky130_fd_sc_hd__buf_8 fanout223 (.A(net974),
    .X(net973));
 sky130_fd_sc_hd__buf_12 fanout224 (.A(net21),
    .X(net974));
 sky130_fd_sc_hd__buf_8 fanout225 (.A(net20),
    .X(net975));
 sky130_fd_sc_hd__clkbuf_4 fanout226 (.A(net20),
    .X(net976));
 sky130_fd_sc_hd__buf_12 fanout227 (.A(net978),
    .X(net977));
 sky130_fd_sc_hd__buf_12 fanout228 (.A(net851),
    .X(net978));
 sky130_fd_sc_hd__buf_8 fanout229 (.A(net19),
    .X(net979));
 sky130_fd_sc_hd__buf_6 fanout230 (.A(net16),
    .X(net980));
 sky130_fd_sc_hd__buf_2 max_cap231 (.A(net685),
    .X(net981));
 sky130_fd_sc_hd__clkbuf_4 fanout232 (.A(net671),
    .X(net982));
 sky130_fd_sc_hd__clkbuf_4 fanout233 (.A(net664),
    .X(net983));
 sky130_fd_sc_hd__buf_2 fanout234 (.A(net664),
    .X(net984));
 sky130_fd_sc_hd__buf_4 fanout235 (.A(net655),
    .X(net985));
 sky130_fd_sc_hd__clkbuf_4 fanout236 (.A(net987),
    .X(net986));
 sky130_fd_sc_hd__buf_2 fanout237 (.A(net988),
    .X(net987));
 sky130_fd_sc_hd__clkbuf_4 fanout238 (.A(net653),
    .X(net988));
 sky130_fd_sc_hd__clkbuf_4 max_cap239 (.A(net608),
    .X(net989));
 sky130_fd_sc_hd__buf_4 max_cap240 (.A(net566),
    .X(net990));
 sky130_fd_sc_hd__buf_12 fanout241 (.A(net922),
    .X(net991));
 sky130_fd_sc_hd__buf_4 fanout242 (.A(net840),
    .X(net992));
 sky130_fd_sc_hd__clkbuf_4 fanout243 (.A(net759),
    .X(net993));
 sky130_fd_sc_hd__buf_12 fanout244 (.A(net758),
    .X(net994));
 sky130_fd_sc_hd__clkbuf_2 fanout245 (.A(net758),
    .X(net995));
 sky130_fd_sc_hd__buf_4 fanout246 (.A(net829),
    .X(net996));
 sky130_fd_sc_hd__clkbuf_2 fanout247 (.A(net829),
    .X(net997));
 sky130_fd_sc_hd__buf_6 fanout248 (.A(net757),
    .X(net998));
 sky130_fd_sc_hd__buf_4 fanout249 (.A(net818),
    .X(net999));
 sky130_fd_sc_hd__buf_2 fanout250 (.A(net818),
    .X(net1000));
 sky130_fd_sc_hd__buf_4 fanout251 (.A(net807),
    .X(net1001));
 sky130_fd_sc_hd__buf_2 fanout252 (.A(net807),
    .X(net1002));
 sky130_fd_sc_hd__buf_4 fanout253 (.A(net755),
    .X(net1003));
 sky130_fd_sc_hd__buf_2 fanout254 (.A(net755),
    .X(net1004));
 sky130_fd_sc_hd__buf_4 fanout255 (.A(net796),
    .X(net1005));
 sky130_fd_sc_hd__buf_4 fanout256 (.A(net754),
    .X(net1006));
 sky130_fd_sc_hd__buf_12 fanout257 (.A(net785),
    .X(net1007));
 sky130_fd_sc_hd__buf_4 fanout258 (.A(net782),
    .X(net1008));
 sky130_fd_sc_hd__buf_4 fanout259 (.A(net775),
    .X(net1009));
 sky130_fd_sc_hd__buf_12 fanout260 (.A(net1011),
    .X(net1010));
 sky130_fd_sc_hd__buf_12 fanout261 (.A(net1013),
    .X(net1011));
 sky130_fd_sc_hd__clkbuf_4 fanout262 (.A(net1013),
    .X(net1012));
 sky130_fd_sc_hd__buf_8 fanout263 (.A(net774),
    .X(net1013));
 sky130_fd_sc_hd__clkbuf_4 fanout264 (.A(net1015),
    .X(net1014));
 sky130_fd_sc_hd__buf_2 fanout265 (.A(net774),
    .X(net1015));
 sky130_fd_sc_hd__buf_4 fanout266 (.A(net752),
    .X(net1016));
 sky130_fd_sc_hd__clkbuf_8 fanout267 (.A(net769),
    .X(net1017));
 sky130_fd_sc_hd__buf_2 fanout268 (.A(net769),
    .X(net1018));
 sky130_fd_sc_hd__clkbuf_4 fanout269 (.A(net768),
    .X(net1019));
 sky130_fd_sc_hd__buf_4 fanout270 (.A(net765),
    .X(net1020));
 sky130_fd_sc_hd__buf_4 fanout271 (.A(net764),
    .X(net1021));
 sky130_fd_sc_hd__buf_4 fanout272 (.A(net763),
    .X(net1022));
 sky130_fd_sc_hd__buf_4 fanout273 (.A(net762),
    .X(net1023));
 sky130_fd_sc_hd__buf_6 fanout274 (.A(net761),
    .X(net1024));
 sky130_fd_sc_hd__clkbuf_8 fanout275 (.A(net760),
    .X(net1025));
 sky130_fd_sc_hd__buf_4 fanout276 (.A(net194),
    .X(net1026));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net734 (.A(net734),
    .X(clknet_0_net734));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net734 (.A(clknet_0_net734),
    .X(clknet_1_0__leaf_net734));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net734 (.A(clknet_0_net734),
    .X(clknet_1_1__leaf_net734));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net733 (.A(net733),
    .X(clknet_0_net733));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net733 (.A(clknet_0_net733),
    .X(clknet_1_0__leaf_net733));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net733 (.A(clknet_0_net733),
    .X(clknet_1_1__leaf_net733));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net732 (.A(net732),
    .X(clknet_0_net732));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net732 (.A(clknet_0_net732),
    .X(clknet_1_0__leaf_net732));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net732 (.A(clknet_0_net732),
    .X(clknet_1_1__leaf_net732));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net429 (.A(net429),
    .X(clknet_0_net429));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net429 (.A(clknet_0_net429),
    .X(clknet_1_0__leaf_net429));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net429 (.A(clknet_0_net429),
    .X(clknet_1_1__leaf_net429));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net715 (.A(net715),
    .X(clknet_0_net715));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net715 (.A(clknet_0_net715),
    .X(clknet_1_0__leaf_net715));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net715 (.A(clknet_0_net715),
    .X(clknet_1_1__leaf_net715));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net380 (.A(net380),
    .X(clknet_0_net380));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net380 (.A(clknet_0_net380),
    .X(clknet_1_0__leaf_net380));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net380 (.A(clknet_0_net380),
    .X(clknet_1_1__leaf_net380));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net377 (.A(net377),
    .X(clknet_0_net377));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net377 (.A(clknet_0_net377),
    .X(clknet_1_0__leaf_net377));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net377 (.A(clknet_0_net377),
    .X(clknet_1_1__leaf_net377));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net375 (.A(net375),
    .X(clknet_0_net375));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net375 (.A(clknet_0_net375),
    .X(clknet_1_0__leaf_net375));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net375 (.A(clknet_0_net375),
    .X(clknet_1_1__leaf_net375));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net714 (.A(net714),
    .X(clknet_0_net714));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net714 (.A(clknet_0_net714),
    .X(clknet_1_0__leaf_net714));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net714 (.A(clknet_0_net714),
    .X(clknet_1_1__leaf_net714));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net407 (.A(net407),
    .X(clknet_0_net407));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net407 (.A(clknet_0_net407),
    .X(clknet_1_0__leaf_net407));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net407 (.A(clknet_0_net407),
    .X(clknet_1_1__leaf_net407));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net713 (.A(net713),
    .X(clknet_0_net713));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net713 (.A(clknet_0_net713),
    .X(clknet_1_0__leaf_net713));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net713 (.A(clknet_0_net713),
    .X(clknet_1_1__leaf_net713));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net372 (.A(net372),
    .X(clknet_0_net372));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net372 (.A(clknet_0_net372),
    .X(clknet_1_0__leaf_net372));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net372 (.A(clknet_0_net372),
    .X(clknet_1_1__leaf_net372));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net695 (.A(net695),
    .X(clknet_0_net695));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net695 (.A(clknet_0_net695),
    .X(clknet_1_0__leaf_net695));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net695 (.A(clknet_0_net695),
    .X(clknet_1_1__leaf_net695));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net310 (.A(net310),
    .X(clknet_0_net310));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net310 (.A(clknet_0_net310),
    .X(clknet_1_0__leaf_net310));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net310 (.A(clknet_0_net310),
    .X(clknet_1_1__leaf_net310));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net527 (.A(net527),
    .X(clknet_0_net527));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net527 (.A(clknet_0_net527),
    .X(clknet_1_0__leaf_net527));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net527 (.A(clknet_0_net527),
    .X(clknet_1_1__leaf_net527));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net694 (.A(net694),
    .X(clknet_0_net694));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net694 (.A(clknet_0_net694),
    .X(clknet_1_0__leaf_net694));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net694 (.A(clknet_0_net694),
    .X(clknet_1_1__leaf_net694));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net868 (.A(net868),
    .X(clknet_0_net868));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net868 (.A(clknet_0_net868),
    .X(clknet_1_0__leaf_net868));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net868 (.A(clknet_0_net868),
    .X(clknet_1_1__leaf_net868));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net302 (.A(net302),
    .X(clknet_0_net302));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net302 (.A(clknet_0_net302),
    .X(clknet_1_0__leaf_net302));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net302 (.A(clknet_0_net302),
    .X(clknet_1_1__leaf_net302));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net882 (.A(net882),
    .X(clknet_0_net882));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net882 (.A(clknet_0_net882),
    .X(clknet_1_0__leaf_net882));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net882 (.A(clknet_0_net882),
    .X(clknet_1_1__leaf_net882));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net693 (.A(net693),
    .X(clknet_0_net693));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net693 (.A(clknet_0_net693),
    .X(clknet_1_0__leaf_net693));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net693 (.A(clknet_0_net693),
    .X(clknet_1_1__leaf_net693));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net675 (.A(net675),
    .X(clknet_0_net675));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net675 (.A(clknet_0_net675),
    .X(clknet_1_0__leaf_net675));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net675 (.A(clknet_0_net675),
    .X(clknet_1_1__leaf_net675));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net913 (.A(net913),
    .X(clknet_0_net913));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net913 (.A(clknet_0_net913),
    .X(clknet_1_0__leaf_net913));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net913 (.A(clknet_0_net913),
    .X(clknet_1_1__leaf_net913));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net521 (.A(net521),
    .X(clknet_0_net521));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net521 (.A(clknet_0_net521),
    .X(clknet_1_0__leaf_net521));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net521 (.A(clknet_0_net521),
    .X(clknet_1_1__leaf_net521));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net495 (.A(net495),
    .X(clknet_0_net495));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net495 (.A(clknet_0_net495),
    .X(clknet_1_0__leaf_net495));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net495 (.A(clknet_0_net495),
    .X(clknet_1_1__leaf_net495));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net451 (.A(net451),
    .X(clknet_0_net451));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net451 (.A(clknet_0_net451),
    .X(clknet_1_0__leaf_net451));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net451 (.A(clknet_0_net451),
    .X(clknet_1_1__leaf_net451));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net469 (.A(net469),
    .X(clknet_0_net469));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net469 (.A(clknet_0_net469),
    .X(clknet_1_0__leaf_net469));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net469 (.A(clknet_0_net469),
    .X(clknet_1_1__leaf_net469));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net455 (.A(net455),
    .X(clknet_0_net455));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net455 (.A(clknet_0_net455),
    .X(clknet_1_0__leaf_net455));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net455 (.A(clknet_0_net455),
    .X(clknet_1_1__leaf_net455));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net499 (.A(net499),
    .X(clknet_0_net499));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net499 (.A(clknet_0_net499),
    .X(clknet_1_0__leaf_net499));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net499 (.A(clknet_0_net499),
    .X(clknet_1_1__leaf_net499));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net502 (.A(net502),
    .X(clknet_0_net502));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net502 (.A(clknet_0_net502),
    .X(clknet_1_0__leaf_net502));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net502 (.A(clknet_0_net502),
    .X(clknet_1_1__leaf_net502));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net489 (.A(net489),
    .X(clknet_0_net489));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net489 (.A(clknet_0_net489),
    .X(clknet_1_0__leaf_net489));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net489 (.A(clknet_0_net489),
    .X(clknet_1_1__leaf_net489));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net458 (.A(net458),
    .X(clknet_0_net458));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net458 (.A(clknet_0_net458),
    .X(clknet_1_0__leaf_net458));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net458 (.A(clknet_0_net458),
    .X(clknet_1_1__leaf_net458));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net457 (.A(net457),
    .X(clknet_0_net457));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net457 (.A(clknet_0_net457),
    .X(clknet_1_0__leaf_net457));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net457 (.A(clknet_0_net457),
    .X(clknet_1_1__leaf_net457));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net463 (.A(net463),
    .X(clknet_0_net463));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net463 (.A(clknet_0_net463),
    .X(clknet_1_0__leaf_net463));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net463 (.A(clknet_0_net463),
    .X(clknet_1_1__leaf_net463));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net250 (.A(net250),
    .X(clknet_0_net250));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net250 (.A(clknet_0_net250),
    .X(clknet_1_0__leaf_net250));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net250 (.A(clknet_0_net250),
    .X(clknet_1_1__leaf_net250));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net456 (.A(net456),
    .X(clknet_0_net456));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net456 (.A(clknet_0_net456),
    .X(clknet_1_0__leaf_net456));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net456 (.A(clknet_0_net456),
    .X(clknet_1_1__leaf_net456));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net446 (.A(net446),
    .X(clknet_0_net446));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net446 (.A(clknet_0_net446),
    .X(clknet_1_0__leaf_net446));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net446 (.A(clknet_0_net446),
    .X(clknet_1_1__leaf_net446));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net481 (.A(net481),
    .X(clknet_0_net481));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net481 (.A(clknet_0_net481),
    .X(clknet_1_0__leaf_net481));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net481 (.A(clknet_0_net481),
    .X(clknet_1_1__leaf_net481));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net447 (.A(net447),
    .X(clknet_0_net447));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net447 (.A(clknet_0_net447),
    .X(clknet_1_0__leaf_net447));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net447 (.A(clknet_0_net447),
    .X(clknet_1_1__leaf_net447));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net443 (.A(net443),
    .X(clknet_0_net443));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net443 (.A(clknet_0_net443),
    .X(clknet_1_0__leaf_net443));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net443 (.A(clknet_0_net443),
    .X(clknet_1_1__leaf_net443));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net349 (.A(net349),
    .X(clknet_0_net349));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net349 (.A(clknet_0_net349),
    .X(clknet_1_0__leaf_net349));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net349 (.A(clknet_0_net349),
    .X(clknet_1_1__leaf_net349));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net674 (.A(net674),
    .X(clknet_0_net674));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net674 (.A(clknet_0_net674),
    .X(clknet_1_0__leaf_net674));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net674 (.A(clknet_0_net674),
    .X(clknet_1_1__leaf_net674));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net352 (.A(net352),
    .X(clknet_0_net352));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net352 (.A(clknet_0_net352),
    .X(clknet_1_0__leaf_net352));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net352 (.A(clknet_0_net352),
    .X(clknet_1_1__leaf_net352));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net523 (.A(net523),
    .X(clknet_0_net523));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net523 (.A(clknet_0_net523),
    .X(clknet_1_0__leaf_net523));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net523 (.A(clknet_0_net523),
    .X(clknet_1_1__leaf_net523));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net643 (.A(net643),
    .X(clknet_0_net643));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net643 (.A(clknet_0_net643),
    .X(clknet_1_0__leaf_net643));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net643 (.A(clknet_0_net643),
    .X(clknet_1_1__leaf_net643));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net528 (.A(net528),
    .X(clknet_0_net528));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net528 (.A(clknet_0_net528),
    .X(clknet_1_0__leaf_net528));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net528 (.A(clknet_0_net528),
    .X(clknet_1_1__leaf_net528));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net877 (.A(net877),
    .X(clknet_0_net877));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net877 (.A(clknet_0_net877),
    .X(clknet_1_0__leaf_net877));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net877 (.A(clknet_0_net877),
    .X(clknet_1_1__leaf_net877));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net358 (.A(net358),
    .X(clknet_0_net358));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net358 (.A(clknet_0_net358),
    .X(clknet_1_0__leaf_net358));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net358 (.A(clknet_0_net358),
    .X(clknet_1_1__leaf_net358));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net492 (.A(net492),
    .X(clknet_0_net492));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net492 (.A(clknet_0_net492),
    .X(clknet_1_0__leaf_net492));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net492 (.A(clknet_0_net492),
    .X(clknet_1_1__leaf_net492));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net509 (.A(net509),
    .X(clknet_0_net509));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net509 (.A(clknet_0_net509),
    .X(clknet_1_0__leaf_net509));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net509 (.A(clknet_0_net509),
    .X(clknet_1_1__leaf_net509));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net357 (.A(net357),
    .X(clknet_0_net357));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net357 (.A(clknet_0_net357),
    .X(clknet_1_0__leaf_net357));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net357 (.A(clknet_0_net357),
    .X(clknet_1_1__leaf_net357));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net353 (.A(net353),
    .X(clknet_0_net353));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net353 (.A(clknet_0_net353),
    .X(clknet_1_0__leaf_net353));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net353 (.A(clknet_0_net353),
    .X(clknet_1_1__leaf_net353));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net348 (.A(net348),
    .X(clknet_0_net348));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net348 (.A(clknet_0_net348),
    .X(clknet_1_0__leaf_net348));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net348 (.A(clknet_0_net348),
    .X(clknet_1_1__leaf_net348));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net370 (.A(net370),
    .X(clknet_0_net370));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net370 (.A(clknet_0_net370),
    .X(clknet_1_0__leaf_net370));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net370 (.A(clknet_0_net370),
    .X(clknet_1_1__leaf_net370));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net403 (.A(net403),
    .X(clknet_0_net403));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net403 (.A(clknet_0_net403),
    .X(clknet_1_0__leaf_net403));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net403 (.A(clknet_0_net403),
    .X(clknet_1_1__leaf_net403));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net366 (.A(net366),
    .X(clknet_0_net366));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net366 (.A(clknet_0_net366),
    .X(clknet_1_0__leaf_net366));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net366 (.A(clknet_0_net366),
    .X(clknet_1_1__leaf_net366));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net342 (.A(net342),
    .X(clknet_0_net342));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net342 (.A(clknet_0_net342),
    .X(clknet_1_0__leaf_net342));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net342 (.A(clknet_0_net342),
    .X(clknet_1_1__leaf_net342));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net444 (.A(net444),
    .X(clknet_0_net444));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net444 (.A(clknet_0_net444),
    .X(clknet_1_0__leaf_net444));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net444 (.A(clknet_0_net444),
    .X(clknet_1_1__leaf_net444));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net347 (.A(net347),
    .X(clknet_0_net347));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net347 (.A(clknet_0_net347),
    .X(clknet_1_0__leaf_net347));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net347 (.A(clknet_0_net347),
    .X(clknet_1_1__leaf_net347));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net343 (.A(net343),
    .X(clknet_0_net343));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net343 (.A(clknet_0_net343),
    .X(clknet_1_0__leaf_net343));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net343 (.A(clknet_0_net343),
    .X(clknet_1_1__leaf_net343));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net246 (.A(net246),
    .X(clknet_0_net246));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net246 (.A(clknet_0_net246),
    .X(clknet_1_0__leaf_net246));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net246 (.A(clknet_0_net246),
    .X(clknet_1_1__leaf_net246));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net673 (.A(net673),
    .X(clknet_0_net673));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net673 (.A(clknet_0_net673),
    .X(clknet_1_0__leaf_net673));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net673 (.A(clknet_0_net673),
    .X(clknet_1_1__leaf_net673));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net341 (.A(net341),
    .X(clknet_0_net341));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net341 (.A(clknet_0_net341),
    .X(clknet_1_0__leaf_net341));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net341 (.A(clknet_0_net341),
    .X(clknet_1_1__leaf_net341));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net367 (.A(net367),
    .X(clknet_0_net367));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net367 (.A(clknet_0_net367),
    .X(clknet_1_0__leaf_net367));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net367 (.A(clknet_0_net367),
    .X(clknet_1_1__leaf_net367));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net658 (.A(net658),
    .X(clknet_0_net658));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net658 (.A(clknet_0_net658),
    .X(clknet_1_0__leaf_net658));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net658 (.A(clknet_0_net658),
    .X(clknet_1_1__leaf_net658));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net907 (.A(net907),
    .X(clknet_0_net907));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net907 (.A(clknet_0_net907),
    .X(clknet_1_0__leaf_net907));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net907 (.A(clknet_0_net907),
    .X(clknet_1_1__leaf_net907));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net107 (.A(net107),
    .X(clknet_0_net107));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net107 (.A(clknet_0_net107),
    .X(clknet_1_0__leaf_net107));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net107 (.A(clknet_0_net107),
    .X(clknet_1_1__leaf_net107));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net318 (.A(net318),
    .X(clknet_0_net318));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net318 (.A(clknet_0_net318),
    .X(clknet_1_0__leaf_net318));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net318 (.A(clknet_0_net318),
    .X(clknet_1_1__leaf_net318));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net205 (.A(net205),
    .X(clknet_0_net205));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net205 (.A(clknet_0_net205),
    .X(clknet_1_0__leaf_net205));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net205 (.A(clknet_0_net205),
    .X(clknet_1_1__leaf_net205));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net109 (.A(net109),
    .X(clknet_0_net109));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net109 (.A(clknet_0_net109),
    .X(clknet_1_0__leaf_net109));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net109 (.A(clknet_0_net109),
    .X(clknet_1_1__leaf_net109));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net105 (.A(net105),
    .X(clknet_0_net105));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net105 (.A(clknet_0_net105),
    .X(clknet_1_0__leaf_net105));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net105 (.A(clknet_0_net105),
    .X(clknet_1_1__leaf_net105));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net921 (.A(net921),
    .X(clknet_0_net921));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net921 (.A(clknet_0_net921),
    .X(clknet_1_0__leaf_net921));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net921 (.A(clknet_0_net921),
    .X(clknet_1_1__leaf_net921));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net657 (.A(net657),
    .X(clknet_0_net657));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net657 (.A(clknet_0_net657),
    .X(clknet_1_0__leaf_net657));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net657 (.A(clknet_0_net657),
    .X(clknet_1_1__leaf_net657));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net656 (.A(net656),
    .X(clknet_0_net656));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net656 (.A(clknet_0_net656),
    .X(clknet_1_0__leaf_net656));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net656 (.A(clknet_0_net656),
    .X(clknet_1_1__leaf_net656));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net316 (.A(net316),
    .X(clknet_0_net316));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net316 (.A(clknet_0_net316),
    .X(clknet_1_0__leaf_net316));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net316 (.A(clknet_0_net316),
    .X(clknet_1_1__leaf_net316));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net644 (.A(net644),
    .X(clknet_0_net644));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net644 (.A(clknet_0_net644),
    .X(clknet_1_0__leaf_net644));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net644 (.A(clknet_0_net644),
    .X(clknet_1_1__leaf_net644));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net216 (.A(net216),
    .X(clknet_0_net216));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net216 (.A(clknet_0_net216),
    .X(clknet_1_0__leaf_net216));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net216 (.A(clknet_0_net216),
    .X(clknet_1_1__leaf_net216));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net912 (.A(net912),
    .X(clknet_0_net912));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net912 (.A(clknet_0_net912),
    .X(clknet_1_0__leaf_net912));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net912 (.A(clknet_0_net912),
    .X(clknet_1_1__leaf_net912));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net887 (.A(net887),
    .X(clknet_0_net887));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net887 (.A(clknet_0_net887),
    .X(clknet_1_0__leaf_net887));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net887 (.A(clknet_0_net887),
    .X(clknet_1_1__leaf_net887));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net319 (.A(net319),
    .X(clknet_0_net319));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net319 (.A(clknet_0_net319),
    .X(clknet_1_0__leaf_net319));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net319 (.A(clknet_0_net319),
    .X(clknet_1_1__leaf_net319));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net203 (.A(net203),
    .X(clknet_0_net203));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net203 (.A(clknet_0_net203),
    .X(clknet_1_0__leaf_net203));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net203 (.A(clknet_0_net203),
    .X(clknet_1_1__leaf_net203));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer1 (.A(net42),
    .X(net1027));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer2 (.A(net1027),
    .X(net1028));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer3 (.A(net1027),
    .X(net1029));
 sky130_fd_sc_hd__buf_2 rebuffer4 (.A(net1029),
    .X(net1030));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer5 (.A(net42),
    .X(net1031));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer6 (.A(net46),
    .X(net1032));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer7 (.A(net1032),
    .X(net1033));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer8 (.A(net1033),
    .X(net1034));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer9 (.A(net1136),
    .X(net1035));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer10 (.A(net48),
    .X(net1036));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer11 (.A(net1036),
    .X(net1037));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer12 (.A(net1039),
    .X(net1038));
 sky130_fd_sc_hd__mux4_1 clone13 (.A0(net1118),
    .A1(net1135),
    .A2(net1052),
    .A3(net1161),
    .S0(net1026),
    .S1(net1023),
    .X(net1039));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer14 (.A(net49),
    .X(net1040));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer15 (.A(net1040),
    .X(net1041));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer16 (.A(net879),
    .X(net1042));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer17 (.A(net1042),
    .X(net1043));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer18 (.A(net1043),
    .X(net1044));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer19 (.A(net1043),
    .X(net1045));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer20 (.A(net295),
    .X(net1046));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer21 (.A(net1046),
    .X(net1047));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer22 (.A(net295),
    .X(net1048));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer23 (.A(net1139),
    .X(net1049));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer24 (.A(net28),
    .X(net1050));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer25 (.A(net1052),
    .X(net1051));
 sky130_fd_sc_hd__mux4_1 clone26 (.A0(net1081),
    .A1(net24),
    .A2(net1132),
    .A3(net1160),
    .S0(net1117),
    .S1(net1121),
    .X(net1052));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer27 (.A(net47),
    .X(net1053));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer28 (.A(net1053),
    .X(net1054));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer29 (.A(net40),
    .X(net1055));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer30 (.A(net1055),
    .X(net1056));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer31 (.A(net30),
    .X(net1057));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer32 (.A(net23),
    .X(net1058));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer33 (.A(net32),
    .X(net1059));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer34 (.A(net137),
    .X(net1060));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer35 (.A(net1060),
    .X(net1061));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer36 (.A(net74),
    .X(net1062));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer37 (.A(net1062),
    .X(net1063));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer38 (.A(net31),
    .X(net1064));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer39 (.A(net128),
    .X(net1065));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer40 (.A(net128),
    .X(net1066));
 sky130_fd_sc_hd__dlygate4sd3_1 rebuffer41 (.A(net135),
    .X(net1067));
 sky130_fd_sc_hd__clkbuf_4 rebuffer42 (.A(net1067),
    .X(net1068));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer43 (.A(net1068),
    .X(net1069));
 sky130_fd_sc_hd__dlymetal6s4s_1 rebuffer44 (.A(net1067),
    .X(net1070));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer45 (.A(net134),
    .X(net1071));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer46 (.A(net1071),
    .X(net1072));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer47 (.A(net1072),
    .X(net1073));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer48 (.A(net134),
    .X(net1074));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer49 (.A(net188),
    .X(net1075));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer50 (.A(net190),
    .X(net1076));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer51 (.A(net133),
    .X(net1077));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer52 (.A(net1077),
    .X(net1078));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer53 (.A(net1077),
    .X(net1079));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer54 (.A(net26),
    .X(net1080));
 sky130_fd_sc_hd__clkbuf_1 clone55 (.A(net23),
    .X(net1081));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer56 (.A(net126),
    .X(net1082));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer57 (.A(net1082),
    .X(net1083));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer58 (.A(net1083),
    .X(net1084));
 sky130_fd_sc_hd__clkbuf_4 clone59 (.A(net40),
    .X(net1085));
 sky130_fd_sc_hd__clkbuf_1 clone60 (.A(net28),
    .X(net1086));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer61 (.A(net935),
    .X(net1087));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer62 (.A(net1087),
    .X(net1088));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer63 (.A(net935),
    .X(net1089));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer64 (.A(net955),
    .X(net1090));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer65 (.A(net1090),
    .X(net1091));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer66 (.A(net1090),
    .X(net1092));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer67 (.A(net1092),
    .X(net1093));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer68 (.A(net958),
    .X(net1094));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer69 (.A(net958),
    .X(net1095));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer70 (.A(net1095),
    .X(net1096));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer71 (.A(net1096),
    .X(net1097));
 sky130_fd_sc_hd__clkbuf_1 clone72 (.A(net30),
    .X(net1098));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer73 (.A(net193),
    .X(net1099));
 sky130_fd_sc_hd__a41o_1 clone74 (.A1(net971),
    .A2(net753),
    .A3(net18),
    .A4(net1160),
    .B1(net1121),
    .X(net1100));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer75 (.A(net978),
    .X(net1101));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer76 (.A(net1105),
    .X(net1102));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer77 (.A(net635),
    .X(net1103));
 sky130_fd_sc_hd__clkbuf_1 clone78 (.A(net27),
    .X(net1104));
 sky130_fd_sc_hd__clkbuf_1 clone79 (.A(net922),
    .X(net1105));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer80 (.A(net922),
    .X(net1106));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer81 (.A(net1106),
    .X(net1107));
 sky130_fd_sc_hd__clkbuf_4 clone82 (.A(net43),
    .X(net1108));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer83 (.A(net43),
    .X(net1109));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer84 (.A(net1109),
    .X(net1110));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer85 (.A(net1112),
    .X(net1111));
 sky130_fd_sc_hd__clkbuf_1 clone86 (.A(net35),
    .X(net1112));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer87 (.A(net974),
    .X(net1113));
 sky130_fd_sc_hd__clkbuf_1 clone88 (.A(net898),
    .X(net1114));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer89 (.A(net898),
    .X(net1115));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer90 (.A(net1013),
    .X(net1116));
 sky130_fd_sc_hd__clkbuf_1 clone91 (.A(net1011),
    .X(net1117));
 sky130_fd_sc_hd__clkbuf_1 clone92 (.A(net978),
    .X(net1118));
 sky130_fd_sc_hd__clkbuf_1 clone93 (.A(net945),
    .X(net1119));
 sky130_fd_sc_hd__clkbuf_1 clone94 (.A(net1013),
    .X(net1120));
 sky130_fd_sc_hd__clkbuf_1 clone95 (.A(net973),
    .X(net1121));
 sky130_fd_sc_hd__dlygate4sd3_1 hold96 (.A(net870),
    .X(net1122));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(net983),
    .X(net1123));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(net985),
    .X(net1124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(net982),
    .X(net1125));
 sky130_fd_sc_hd__dlygate4sd3_1 hold100 (.A(net749),
    .X(net1126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold101 (.A(net691),
    .X(net1127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold102 (.A(net654),
    .X(net1128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold103 (.A(net684),
    .X(net1129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold104 (.A(net632),
    .X(net1130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold105 (.A(net620),
    .X(net1131));
 sky130_fd_sc_hd__buf_12 fanout1 (.A(net975),
    .X(net1132));
 sky130_fd_sc_hd__clkbuf_1 fanout2 (.A(net1026),
    .X(net1133));
 sky130_fd_sc_hd__buf_4 fanout3 (.A(net1023),
    .X(net1134));
 sky130_fd_sc_hd__buf_8 fanout4 (.A(net992),
    .X(net1135));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_A (.DIODE(clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(in0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(in1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(in10));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(in11));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(in12));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(in13));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(in14));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(in15));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(in16));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(in17));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(in18));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(in19));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(in2));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(in20));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(in21));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(in22));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(in23));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(in24));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(in25));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(in26));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(in27));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_A (.DIODE(in28));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_A (.DIODE(in29));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_A (.DIODE(in3));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_A (.DIODE(in30));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_A (.DIODE(in31));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_A (.DIODE(in32));
 sky130_fd_sc_hd__diode_2 ANTENNA_input28_A (.DIODE(in33));
 sky130_fd_sc_hd__diode_2 ANTENNA_input29_A (.DIODE(in34));
 sky130_fd_sc_hd__diode_2 ANTENNA_input30_A (.DIODE(in35));
 sky130_fd_sc_hd__diode_2 ANTENNA_input31_A (.DIODE(in36));
 sky130_fd_sc_hd__diode_2 ANTENNA_input32_A (.DIODE(in37));
 sky130_fd_sc_hd__diode_2 ANTENNA_input33_A (.DIODE(in38));
 sky130_fd_sc_hd__diode_2 ANTENNA_input34_A (.DIODE(in39));
 sky130_fd_sc_hd__diode_2 ANTENNA_input35_A (.DIODE(in4));
 sky130_fd_sc_hd__diode_2 ANTENNA_input36_A (.DIODE(in40));
 sky130_fd_sc_hd__diode_2 ANTENNA_input37_A (.DIODE(in41));
 sky130_fd_sc_hd__diode_2 ANTENNA_input38_A (.DIODE(in42));
 sky130_fd_sc_hd__diode_2 ANTENNA_input39_A (.DIODE(in43));
 sky130_fd_sc_hd__diode_2 ANTENNA_input40_A (.DIODE(in44));
 sky130_fd_sc_hd__diode_2 ANTENNA_input41_A (.DIODE(in45));
 sky130_fd_sc_hd__diode_2 ANTENNA_input42_A (.DIODE(in46));
 sky130_fd_sc_hd__diode_2 ANTENNA_input43_A (.DIODE(in47));
 sky130_fd_sc_hd__diode_2 ANTENNA_input44_A (.DIODE(in48));
 sky130_fd_sc_hd__diode_2 ANTENNA_input45_A (.DIODE(in49));
 sky130_fd_sc_hd__diode_2 ANTENNA_input46_A (.DIODE(in5));
 sky130_fd_sc_hd__diode_2 ANTENNA_input47_A (.DIODE(in50));
 sky130_fd_sc_hd__diode_2 ANTENNA_input48_A (.DIODE(in51));
 sky130_fd_sc_hd__diode_2 ANTENNA_input49_A (.DIODE(in52));
 sky130_fd_sc_hd__diode_2 ANTENNA_input50_A (.DIODE(in53));
 sky130_fd_sc_hd__diode_2 ANTENNA_input51_A (.DIODE(in54));
 sky130_fd_sc_hd__diode_2 ANTENNA_input52_A (.DIODE(in55));
 sky130_fd_sc_hd__diode_2 ANTENNA_input53_A (.DIODE(in56));
 sky130_fd_sc_hd__diode_2 ANTENNA_input54_A (.DIODE(in57));
 sky130_fd_sc_hd__diode_2 ANTENNA_input55_A (.DIODE(in58));
 sky130_fd_sc_hd__diode_2 ANTENNA_input56_A (.DIODE(in59));
 sky130_fd_sc_hd__diode_2 ANTENNA_input57_A (.DIODE(in6));
 sky130_fd_sc_hd__diode_2 ANTENNA_input58_A (.DIODE(in60));
 sky130_fd_sc_hd__diode_2 ANTENNA_input59_A (.DIODE(in61));
 sky130_fd_sc_hd__diode_2 ANTENNA_input60_A (.DIODE(in62));
 sky130_fd_sc_hd__diode_2 ANTENNA_input61_A (.DIODE(in63));
 sky130_fd_sc_hd__diode_2 ANTENNA_input62_A (.DIODE(in64));
 sky130_fd_sc_hd__diode_2 ANTENNA_input63_A (.DIODE(in65));
 sky130_fd_sc_hd__diode_2 ANTENNA_input64_A (.DIODE(in66));
 sky130_fd_sc_hd__diode_2 ANTENNA_input65_A (.DIODE(in67));
 sky130_fd_sc_hd__diode_2 ANTENNA_input66_A (.DIODE(in68));
 sky130_fd_sc_hd__diode_2 ANTENNA_input67_A (.DIODE(in69));
 sky130_fd_sc_hd__diode_2 ANTENNA_input68_A (.DIODE(in7));
 sky130_fd_sc_hd__diode_2 ANTENNA_input69_A (.DIODE(in70));
 sky130_fd_sc_hd__diode_2 ANTENNA_input70_A (.DIODE(in71));
 sky130_fd_sc_hd__diode_2 ANTENNA_input71_A (.DIODE(in72));
 sky130_fd_sc_hd__diode_2 ANTENNA_input72_A (.DIODE(in73));
 sky130_fd_sc_hd__diode_2 ANTENNA_input73_A (.DIODE(in74));
 sky130_fd_sc_hd__diode_2 ANTENNA_input74_A (.DIODE(in75));
 sky130_fd_sc_hd__diode_2 ANTENNA_input75_A (.DIODE(in76));
 sky130_fd_sc_hd__diode_2 ANTENNA_input76_A (.DIODE(in77));
 sky130_fd_sc_hd__diode_2 ANTENNA_input77_A (.DIODE(in78));
 sky130_fd_sc_hd__diode_2 ANTENNA_input78_A (.DIODE(in79));
 sky130_fd_sc_hd__diode_2 ANTENNA_input79_A (.DIODE(in8));
 sky130_fd_sc_hd__diode_2 ANTENNA_input80_A (.DIODE(in80));
 sky130_fd_sc_hd__diode_2 ANTENNA_input81_A (.DIODE(in81));
 sky130_fd_sc_hd__diode_2 ANTENNA_input82_A (.DIODE(in82));
 sky130_fd_sc_hd__diode_2 ANTENNA_input83_A (.DIODE(in83));
 sky130_fd_sc_hd__diode_2 ANTENNA_input84_A (.DIODE(in84));
 sky130_fd_sc_hd__diode_2 ANTENNA_input85_A (.DIODE(in85));
 sky130_fd_sc_hd__diode_2 ANTENNA_input86_A (.DIODE(in86));
 sky130_fd_sc_hd__diode_2 ANTENNA_input87_A (.DIODE(in87));
 sky130_fd_sc_hd__diode_2 ANTENNA_input88_A (.DIODE(in88));
 sky130_fd_sc_hd__diode_2 ANTENNA_input89_A (.DIODE(in89));
 sky130_fd_sc_hd__diode_2 ANTENNA_input90_A (.DIODE(in9));
 sky130_fd_sc_hd__diode_2 ANTENNA_input91_A (.DIODE(in90));
 sky130_fd_sc_hd__diode_2 ANTENNA_input92_A (.DIODE(in91));
 sky130_fd_sc_hd__diode_2 ANTENNA_input93_A (.DIODE(in92));
 sky130_fd_sc_hd__diode_2 ANTENNA_input94_A (.DIODE(in93));
 sky130_fd_sc_hd__diode_2 ANTENNA_input95_A (.DIODE(in94));
 sky130_fd_sc_hd__diode_2 ANTENNA_input96_A (.DIODE(in95));
 sky130_fd_sc_hd__diode_2 ANTENNA_input97_A (.DIODE(in96));
 sky130_fd_sc_hd__diode_2 ANTENNA_input98_A (.DIODE(in97));
 sky130_fd_sc_hd__diode_2 ANTENNA_input99_A (.DIODE(in98));
 sky130_fd_sc_hd__diode_2 ANTENNA_input100_A (.DIODE(in99));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_A0 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_S1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_S1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c271_A2 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c270_A4 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c269_A1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_A2 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c267_B1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c264_X (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_A0 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c558_A3 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c532_D (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c404_A4 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_A0 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_A4 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c273_A2 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c267_X (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_A0 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_A3 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c557_A2 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_A2 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_A1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_A3 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c270_A1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_X (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c340_A0 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_A3 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_A0 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_A4 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c276_A2 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c275_A4 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c274_A1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c270_X (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c672_A3 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c670_S0 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c667_A1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c662_S0 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c546_D (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c404_A2 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c279_A2 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c275_X (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_A0 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_c398_A3 (.DIODE(net1143));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_A0 (.DIODE(net1143));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_A2 (.DIODE(net1143));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_A3 (.DIODE(net1143));
 sky130_fd_sc_hd__diode_2 ANTENNA_c283_A0 (.DIODE(net1143));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_A2 (.DIODE(net1143));
 sky130_fd_sc_hd__diode_2 ANTENNA_c278_X (.DIODE(net1143));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_A2 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA_c530_A1 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_A3 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_A0 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_A3 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA_c279_X (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_A0 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_c544_A1 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_A1 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_A0 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_X (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_c559_S0 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_A0 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_S0 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_S0 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_c286_X (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_A2 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_c614_A2 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_c556_S1 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_A0 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_A0 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_A0 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_A2 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_B1 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_c295_A2 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_X (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_A0 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_A2 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_c587_S0 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_c555_A1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_A2 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_A3 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_A3 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_A2 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_X (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_A0 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_A1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_A1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_S0 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_A1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_X (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c370_A1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_S0 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_A2 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_SCD (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA_c295_A3 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_A0 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_X (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_A0 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_A2 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_A1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_S0 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_S0 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_A0 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_S1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_X (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_A2 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_A4 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_A2 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_A3 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_S0 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_Q_N (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_A0 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_A1 (.DIODE(net1142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c279_A4 (.DIODE(net1142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c265_A2 (.DIODE(net1142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_A2 (.DIODE(net1142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_A3 (.DIODE(net1142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_A2 (.DIODE(net1142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_A1 (.DIODE(net1142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_X (.DIODE(net1142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_A2 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_A2 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_c561_A1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_c554_A1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_A3 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_A2 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_c311_A1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_A2 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_A2 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_A0 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_c297_X (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_c700_A0 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_A3 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_A0 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_A3 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_A0 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_S0 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_X (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_A0 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_c703_A1 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_A3 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_S1 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_A2 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_X (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_c496_A0 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA_c494_A2 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_A0 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA_c446_A0 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_A4 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_A2 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_X (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA_c564_A1 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA_c562_A2 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA_c556_A0 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_A0 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_X (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_A0 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_A3 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_A2 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_X (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout230_A (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c428_A2 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_A4 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_X (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_A0 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_A1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_S1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_A0 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_A1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_A1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c323_A3 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_A2 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_A3 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_X (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_A1 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_A2 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_A3 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_A1 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_A0 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_A1 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_A2 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_A1 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_X (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA_c366_A0 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_S0 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_A1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_A2 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_A2 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_A0 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA_c321_A2 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_S0 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_S0 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA_c313_A1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_X (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_A1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_A3 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_A0 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_A1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA_c321_A0 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_A1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_X (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_A0 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_A0 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_X (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA_c138_A1 (.DIODE(net1141));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_A0 (.DIODE(net1141));
 sky130_fd_sc_hd__diode_2 ANTENNA_c264_A4 (.DIODE(net1141));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_A1 (.DIODE(net1141));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_A0 (.DIODE(net1141));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_S0 (.DIODE(net1141));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_A1 (.DIODE(net1141));
 sky130_fd_sc_hd__diode_2 ANTENNA_c136_A1 (.DIODE(net1141));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_X (.DIODE(net1141));
 sky130_fd_sc_hd__diode_2 ANTENNA_c582_A3 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_A3 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_A0 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_A1 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_A3 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_A3 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA_c321_S0 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_X (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_A0 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_c364_A1 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_A3 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_A1 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_A1 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_A1 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_X (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_A0 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_A0 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_A0 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_A3 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA_c346_A1 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_A3 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_A0 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_A2 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_X (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_A0 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_A1 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_X (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone74_A3 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_A4 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_A0 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_A3 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_A1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_S0 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_A2 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_c143_A3 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_c140_B1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_c136_X (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A0 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA_c340_S0 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_X (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout229_A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A0 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c761_S0 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_X (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_A0 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_A1 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_A3 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA_c350_A3 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_A1 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA_c346_A2 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_X (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout226_A (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout225_A (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_X (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout224_A (.DIODE(net1156));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_A1 (.DIODE(net1156));
 sky130_fd_sc_hd__diode_2 ANTENNA_c582_A2 (.DIODE(net1156));
 sky130_fd_sc_hd__diode_2 ANTENNA_c140_X (.DIODE(net1156));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout191_A (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_A2 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_X (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_A0 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_A1 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA_c529_A2 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_A2 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA_c413_A1 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA_c405_SCD (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA_c403_A3 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA_c397_X (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_A0 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_A2 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA_c700_A2 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_A2 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA_c586_A1 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA_c554_A2 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_A3 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_S0 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_A3 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA_c404_A1 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA_c399_X (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_A1 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_A2 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_A1 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_A1 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_c412_A1 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_c406_D (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_c402_D (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_c401_X (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_c548_A0 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA_c408_D (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA_c406_SCD (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA_c403_A1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA_c402_Q (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone55_A (.DIODE(net1137));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer32_A (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout221_A (.DIODE(net1137));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_A3 (.DIODE(net1137));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_X (.DIODE(net1137));
 sky130_fd_sc_hd__diode_2 ANTENNA_c662_A0 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA_c415_RESET_B (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA_c409_RESET_B (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA_c407_RESET_B (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA_c405_Q (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA_c693_A1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_A3 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_c663_B1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_c531_A3 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_A3 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_c409_SET_B (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_c406_Q_N (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_c761_A0 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_A3 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA_c669_RESET_B (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_A3 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_A2 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_A3 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA_c416_A1 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA_c406_Q (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA_c586_A0 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_S0 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c424_A4 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c413_A2 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c408_SCD (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c407_Q_N (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_A0 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA_c555_S0 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_A1 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_A1 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_A2 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA_c411_A1 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA_c407_Q (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_A2 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c686_S0 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_S0 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c414_A1 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c411_A3 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c408_Q_N (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c765_A0 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_c739_S0 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_S0 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_A2 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_c410_A1 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_c408_Q (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_A2 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA_c561_A3 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_A3 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_A0 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA_c416_A3 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA_c409_Q_N (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_A2 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_A0 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA_c555_A3 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA_c531_A1 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_A2 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_A1 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA_c409_Q (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_A2 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_A4 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_A4 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_A2 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c416_S0 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c415_Q_N (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_A0 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_A2 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA_c554_A3 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_A2 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_A1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_A1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA_c415_Q (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA_c496_A1 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_c428_A3 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_A3 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_c424_A1 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_A2 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_A2 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_X (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_A2 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_A1 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA_c587_A3 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA_c554_S0 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_A3 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_A0 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA_c434_A2 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_A1 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA_c431_A0 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_X (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_A0 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_A1 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_A0 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_A2 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_A0 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_X (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout182_A (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_S0 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_S0 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A0 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA_c424_X (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_A0 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_A2 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_A0 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_A3 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_c428_X (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_A1 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_A0 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_A2 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_A3 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_A1 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_A2 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_c437_A0 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_X (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone78_A (.DIODE(net1138));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout216_A (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_S1 (.DIODE(net1138));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_A0 (.DIODE(net1138));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_X (.DIODE(net1138));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_A1 (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_A1 (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_A2 (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_A0 (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_X (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone60_A (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer24_A (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout220_A (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_X (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A1 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_A2 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_A0 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_A2 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_A2 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_S0 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_A2 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_A3 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_A2 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_A2 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_X (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_A1 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_A3 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA_c577_A1 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA_c458_A0 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_A1 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_X (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout215_A (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_A3 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_c760_A1 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_X (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer23_A (.DIODE(net1139));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer22_A (.DIODE(net1140));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer20_A (.DIODE(net1140));
 sky130_fd_sc_hd__diode_2 ANTENNA_c746_A0 (.DIODE(net1140));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_A3 (.DIODE(net1140));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_X (.DIODE(net1140));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_A0 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_A2 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_A3 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_A3 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_A3 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_A2 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_X (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA_c368_A0 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_A3 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_A1 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c221_A2 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c109_A3 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c106_A2 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c105_X (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone72_A (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer31_A (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout213_A (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_X (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_A2 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_A3 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA_c669_SCD (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA_c562_A0 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA_c538_SET_B (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA_c528_Q_N (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_A1 (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA_c702_A2 (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA_c663_A2 (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA_c543_A1 (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA_c540_A0 (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA_c528_Q (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA_c769_A2 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_A1 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_A3 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_A3 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_A0 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_A1 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_A2 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_B1 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_A3 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_X (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone86_A (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout214_A (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_c431_A1 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_A2 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_A0 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_A2 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_X (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net352_A (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA_c543_X (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net357_A (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA_c547_X (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_A1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_A1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c458_S0 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c434_A3 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_A1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c297_A2 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c184_S1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_A4 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_A3 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c159_B1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_X (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c557_A1 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_c554_A0 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_A1 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_A3 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_A0 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_A2 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_c159_X (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_c745_S0 (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_A0 (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_A3 (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_A1 (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_S0 (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_S0 (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_A2 (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_A2 (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_X (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_A0 (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_A2 (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_A1 (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_X (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout204_A (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_A0 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_A1 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_A3 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_X (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_A0 (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_A2 (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_A1 (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_A2 (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_X (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA_c764_A2 (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA_c759_A1 (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA_c615_A2 (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA_c611_A2 (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_A2 (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_A3 (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_X (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout198_A (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_A3 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_A2 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_A0 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_X (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer5_A (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer1_A (.DIODE(net1144));
 sky130_fd_sc_hd__diode_2 ANTENNA_c313_A3 (.DIODE(net1144));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_A1 (.DIODE(net1144));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_A1 (.DIODE(net1144));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_X (.DIODE(net1144));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer83_A (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone82_A (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout193_A (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_X (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer9_A (.DIODE(net1136));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_A2 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_c226_A2 (.DIODE(net1136));
 sky130_fd_sc_hd__diode_2 ANTENNA_c198_A0 (.DIODE(net1136));
 sky130_fd_sc_hd__diode_2 ANTENNA_c194_A3 (.DIODE(net1136));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_S0 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_A1 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_X (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_A0 (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_A2 (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA_c669_Q (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA_c739_A2 (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 ANTENNA_c696_A0 (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 ANTENNA_c691_X (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net481_A (.DIODE(net481));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_X (.DIODE(net481));
 sky130_fd_sc_hd__diode_2 ANTENNA_c769_A1 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_A0 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_A2 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_A1 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_A1 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_S0 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_X (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_A2 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_A1 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_A3 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_A0 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_A3 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_A1 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_A3 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_X (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_A0 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_A3 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_A3 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_c263_A3 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_c262_A0 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_c232_A2 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_S0 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_S0 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_X (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_A0 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_A2 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_A1 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_A1 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA_c238_A1 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA_c236_A1 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_A2 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_A2 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_A3 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_A4 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_X (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_A3 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_A0 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_A3 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_A1 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_A3 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_A1 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_A2 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA_c184_A3 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_X (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge795_Q_N (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_A3 (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA_c691_A2 (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA_c562_S0 (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA_c535_A4 (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap240_A (.DIODE(net566));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge799_Q (.DIODE(net566));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_S0 (.DIODE(net566));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_S0 (.DIODE(net566));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_A1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_c610_A0 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_A3 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_A2 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_c372_A0 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_c232_A1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_c220_A1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_c184_A1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_X (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge806_Q (.DIODE(net573));
 sky130_fd_sc_hd__diode_2 ANTENNA_c691_A3 (.DIODE(net573));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_A3 (.DIODE(net573));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_A3 (.DIODE(net573));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_S0 (.DIODE(net573));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_A3 (.DIODE(net573));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_S0 (.DIODE(net573));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge808_Q (.DIODE(net576));
 sky130_fd_sc_hd__diode_2 ANTENNA_c430_SCE (.DIODE(net576));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_S1 (.DIODE(net576));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_S1 (.DIODE(net576));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_A3 (.DIODE(net576));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_A0 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA_c203_A1 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_A3 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA_c190_A0 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA_c182_X (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge813_Q (.DIODE(net580));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_A4 (.DIODE(net580));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_S0 (.DIODE(net580));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_S1 (.DIODE(net580));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_S0 (.DIODE(net581));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_A3 (.DIODE(net581));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_A3 (.DIODE(net581));
 sky130_fd_sc_hd__diode_2 ANTENNA_c313_S1 (.DIODE(net581));
 sky130_fd_sc_hd__diode_2 ANTENNA_c311_B1 (.DIODE(net581));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_S1 (.DIODE(net581));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_S1 (.DIODE(net581));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_S0 (.DIODE(net581));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_S1 (.DIODE(net581));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_A1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_A2 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA_c198_S0 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_A0 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_X (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge839_Q (.DIODE(net605));
 sky130_fd_sc_hd__diode_2 ANTENNA_c610_S0 (.DIODE(net605));
 sky130_fd_sc_hd__diode_2 ANTENNA_c560_A3 (.DIODE(net605));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_S0 (.DIODE(net605));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_A3 (.DIODE(net605));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_S0 (.DIODE(net605));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_S0 (.DIODE(net605));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge840_Q_N (.DIODE(net606));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_A3 (.DIODE(net606));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_S0 (.DIODE(net606));
 sky130_fd_sc_hd__diode_2 ANTENNA_c428_B1 (.DIODE(net606));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge840_Q (.DIODE(net607));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_S1 (.DIODE(net607));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_S0 (.DIODE(net607));
 sky130_fd_sc_hd__diode_2 ANTENNA_c446_S0 (.DIODE(net607));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_S0 (.DIODE(net607));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_A0 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_A3 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_S1 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_A2 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA_c230_A3 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA_c226_A0 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_X (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA_c765_A2 (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA_c747_S1 (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_S1 (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_A3 (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_S0 (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge852_Q (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_A3 (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_A2 (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_S0 (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA_c494_S0 (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_S0 (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA_c763_A1 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_A1 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_S0 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_A1 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_S0 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_B1 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA_c237_A1 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_A0 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_S0 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_A2 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_X (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge858_Q (.DIODE(net622));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_A3 (.DIODE(net622));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_S1 (.DIODE(net622));
 sky130_fd_sc_hd__diode_2 ANTENNA_c373_A3 (.DIODE(net622));
 sky130_fd_sc_hd__diode_2 ANTENNA_c372_A3 (.DIODE(net622));
 sky130_fd_sc_hd__diode_2 ANTENNA_c364_S0 (.DIODE(net622));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge862_Q (.DIODE(net627));
 sky130_fd_sc_hd__diode_2 ANTENNA_c769_A3 (.DIODE(net627));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_S0 (.DIODE(net627));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_A3 (.DIODE(net627));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_S0 (.DIODE(net627));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_S1 (.DIODE(net627));
 sky130_fd_sc_hd__diode_2 ANTENNA_c587_S1 (.DIODE(net627));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge863_Q (.DIODE(net628));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_A3 (.DIODE(net628));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_S1 (.DIODE(net628));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_S1 (.DIODE(net628));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_A3 (.DIODE(net628));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_S1 (.DIODE(net628));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge868_Q (.DIODE(net637));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_A3 (.DIODE(net637));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_S0 (.DIODE(net637));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_A3 (.DIODE(net637));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_S1 (.DIODE(net637));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_S1 (.DIODE(net637));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_S0 (.DIODE(net637));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_S0 (.DIODE(net637));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_A3 (.DIODE(net637));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_S1 (.DIODE(net639));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_S0 (.DIODE(net639));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_A3 (.DIODE(net639));
 sky130_fd_sc_hd__diode_2 ANTENNA_c365_S1 (.DIODE(net639));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_S1 (.DIODE(net639));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge880_Q (.DIODE(net647));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_S1 (.DIODE(net647));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_S1 (.DIODE(net647));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_S1 (.DIODE(net647));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_S1 (.DIODE(net647));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_A4 (.DIODE(net647));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_S0 (.DIODE(net647));
 sky130_fd_sc_hd__diode_2 ANTENNA_s884_Q_N (.DIODE(net649));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_A3 (.DIODE(net649));
 sky130_fd_sc_hd__diode_2 ANTENNA_c190_S1 (.DIODE(net649));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_S1 (.DIODE(net649));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_B1 (.DIODE(net649));
 sky130_fd_sc_hd__diode_2 ANTENNA_c743_A1 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_S0 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_S1 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_A2 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_A1 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA_c191_A0 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA_c190_X (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA_s884_Q (.DIODE(net650));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_S1 (.DIODE(net650));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_S1 (.DIODE(net650));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_S1 (.DIODE(net650));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_S0 (.DIODE(net650));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_S1 (.DIODE(net650));
 sky130_fd_sc_hd__diode_2 ANTENNA_s885_Q_N (.DIODE(net651));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_A3 (.DIODE(net651));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_S0 (.DIODE(net651));
 sky130_fd_sc_hd__diode_2 ANTENNA_c239_S1 (.DIODE(net651));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_S1 (.DIODE(net651));
 sky130_fd_sc_hd__diode_2 ANTENNA_s885_Q (.DIODE(net652));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_S0 (.DIODE(net652));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_S0 (.DIODE(net652));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_S1 (.DIODE(net652));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_S0 (.DIODE(net652));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold102_A (.DIODE(net654));
 sky130_fd_sc_hd__diode_2 ANTENNA_s887_Q (.DIODE(net654));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_A3 (.DIODE(net654));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_S0 (.DIODE(net654));
 sky130_fd_sc_hd__diode_2 ANTENNA_c218_S0 (.DIODE(net654));
 sky130_fd_sc_hd__diode_2 ANTENNA_c216_S1 (.DIODE(net654));
 sky130_fd_sc_hd__diode_2 ANTENNA_c208_S1 (.DIODE(net654));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout235_A (.DIODE(net655));
 sky130_fd_sc_hd__diode_2 ANTENNA_c762_S0 (.DIODE(net655));
 sky130_fd_sc_hd__diode_2 ANTENNA_s888_Q (.DIODE(net655));
 sky130_fd_sc_hd__diode_2 ANTENNA_s892_Q_N (.DIODE(net659));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_A3 (.DIODE(net659));
 sky130_fd_sc_hd__diode_2 ANTENNA_c258_S0 (.DIODE(net659));
 sky130_fd_sc_hd__diode_2 ANTENNA_c235_S1 (.DIODE(net659));
 sky130_fd_sc_hd__diode_2 ANTENNA_c231_S1 (.DIODE(net659));
 sky130_fd_sc_hd__diode_2 ANTENNA_c371_A0 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_A2 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_A2 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_A2 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_A2 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_S0 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_c191_X (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_s893_Q_N (.DIODE(net660));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_A3 (.DIODE(net660));
 sky130_fd_sc_hd__diode_2 ANTENNA_c238_S1 (.DIODE(net660));
 sky130_fd_sc_hd__diode_2 ANTENNA_s895_Q (.DIODE(net663));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_S0 (.DIODE(net663));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_A3 (.DIODE(net663));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_S0 (.DIODE(net663));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_S1 (.DIODE(net663));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_A3 (.DIODE(net663));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_S0 (.DIODE(net663));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_S1 (.DIODE(net663));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_S0 (.DIODE(net663));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_S1 (.DIODE(net663));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout234_A (.DIODE(net664));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout233_A (.DIODE(net664));
 sky130_fd_sc_hd__diode_2 ANTENNA_s896_Q (.DIODE(net664));
 sky130_fd_sc_hd__diode_2 ANTENNA_s897_Q (.DIODE(net665));
 sky130_fd_sc_hd__diode_2 ANTENNA_c764_A3 (.DIODE(net665));
 sky130_fd_sc_hd__diode_2 ANTENNA_c759_S0 (.DIODE(net665));
 sky130_fd_sc_hd__diode_2 ANTENNA_c742_S0 (.DIODE(net665));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_S0 (.DIODE(net665));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_A3 (.DIODE(net665));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_B1 (.DIODE(net665));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_S1 (.DIODE(net665));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_S1 (.DIODE(net665));
 sky130_fd_sc_hd__diode_2 ANTENNA_s898_Q (.DIODE(net666));
 sky130_fd_sc_hd__diode_2 ANTENNA_c372_S1 (.DIODE(net666));
 sky130_fd_sc_hd__diode_2 ANTENNA_c366_S1 (.DIODE(net666));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_S1 (.DIODE(net666));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_S0 (.DIODE(net666));
 sky130_fd_sc_hd__diode_2 ANTENNA_c346_S1 (.DIODE(net666));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_S0 (.DIODE(net666));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_S0 (.DIODE(net666));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_A1 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA_c220_A3 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_A0 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA_c194_S0 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_A3 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_X (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA_s902_Q (.DIODE(net670));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_S0 (.DIODE(net670));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_S1 (.DIODE(net670));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_S0 (.DIODE(net670));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A3 (.DIODE(net670));
 sky130_fd_sc_hd__diode_2 ANTENNA_c633_S0 (.DIODE(net670));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_S1 (.DIODE(net670));
 sky130_fd_sc_hd__diode_2 ANTENNA_c610_S1 (.DIODE(net670));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_S1 (.DIODE(net670));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net675_A (.DIODE(net675));
 sky130_fd_sc_hd__diode_2 ANTENNA_s907_GCLK (.DIODE(net675));
 sky130_fd_sc_hd__diode_2 ANTENNA_s908_Q (.DIODE(net677));
 sky130_fd_sc_hd__diode_2 ANTENNA_c723_S0 (.DIODE(net677));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_A3 (.DIODE(net677));
 sky130_fd_sc_hd__diode_2 ANTENNA_c427_B1 (.DIODE(net677));
 sky130_fd_sc_hd__diode_2 ANTENNA_s909_Q_N (.DIODE(net678));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_S1 (.DIODE(net678));
 sky130_fd_sc_hd__diode_2 ANTENNA_c431_S1 (.DIODE(net678));
 sky130_fd_sc_hd__diode_2 ANTENNA_c424_B1 (.DIODE(net678));
 sky130_fd_sc_hd__diode_2 ANTENNA_s909_Q (.DIODE(net679));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_S0 (.DIODE(net679));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_A3 (.DIODE(net679));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_S1 (.DIODE(net679));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_S1 (.DIODE(net679));
 sky130_fd_sc_hd__diode_2 ANTENNA_c766_S0 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_A2 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_A3 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_A1 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_A2 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c371_A3 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_A0 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_S0 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c194_A0 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_X (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_s911_Q (.DIODE(net682));
 sky130_fd_sc_hd__diode_2 ANTENNA_c769_B1 (.DIODE(net682));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_S0 (.DIODE(net682));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_S0 (.DIODE(net682));
 sky130_fd_sc_hd__diode_2 ANTENNA_c434_S1 (.DIODE(net682));
 sky130_fd_sc_hd__diode_2 ANTENNA_c430_SET_B (.DIODE(net682));
 sky130_fd_sc_hd__diode_2 ANTENNA_s912_Q (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_S0 (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA_c696_A2 (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA_c687_A2 (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_A3 (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_S1 (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_S1 (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_S1 (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold103_A (.DIODE(net684));
 sky130_fd_sc_hd__diode_2 ANTENNA_s913_Q (.DIODE(net684));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_S1 (.DIODE(net684));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_S0 (.DIODE(net684));
 sky130_fd_sc_hd__diode_2 ANTENNA_c686_S1 (.DIODE(net684));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_A3 (.DIODE(net684));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_S0 (.DIODE(net684));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_S0 (.DIODE(net684));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_S1 (.DIODE(net684));
 sky130_fd_sc_hd__diode_2 ANTENNA_c437_S1 (.DIODE(net684));
 sky130_fd_sc_hd__diode_2 ANTENNA_s915_Q (.DIODE(net686));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_B1 (.DIODE(net686));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_S0 (.DIODE(net686));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_S1 (.DIODE(net686));
 sky130_fd_sc_hd__diode_2 ANTENNA_c446_S1 (.DIODE(net686));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_S1 (.DIODE(net686));
 sky130_fd_sc_hd__diode_2 ANTENNA_s918_Q (.DIODE(net690));
 sky130_fd_sc_hd__diode_2 ANTENNA_c763_S0 (.DIODE(net690));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_S1 (.DIODE(net690));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_S1 (.DIODE(net690));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_S1 (.DIODE(net690));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_S0 (.DIODE(net690));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_S1 (.DIODE(net690));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_S1 (.DIODE(net690));
 sky130_fd_sc_hd__diode_2 ANTENNA_s920_Q (.DIODE(net692));
 sky130_fd_sc_hd__diode_2 ANTENNA_c764_S0 (.DIODE(net692));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_S1 (.DIODE(net692));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_S0 (.DIODE(net692));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_S0 (.DIODE(net692));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_S0 (.DIODE(net692));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_S1 (.DIODE(net692));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_S1 (.DIODE(net692));
 sky130_fd_sc_hd__diode_2 ANTENNA_s932_Q (.DIODE(net708));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_S1 (.DIODE(net708));
 sky130_fd_sc_hd__diode_2 ANTENNA_c698_S0 (.DIODE(net708));
 sky130_fd_sc_hd__diode_2 ANTENNA_c577_S1 (.DIODE(net708));
 sky130_fd_sc_hd__diode_2 ANTENNA_s933_Q_N (.DIODE(net709));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_S0 (.DIODE(net709));
 sky130_fd_sc_hd__diode_2 ANTENNA_c703_S0 (.DIODE(net709));
 sky130_fd_sc_hd__diode_2 ANTENNA_c685_S1 (.DIODE(net709));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_S1 (.DIODE(net709));
 sky130_fd_sc_hd__diode_2 ANTENNA_c560_S0 (.DIODE(net709));
 sky130_fd_sc_hd__diode_2 ANTENNA_c557_S1 (.DIODE(net709));
 sky130_fd_sc_hd__diode_2 ANTENNA_c555_S1 (.DIODE(net709));
 sky130_fd_sc_hd__diode_2 ANTENNA_c554_S1 (.DIODE(net709));
 sky130_fd_sc_hd__diode_2 ANTENNA_s934_Q (.DIODE(net710));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_S0 (.DIODE(net710));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_S1 (.DIODE(net710));
 sky130_fd_sc_hd__diode_2 ANTENNA_c696_A3 (.DIODE(net710));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_S0 (.DIODE(net710));
 sky130_fd_sc_hd__diode_2 ANTENNA_s935_Q (.DIODE(net711));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_S0 (.DIODE(net711));
 sky130_fd_sc_hd__diode_2 ANTENNA_c693_A3 (.DIODE(net711));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_S0 (.DIODE(net711));
 sky130_fd_sc_hd__diode_2 ANTENNA_c687_A3 (.DIODE(net711));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_S1 (.DIODE(net711));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net714_A (.DIODE(net714));
 sky130_fd_sc_hd__diode_2 ANTENNA_s938_GCLK (.DIODE(net714));
 sky130_fd_sc_hd__diode_2 ANTENNA_s940_Q (.DIODE(net717));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_S1 (.DIODE(net717));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_A4 (.DIODE(net717));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_S0 (.DIODE(net717));
 sky130_fd_sc_hd__diode_2 ANTENNA_s942_Q_N (.DIODE(net720));
 sky130_fd_sc_hd__diode_2 ANTENNA_c687_S0 (.DIODE(net720));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_S1 (.DIODE(net720));
 sky130_fd_sc_hd__diode_2 ANTENNA_c571_S1 (.DIODE(net720));
 sky130_fd_sc_hd__diode_2 ANTENNA_s942_Q (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_S0 (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_S1 (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_A3 (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_S1 (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA_s943_Q (.DIODE(net722));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_S1 (.DIODE(net722));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_S1 (.DIODE(net722));
 sky130_fd_sc_hd__diode_2 ANTENNA_c586_A3 (.DIODE(net722));
 sky130_fd_sc_hd__diode_2 ANTENNA_s948_Q_N (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA_c762_S1 (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_S1 (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_S0 (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA_s948_Q (.DIODE(net726));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_S0 (.DIODE(net726));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_A3 (.DIODE(net726));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_S1 (.DIODE(net726));
 sky130_fd_sc_hd__diode_2 ANTENNA_s952_Q (.DIODE(net731));
 sky130_fd_sc_hd__diode_2 ANTENNA_c760_S1 (.DIODE(net731));
 sky130_fd_sc_hd__diode_2 ANTENNA_c759_S1 (.DIODE(net731));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_S1 (.DIODE(net731));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_S1 (.DIODE(net731));
 sky130_fd_sc_hd__diode_2 ANTENNA_s961_Q (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA_c764_S1 (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA_c742_S1 (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_S0 (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA_c687_S1 (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA_s964_Q (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA_c767_S1 (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA_c765_S1 (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_S1 (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA_c700_S1 (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_S1 (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_A3 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_A0 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_S0 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_A0 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_A3 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_A1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_X (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_A1 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_A3 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_c371_A1 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_S0 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_A2 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_A0 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_S0 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_A2 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_X (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_c765_A1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_A0 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_A2 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_A2 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_A1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_A2 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_A2 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_A3 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_X (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c502_A0 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_A1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_c370_S0 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_A3 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_c206_A1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_c205_A2 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_c203_X (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_A1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_A3 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_A3 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_A0 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_c208_X (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout183_A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_A2 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_c218_X (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_A0 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_c369_A1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_c366_A1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_A2 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_A2 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_X (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_A1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_A0 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_A3 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_c240_A2 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_c236_A0 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_A2 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_c232_A0 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_X (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_A0 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA_c502_A3 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_A2 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_A2 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_A3 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA_c226_X (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout276_A (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_X (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_A0 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_A2 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_A0 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_A1 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout266_A (.DIODE(net752));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_X (.DIODE(net752));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_A1 (.DIODE(net752));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone74_A2 (.DIODE(net753));
 sky130_fd_sc_hd__diode_2 ANTENNA_c143_A2 (.DIODE(net753));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_X (.DIODE(net753));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_A0 (.DIODE(net753));
 sky130_fd_sc_hd__diode_2 ANTENNA_c403_A2 (.DIODE(net753));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_S1 (.DIODE(net753));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_A1 (.DIODE(net753));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_A3 (.DIODE(net753));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_A1 (.DIODE(net753));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_A1 (.DIODE(net753));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout256_A (.DIODE(net754));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_X (.DIODE(net754));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_A2 (.DIODE(net754));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_S0 (.DIODE(net754));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_A3 (.DIODE(net754));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout254_A (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout253_A (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_X (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_A3 (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_X (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA_c412_A0 (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_A3 (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA_c275_A2 (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_A2 (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_A0 (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_A2 (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA_c134_A2 (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout248_A (.DIODE(net757));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_X (.DIODE(net757));
 sky130_fd_sc_hd__diode_2 ANTENNA_c760_A0 (.DIODE(net757));
 sky130_fd_sc_hd__diode_2 ANTENNA_c759_A3 (.DIODE(net757));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_A3 (.DIODE(net757));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_S1 (.DIODE(net757));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout245_A (.DIODE(net758));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout244_A (.DIODE(net758));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_X (.DIODE(net758));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout243_A (.DIODE(net759));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_X (.DIODE(net759));
 sky130_fd_sc_hd__diode_2 ANTENNA_c537_A0 (.DIODE(net759));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout275_A (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_X (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_A2 (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_S0 (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_A3 (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_A3 (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout274_A (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_X (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_c239_S0 (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout273_A (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_X (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_A0 (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA_c400_B1 (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout272_A (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_X (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_A0 (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_A1 (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_S0 (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout271_A (.DIODE(net764));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_X (.DIODE(net764));
 sky130_fd_sc_hd__diode_2 ANTENNA_c365_A2 (.DIODE(net764));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_A2 (.DIODE(net764));
 sky130_fd_sc_hd__diode_2 ANTENNA_c231_A2 (.DIODE(net764));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_A1 (.DIODE(net764));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout270_A (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_X (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_A1 (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_c615_A1 (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_c502_S1 (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_A3 (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_X (.DIODE(net766));
 sky130_fd_sc_hd__diode_2 ANTENNA_c297_A3 (.DIODE(net766));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_SCE (.DIODE(net766));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_S0 (.DIODE(net766));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_A1 (.DIODE(net766));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_A3 (.DIODE(net766));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_X (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_A0 (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_A3 (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_c216_A2 (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_A3 (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_c108_A1 (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout269_A (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_X (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_A3 (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout268_A (.DIODE(net769));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout267_A (.DIODE(net769));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_X (.DIODE(net769));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_X (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_c208_A0 (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_c184_A0 (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_S1 (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_A2 (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_A1 (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_X (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_A0 (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_A3 (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_A0 (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_S0 (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_A3 (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_A2 (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_X (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_S0 (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA_c323_A1 (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_A1 (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_A1 (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_S0 (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA_c116_B1 (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout265_A (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout263_A (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_X (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A3 (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout259_A (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_X (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_c757_A1 (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_X (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_A0 (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_S0 (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_A3 (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c260_A0 (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c256_S1 (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c226_S0 (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c111_A1 (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_X (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_A0 (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_A1 (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_c696_A1 (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_A2 (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_A1 (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_input28_X (.DIODE(net778));
 sky130_fd_sc_hd__diode_2 ANTENNA_c558_A2 (.DIODE(net778));
 sky130_fd_sc_hd__diode_2 ANTENNA_c557_A0 (.DIODE(net778));
 sky130_fd_sc_hd__diode_2 ANTENNA_c424_A3 (.DIODE(net778));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_A2 (.DIODE(net778));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_A4 (.DIODE(net778));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_S1 (.DIODE(net778));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_S1 (.DIODE(net778));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_A1 (.DIODE(net778));
 sky130_fd_sc_hd__diode_2 ANTENNA_input30_X (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_S0 (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_A0 (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_A3 (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_A1 (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_A1 (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA_input31_X (.DIODE(net781));
 sky130_fd_sc_hd__diode_2 ANTENNA_c458_A2 (.DIODE(net781));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_A0 (.DIODE(net781));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_A0 (.DIODE(net781));
 sky130_fd_sc_hd__diode_2 ANTENNA_c313_A2 (.DIODE(net781));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_A3 (.DIODE(net781));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout258_A (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_input32_X (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_A0 (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_input33_X (.DIODE(net783));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_A0 (.DIODE(net783));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_A1 (.DIODE(net783));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_A3 (.DIODE(net783));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_A1 (.DIODE(net783));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_A3 (.DIODE(net783));
 sky130_fd_sc_hd__diode_2 ANTENNA_input34_X (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA_c194_A2 (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_S0 (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_A1 (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_A1 (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA_c158_B1 (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout257_A (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_input35_X (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_c768_A1 (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_A2 (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_c702_A3 (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_input36_X (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_A1 (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_S0 (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A1 (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_A2 (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_c557_A3 (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_A1 (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_S1 (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_S0 (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_c263_S0 (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_S0 (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_input37_X (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_A3 (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_A0 (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_S0 (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_B1 (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_A3 (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_A1 (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_A2 (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c121_A3 (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_input38_X (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_A1 (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_A0 (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_A2 (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_A0 (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_A2 (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_A3 (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA_input39_X (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_A0 (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_A1 (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_A1 (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_A2 (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_A3 (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_S1 (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_A1 (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_A3 (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_input40_X (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_A0 (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA_c321_A1 (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_A2 (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_A1 (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA_c180_A3 (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA_input41_X (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_c759_A0 (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_A1 (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_A2 (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_A2 (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_S0 (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_S0 (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_A2 (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_A3 (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_input42_X (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_A0 (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_A2 (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_A0 (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_c458_A1 (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_A2 (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_c344_A2 (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_c212_A1 (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_A1 (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_input44_X (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_A0 (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_S0 (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_A1 (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_A3 (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_c183_S0 (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_A1 (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout255_A (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA_input46_X (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA_c764_A1 (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA_input48_X (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_A1 (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA_c313_S0 (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_S0 (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_A3 (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA_c122_A2 (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA_input49_X (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c365_A1 (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_A0 (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_A1 (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_A1 (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_S0 (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_A1 (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c106_S0 (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_input50_X (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_A0 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_A2 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_A3 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_A2 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c183_A3 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_A1 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_A2 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_input53_X (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_A2 (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_A1 (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_A2 (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_A1 (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_A1 (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_S0 (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_A2 (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_S1 (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA_c126_A2 (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA_input54_X (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c344_S0 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c124_A3 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c120_A4 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c119_B1 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c117_S1 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c110_A2 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_input55_X (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_A2 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_A3 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_c577_A2 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_S0 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_A3 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_c230_A0 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_S1 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_c129_B1 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_c113_B1 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_c111_A3 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout252_A (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout251_A (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_input57_X (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_input58_X (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_A2 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c311_A2 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_A0 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_S0 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c182_A2 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_A3 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_input59_X (.DIODE(net809));
 sky130_fd_sc_hd__diode_2 ANTENNA_c261_A0 (.DIODE(net809));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_A1 (.DIODE(net809));
 sky130_fd_sc_hd__diode_2 ANTENNA_c180_A4 (.DIODE(net809));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_S0 (.DIODE(net809));
 sky130_fd_sc_hd__diode_2 ANTENNA_c122_A1 (.DIODE(net809));
 sky130_fd_sc_hd__diode_2 ANTENNA_input60_X (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_A1 (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_S0 (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_A2 (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_A3 (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_S0 (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_A2 (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_c369_A0 (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_S1 (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_A0 (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_A1 (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_input62_X (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_A0 (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_S0 (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_A2 (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_c183_A2 (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_c180_A2 (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_input67_X (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_S1 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_A2 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c257_S1 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_A2 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_A1 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c119_A3 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c115_A1 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c111_A2 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c107_S0 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout250_A (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout249_A (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_input68_X (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_input69_X (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_c502_A1 (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_A1 (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_A0 (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_A1 (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_c120_B1 (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_c118_A0 (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_c113_A2 (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_c101_S1 (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_c100_S1 (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_input71_X (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_A0 (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_A2 (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_A3 (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_A1 (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_c236_A2 (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_A1 (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_c108_S0 (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_input73_X (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_A0 (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_A1 (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_A3 (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_A2 (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_A1 (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_A0 (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_S1 (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_A1 (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_c205_A0 (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_input74_X (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_c742_A3 (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_A1 (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_A2 (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_A2 (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_S0 (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_A3 (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_A1 (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_A0 (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_c203_A2 (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_input75_X (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_c260_A1 (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_c257_A0 (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_c240_A3 (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_c234_A3 (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_c220_A2 (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_c126_S0 (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_c104_S1 (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout247_A (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout246_A (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_input79_X (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_input82_X (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c766_A1 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A1 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_A0 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_A3 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c611_A3 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_A0 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_A2 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_A2 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_A2 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_input83_X (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_c127_A3 (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_c125_S0 (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_c121_A1 (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_c114_B1 (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_c113_A3 (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_c102_S0 (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout242_A (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_input90_X (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_S0 (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_c434_A0 (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_c427_A4 (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_A3 (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_input92_X (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_A2 (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_A2 (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_A1 (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_A3 (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_c107_A0 (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_c105_A3 (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_c103_A2 (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_c102_A1 (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_c101_S0 (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_input93_X (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_A2 (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_A0 (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_A3 (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c222_S0 (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c105_A1 (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c103_A0 (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c102_A2 (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c101_A2 (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c100_A1 (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_input94_X (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_A3 (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_A3 (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_A3 (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_S0 (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c262_A2 (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c115_A3 (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c108_A3 (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c106_A1 (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c105_S0 (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c103_S0 (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_input95_X (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_A2 (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_S0 (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_S1 (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_A1 (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_c260_A2 (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_c124_S0 (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_input99_X (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c368_A3 (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_A0 (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_A3 (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c108_A2 (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_output102_A (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_s947_Q (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_S1 (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_S1 (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_output103_A (.DIODE(net853));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge861_Q (.DIODE(net853));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_A3 (.DIODE(net853));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_A3 (.DIODE(net853));
 sky130_fd_sc_hd__diode_2 ANTENNA_output104_A (.DIODE(net854));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_A1 (.DIODE(net854));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_A2 (.DIODE(net854));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_X (.DIODE(net854));
 sky130_fd_sc_hd__diode_2 ANTENNA_output105_A (.DIODE(net855));
 sky130_fd_sc_hd__diode_2 ANTENNA_s933_Q (.DIODE(net855));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_S0 (.DIODE(net855));
 sky130_fd_sc_hd__diode_2 ANTENNA_c744_S1 (.DIODE(net855));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_S0 (.DIODE(net855));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_S1 (.DIODE(net855));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_A3 (.DIODE(net855));
 sky130_fd_sc_hd__diode_2 ANTENNA_c565_A2 (.DIODE(net855));
 sky130_fd_sc_hd__diode_2 ANTENNA_c563_A3 (.DIODE(net855));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_S1 (.DIODE(net855));
 sky130_fd_sc_hd__diode_2 ANTENNA_output106_A (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge881_Q (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_c746_S1 (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_c633_A3 (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_S0 (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_output108_A (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_c743_A2 (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_A1 (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_A1 (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_A2 (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_X (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_output110_A (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_s967_Q (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_c720_S1 (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_S1 (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout190_A (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_output111_A (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_c434_X (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_output112_A (.DIODE(net862));
 sky130_fd_sc_hd__diode_2 ANTENNA_c559_A2 (.DIODE(net862));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_A3 (.DIODE(net862));
 sky130_fd_sc_hd__diode_2 ANTENNA_c494_A3 (.DIODE(net862));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_A1 (.DIODE(net862));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_A2 (.DIODE(net862));
 sky130_fd_sc_hd__diode_2 ANTENNA_c323_A0 (.DIODE(net862));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_X (.DIODE(net862));
 sky130_fd_sc_hd__diode_2 ANTENNA_output113_A (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge872_Q (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_c760_A3 (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_A3 (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_c614_S0 (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_output114_A (.DIODE(net864));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_A1 (.DIODE(net864));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_S0 (.DIODE(net864));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_X (.DIODE(net864));
 sky130_fd_sc_hd__diode_2 ANTENNA_output115_A (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge812_Q (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_S0 (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout212_A (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_A1 (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_A0 (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_X (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_output119_A (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_A2 (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_S0 (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_A3 (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_c228_A1 (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_c191_A1 (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_c183_X (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold96_A (.DIODE(net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_output120_A (.DIODE(net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_s892_Q (.DIODE(net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_c261_S0 (.DIODE(net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_c237_S1 (.DIODE(net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_S1 (.DIODE(net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_output122_A (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_A3 (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_A1 (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_A3 (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_A3 (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_c586_X (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_output123_A (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_A3 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_A1 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_A2 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_A1 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_A1 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_A2 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_A1 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_A2 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_A3 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_X (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_output124_A (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_A1 (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_A1 (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_c536_A1 (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_c533_X (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_output125_A (.DIODE(net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_s944_Q (.DIODE(net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_S1 (.DIODE(net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_S1 (.DIODE(net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_output130_A (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge793_Q (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_S0 (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_S0 (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_output131_A (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge851_Q (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_A2 (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_S1 (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_output133_A (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge847_Q_N (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_S1 (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_output134_A (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_A2 (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_c350_A2 (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_S0 (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_c215_X (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_output135_A (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_A3 (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_A1 (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_A0 (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_A2 (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_A2 (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_c313_X (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_output136_A (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_S0 (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_c261_A2 (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_S0 (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_A3 (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_S1 (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_B1 (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_A3 (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_S1 (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_c190_S0 (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_output138_A (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_c402_RESET_B (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_A1 (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_A3 (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_c277_A1 (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_c269_A3 (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_c266_A2 (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_c265_X (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_output139_A (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_s901_Q (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_S1 (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_S1 (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_output140_A (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_A3 (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c226_A1 (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c131_A3 (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c109_S1 (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c108_S1 (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c107_X (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_output141_A (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge880_Q_N (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c368_S1 (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_A3 (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_S0 (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_S1 (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_S1 (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_output143_A (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_s916_Q (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_S1 (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_S1 (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_output144_A (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge847_Q (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_S1 (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_output145_A (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_s899_Q (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_S0 (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_c364_S1 (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_S1 (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_output146_A (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_A0 (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_S1 (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_X (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_output147_A (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_A2 (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_A0 (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_A3 (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_X (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_output152_A (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge882_Q (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_S1 (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_S0 (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_A3 (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_c496_A3 (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_c369_S0 (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_c236_S0 (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_output153_A (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_A1 (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_A1 (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_c236_A3 (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_c110_A3 (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_c102_X (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_output154_A (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge818_Q (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_A2 (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_S0 (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_A3 (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_output155_A (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_A2 (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c258_A1 (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c256_S0 (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c228_S0 (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c222_A3 (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c109_X (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_output161_A (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_A2 (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_c297_S0 (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_A2 (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_A2 (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_S0 (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_A1 (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_X (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_output166_A (.DIODE(net916));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge821_Q (.DIODE(net916));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_A3 (.DIODE(net916));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_A3 (.DIODE(net916));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_A3 (.DIODE(net916));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_S0 (.DIODE(net916));
 sky130_fd_sc_hd__diode_2 ANTENNA_c365_A3 (.DIODE(net916));
 sky130_fd_sc_hd__diode_2 ANTENNA_output168_A (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_A0 (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_c259_A1 (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_c222_X (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_output170_A (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge870_Q (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_A3 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_S0 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_c366_S0 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_c262_A3 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_c261_A3 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer80_A (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone79_A (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout241_A (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_c134_X (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_output175_A (.DIODE(net925));
 sky130_fd_sc_hd__diode_2 ANTENNA_c260_A3 (.DIODE(net925));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_A1 (.DIODE(net925));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_S0 (.DIODE(net925));
 sky130_fd_sc_hd__diode_2 ANTENNA_c116_A3 (.DIODE(net925));
 sky130_fd_sc_hd__diode_2 ANTENNA_c103_X (.DIODE(net925));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout182_X (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_A3 (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_A1 (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_c431_A2 (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_c555_A2 (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_A2 (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_S0 (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_A3 (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_c430_RESET_B (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_A2 (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_A3 (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout183_X (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c494_A0 (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c371_S0 (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_S0 (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_S0 (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c231_S0 (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c230_A2 (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_A0 (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_A3 (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_A2 (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_A2 (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout184_X (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_A3 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_A1 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c665_A1 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_A3 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_S1 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c414_A2 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c406_SET_B (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c403_S1 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c401_A4 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c400_A3 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer63_A (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer61_A (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout185_X (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_S1 (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_A2 (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_S0 (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c205_A1 (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c221_A3 (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout186_X (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c566_A2 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c678_SCE (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c747_A3 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_A2 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_A3 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_A2 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_B1 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_S0 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c283_A2 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_A0 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout187_X (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_A1 (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_A3 (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_S0 (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_c412_A3 (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_c400_A2 (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_c399_A4 (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_c283_S0 (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_A2 (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_c397_A4 (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_A2 (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout188_X (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_A1 (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_c670_S1 (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_c668_A0 (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_c666_SCD (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_c664_A4 (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_c661_A1 (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_c660_B1 (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_c408_SCE (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_c533_A4 (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_c530_B1 (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout189_X (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout188_A (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c674_SCE (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_A3 (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_A2 (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_S0 (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_A0 (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout187_A (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout190_X (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_A3 (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_c611_A0 (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_c571_A1 (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_A2 (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_c566_A1 (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_A1 (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_S0 (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_c437_A3 (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_A1 (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_A1 (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout191_X (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_A2 (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_A0 (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_A2 (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c482_A0 (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_A1 (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_A1 (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c409_SCE (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c404_B1 (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c400_A1 (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c398_A1 (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout192_X (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_S1 (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_A1 (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_A3 (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_S0 (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_S0 (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_A1 (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_S1 (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_A3 (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c277_B1 (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_S0 (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout193_X (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_S0 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_A4 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_A1 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c191_S0 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_A2 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout196_X (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c679_A0 (.DIODE(net1158));
 sky130_fd_sc_hd__diode_2 ANTENNA_c661_S0 (.DIODE(net1158));
 sky130_fd_sc_hd__diode_2 ANTENNA_c549_S0 (.DIODE(net1158));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout195_A (.DIODE(net1158));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_A3 (.DIODE(net1158));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_A4 (.DIODE(net1158));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout197_X (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_S0 (.DIODE(net1149));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_A2 (.DIODE(net1149));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_A1 (.DIODE(net1149));
 sky130_fd_sc_hd__diode_2 ANTENNA_c364_A2 (.DIODE(net1149));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_A0 (.DIODE(net1149));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout196_A (.DIODE(net1149));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout198_X (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_A1 (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_A1 (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_A3 (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_A2 (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c286_A2 (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_A3 (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c198_A3 (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_A0 (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_A3 (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_A4 (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout201_X (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_A2 (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_A1 (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_A1 (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_A2 (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout200_A (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_c529_B1 (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_c273_A3 (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout202_X (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c743_S1 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_A1 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_A0 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c677_A3 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c539_A2 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c530_A2 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout201_A (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout204_X (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_S0 (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c437_A2 (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c561_A0 (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_A1 (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_B1 (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c321_A3 (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_A4 (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_A2 (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_A3 (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_A0 (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c271_A1 (.DIODE(net1147));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer64_A (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout205_X (.DIODE(net1147));
 sky130_fd_sc_hd__diode_2 ANTENNA_c587_A1 (.DIODE(net1147));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_S1 (.DIODE(net1147));
 sky130_fd_sc_hd__diode_2 ANTENNA_c532_SCD (.DIODE(net1147));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_S1 (.DIODE(net1147));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_B1 (.DIODE(net1147));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout206_X (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_A1 (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_c237_A2 (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_c226_A3 (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_A0 (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_A0 (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer69_A (.DIODE(net1146));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer68_A (.DIODE(net1146));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout208_X (.DIODE(net1146));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_A2 (.DIODE(net1146));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_A3 (.DIODE(net1146));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_S0 (.DIODE(net1146));
 sky130_fd_sc_hd__diode_2 ANTENNA_c398_A2 (.DIODE(net1146));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_A0 (.DIODE(net1146));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout209_X (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_A0 (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A2 (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_c610_A2 (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_c675_A1 (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_c670_A1 (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_c668_A2 (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_A1 (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout210_X (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c344_A3 (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_A2 (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_RESET_B (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_S0 (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_A0 (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_A4 (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_S0 (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_A4 (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c159_A3 (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout211_X (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c458_A3 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_S1 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_A0 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_A2 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_A1 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_A1 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c205_S0 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout210_A (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout212_X (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_A3 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_S0 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_A1 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_B1 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_S0 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_output116_A (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c542_SCE (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c529_A3 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_A2 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_A2 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout213_X (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c397_A1 (.DIODE(net1145));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_A2 (.DIODE(net1145));
 sky130_fd_sc_hd__diode_2 ANTENNA_c265_B1 (.DIODE(net1145));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_B1 (.DIODE(net1145));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_A1 (.DIODE(net1145));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout215_X (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_A2 (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_A3 (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c539_A3 (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c528_SCD (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c346_A0 (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_A1 (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c297_A0 (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_A3 (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_S1 (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_A4 (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout216_X (.DIODE(net1157));
 sky130_fd_sc_hd__diode_2 ANTENNA_c340_A3 (.DIODE(net1157));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_A2 (.DIODE(net1157));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_A3 (.DIODE(net1157));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_S0 (.DIODE(net1157));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_A0 (.DIODE(net1157));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_A1 (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout217_X (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_output107_A (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_A3 (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c401_A1 (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_A4 (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_S1 (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c273_B1 (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c158_A4 (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_S1 (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_A4 (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout218_X (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_A0 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c662_S1 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_S0 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c534_A1 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c409_SCD (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout219_X (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_A0 (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_A3 (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_c238_A3 (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_c228_S1 (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_S1 (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout217_A (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout218_A (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout220_X (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_c565_A0 (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_c543_A2 (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_S1 (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_A2 (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_c148_A1 (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer87_A (.DIODE(net1155));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout224_X (.DIODE(net1151));
 sky130_fd_sc_hd__diode_2 ANTENNA_c427_A3 (.DIODE(net1151));
 sky130_fd_sc_hd__diode_2 ANTENNA_c547_A1 (.DIODE(net1151));
 sky130_fd_sc_hd__diode_2 ANTENNA_c540_S0 (.DIODE(net1151));
 sky130_fd_sc_hd__diode_2 ANTENNA_c533_B1 (.DIODE(net1151));
 sky130_fd_sc_hd__diode_2 ANTENNA_c397_B1 (.DIODE(net1151));
 sky130_fd_sc_hd__diode_2 ANTENNA_c416_A0 (.DIODE(net1151));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout223_A (.DIODE(net1151));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1_A (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout225_X (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c720_A2 (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c674_SCD (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout226_X (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_A3 (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_A2 (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A1 (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_S0 (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_A0 (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_c666_SCE (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_c140_A1 (.DIODE(net1159));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone74_A4 (.DIODE(net1159));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone26_A3 (.DIODE(net1159));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout227_X (.DIODE(net1159));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_A0 (.DIODE(net1159));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_A3 (.DIODE(net1159));
 sky130_fd_sc_hd__diode_2 ANTENNA_c143_A4 (.DIODE(net1159));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_A3 (.DIODE(net1159));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone92_A (.DIODE(net1150));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer75_A (.DIODE(net1162));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout228_X (.DIODE(net1150));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_A1 (.DIODE(net1150));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_A2 (.DIODE(net1150));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_S0 (.DIODE(net1150));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout227_A (.DIODE(net1150));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout229_X (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_A0 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_A2 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c660_A4 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c532_SET_B (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_A2 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c264_A3 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_B1 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_A1 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_B1 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_A2 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout230_X (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c414_A0 (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c411_A2 (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c399_A1 (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c271_A3 (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c138_B1 (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_A0 (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_A3 (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c136_A2 (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_S0 (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_A3 (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap231_X (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_c611_S1 (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_S0 (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_S1 (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_S0 (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_c458_S1 (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold99_A (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout232_X (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_S1 (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_S1 (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_S1 (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_S1 (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_S1 (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c371_S1 (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c370_S1 (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c369_S1 (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c496_S0 (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold97_A (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout233_X (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_S1 (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_A3 (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_S1 (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_S1 (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_S1 (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_S0 (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c323_S1 (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_S0 (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_S1 (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout234_X (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c760_S0 (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_S0 (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_A3 (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_S0 (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_S0 (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_A3 (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold98_A (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout235_X (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c757_S0 (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c615_S1 (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_S1 (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_S1 (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c218_S1 (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_S1 (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c215_S1 (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_S1 (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c212_S1 (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout237_X (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA_c236_S1 (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA_c220_S1 (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA_c234_S1 (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_S1 (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_S1 (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA_c205_S1 (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout236_A (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout238_X (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_S0 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_A2 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_S1 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_A3 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_S1 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c226_S1 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c203_S1 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout237_A (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap239_X (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_A3 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_S0 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_S1 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c323_S0 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_B1 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_S1 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_S1 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap240_X (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_A2 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c321_S1 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_A0 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_S0 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_S0 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_S0 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_S1 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_A1 (.DIODE(net1152));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout241_X (.DIODE(net1152));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_A0 (.DIODE(net1152));
 sky130_fd_sc_hd__diode_2 ANTENNA_c221_A1 (.DIODE(net1152));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_A0 (.DIODE(net1152));
 sky130_fd_sc_hd__diode_2 ANTENNA_c265_A3 (.DIODE(net1152));
 sky130_fd_sc_hd__diode_2 ANTENNA_c138_A4 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout243_X (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c405_SET_B (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c404_A3 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c399_A3 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_B1 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_A1 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c269_B1 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_A3 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_A2 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_A4 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout244_X (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c111_B1 (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c278_A3 (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c264_A1 (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_A2 (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c159_A4 (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_A2 (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_A0 (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_A2 (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_A2 (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_A4 (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout245_X (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_A2 (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c124_A0 (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c120_A3 (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c115_S1 (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c114_A4 (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout246_X (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c117_A3 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_A2 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c668_A1 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c664_A1 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c663_A4 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_A2 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_S1 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c531_A2 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_A4 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_B1 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout247_X (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c763_A3 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_A2 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_A3 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_A2 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_A2 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_A3 (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c140_A4 (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout248_X (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_A1 (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_A1 (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_A1 (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c256_A3 (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_A3 (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c182_B1 (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_S1 (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_S0 (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout249_X (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c545_A1 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c538_SCE (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c530_A3 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c502_S0 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c446_A2 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c270_B1 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_S1 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_A0 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_A3 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_A1 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout250_X (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_A0 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_S0 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c691_A1 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_A3 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_A2 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout251_X (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_A2 (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_A2 (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_A2 (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_S0 (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_A1 (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_S0 (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_A3 (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_A2 (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_A1 (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_A3 (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout252_X (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c761_A1 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_A0 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c674_SET_B (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_A1 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_S1 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c272_A3 (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout253_X (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c535_A2 (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c397_A2 (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_A4 (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c276_A3 (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_A0 (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_S1 (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_A2 (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c138_A3 (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c105_S1 (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout254_X (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c762_A0 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_A3 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_S1 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_S0 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c540_A2 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout255_X (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_A2 (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_A0 (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_A1 (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_c265_A1 (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_c670_A2 (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_c560_A2 (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_c540_A3 (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_c405_SCE (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_c401_B1 (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_A3 (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout256_X (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_S0 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c203_S0 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_A0 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c119_A4 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c410_A2 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_A1 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_A2 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c286_A1 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_A1 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c136_A3 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_A1 (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout257_X (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_c676_S1 (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_A3 (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_A1 (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_c539_A4 (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_A2 (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_A0 (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_c397_A3 (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_c286_A3 (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_c267_A1 (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout258_X (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_S0 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_A1 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_S0 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c295_A1 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_A0 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c229_A2 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c205_A3 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_A4 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_A2 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_A2 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout259_X (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c702_S0 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_A3 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_A3 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c428_A1 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_A0 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_A2 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_A2 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c206_A3 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c198_A2 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c191_A2 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout262_X (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_A3 (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_A2 (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_A3 (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c671_A2 (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c537_S0 (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c536_S1 (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c535_A3 (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c531_S0 (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c528_SCE (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c408_SET_B (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone94_A (.DIODE(net1154));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer90_A (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout263_X (.DIODE(net1154));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_A0 (.DIODE(net1154));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout262_A (.DIODE(net1154));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout261_A (.DIODE(net1154));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout265_X (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_A0 (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout264_A (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c265_A4 (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c208_A3 (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c198_S1 (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout266_X (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c691_A0 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c686_A0 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c672_A4 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c671_A1 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c661_S1 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c548_S0 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c266_A1 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c182_A1 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_A2 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c136_B1 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout267_X (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c613_A2 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_A2 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c430_SCD (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_S0 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_B1 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c240_S0 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_A3 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_S1 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_S0 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_A3 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout268_X (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_A0 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_A0 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_S0 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_A1 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_A2 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout269_X (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c703_A2 (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_A1 (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c686_A1 (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_S1 (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_A3 (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c180_A1 (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_S1 (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_A2 (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_A3 (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_A3 (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout270_X (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_c237_A3 (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_c228_A3 (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_c693_A2 (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_A1 (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_c675_S1 (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_c667_A3 (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_A2 (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_c542_D (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_c274_A3 (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_c266_A3 (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout271_X (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c203_A3 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c183_A0 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_S1 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c102_A0 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_A1 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_A3 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c274_A0 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c267_A4 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_S0 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_B1 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout272_X (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c203_A0 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c662_A1 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c660_A2 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c561_A2 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c558_S0 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c541_A3 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c405_RESET_B (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_A2 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c279_A1 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_A3 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout3_A (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone13_S1 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout273_X (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_A4 (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout274_X (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_A0 (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_S0 (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_S0 (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_c106_S1 (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_A4 (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_A1 (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_A1 (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_A4 (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_A2 (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout275_X (.DIODE(net1025));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_A2 (.DIODE(net1025));
 sky130_fd_sc_hd__diode_2 ANTENNA_c695_A2 (.DIODE(net1025));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_S0 (.DIODE(net1025));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_S1 (.DIODE(net1025));
 sky130_fd_sc_hd__diode_2 ANTENNA_c366_A3 (.DIODE(net1025));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_S0 (.DIODE(net1025));
 sky130_fd_sc_hd__diode_2 ANTENNA_c276_A0 (.DIODE(net1025));
 sky130_fd_sc_hd__diode_2 ANTENNA_c221_S1 (.DIODE(net1025));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_S0 (.DIODE(net1025));
 sky130_fd_sc_hd__diode_2 ANTENNA_c100_A3 (.DIODE(net1025));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout2_A (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone13_S0 (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout276_X (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_15_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_14_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_13_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_12_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_11_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_10_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_9_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_8_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_7_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_6_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_5_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_4_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_3_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_2_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_1_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_0_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_X (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c402_CLK_N (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c405_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c406_CLK_N (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c407_CLK_N (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge806_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge814_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s905_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s909_GATE_N (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_0_0_clk_X (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_CLK_N (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c430_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge841_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s884_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s895_GATE_N (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s896_GATE_N (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s897_GATE_N (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s911_GATE_N (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_2_0_clk_X (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge840_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge845_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s908_GATE_N (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s912_GATE_N (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s914_GATE (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s915_SLEEP_B (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s918_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s919_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s920_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s936_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s943_GATE_N (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_3_0_clk_X (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c408_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c409_CLK_N (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c528_CLK_N (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c538_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c542_CLK_N (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c546_CLK_N (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c669_CLK_N (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge795_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s931_SLEEP_B (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s932_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s935_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s937_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s938_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s939_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_4_0_clk_X (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c666_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c674_CLK_N (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c678_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge803_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge813_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge816_GATE_N (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s957_GATE_N (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s958_GATE (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s959_GATE_N (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s960_GATE_N (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s961_GATE_N (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s963_SLEEP_B (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s964_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_5_0_clk_X (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge812_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge823_GATE_N (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge838_GATE (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge862_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge883_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s934_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s940_GATE_N (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s941_GATE_N (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s942_GATE (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s944_GATE_N (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s945_GATE_N (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s946_GATE (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s947_SLEEP_B (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s948_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s950_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_6_0_clk_X (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge793_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge799_CLK_N (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge815_GATE_N (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge824_GATE (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge880_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge882_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s886_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s889_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s899_SLEEP_B (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s900_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_8_0_clk_X (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge801_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge818_GATE (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge867_GATE (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge868_GATE_N (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s898_GATE (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s901_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s902_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s916_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_9_0_clk_X (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge809_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge821_GATE_N (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge822_GATE_N (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s887_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s888_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s890_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s891_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s894_GATE (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_10_0_clk_X (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge820_GATE (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge844_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge858_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge870_GATE_N (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge871_GATE (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge878_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s892_GATE_N (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s893_GATE_N (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s903_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s904_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s925_GATE_N (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_11_0_clk_X (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge850_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge860_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge866_GATE (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge872_GATE (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge874_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge875_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge876_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_13_0_clk_X (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c564_S1 (.DIODE(clknet_1_0__leaf_net714));
 sky130_fd_sc_hd__diode_2 ANTENNA_c565_S0 (.DIODE(clknet_1_0__leaf_net714));
 sky130_fd_sc_hd__diode_2 ANTENNA_c566_S0 (.DIODE(clknet_1_0__leaf_net714));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_S0 (.DIODE(clknet_1_0__leaf_net714));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_S1 (.DIODE(clknet_1_0__leaf_net714));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_A2 (.DIODE(clknet_1_0__leaf_net714));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net714_X (.DIODE(clknet_1_0__leaf_net714));
 sky130_fd_sc_hd__diode_2 ANTENNA_c415_SET_B (.DIODE(clknet_1_0__leaf_net675));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_S1 (.DIODE(clknet_1_0__leaf_net675));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_S0 (.DIODE(clknet_1_0__leaf_net675));
 sky130_fd_sc_hd__diode_2 ANTENNA_c531_S1 (.DIODE(clknet_1_0__leaf_net675));
 sky130_fd_sc_hd__diode_2 ANTENNA_c537_S1 (.DIODE(clknet_1_0__leaf_net675));
 sky130_fd_sc_hd__diode_2 ANTENNA_c667_B1 (.DIODE(clknet_1_0__leaf_net675));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net675_X (.DIODE(clknet_1_0__leaf_net675));
 sky130_fd_sc_hd__diode_2 ANTENNA_c544_B1 (.DIODE(clknet_1_0__leaf_net352));
 sky130_fd_sc_hd__diode_2 ANTENNA_c545_S0 (.DIODE(clknet_1_0__leaf_net352));
 sky130_fd_sc_hd__diode_2 ANTENNA_c546_SCE (.DIODE(clknet_1_0__leaf_net352));
 sky130_fd_sc_hd__diode_2 ANTENNA_c547_B1 (.DIODE(clknet_1_0__leaf_net352));
 sky130_fd_sc_hd__diode_2 ANTENNA_c548_A3 (.DIODE(clknet_1_0__leaf_net352));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_S0 (.DIODE(clknet_1_0__leaf_net352));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_S0 (.DIODE(clknet_1_0__leaf_net352));
 sky130_fd_sc_hd__diode_2 ANTENNA_c667_A2 (.DIODE(clknet_1_0__leaf_net352));
 sky130_fd_sc_hd__diode_2 ANTENNA_c676_A3 (.DIODE(clknet_1_0__leaf_net352));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net352_X (.DIODE(clknet_1_0__leaf_net352));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_A3 (.DIODE(clknet_1_1__leaf_net352));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_A1 (.DIODE(clknet_1_1__leaf_net352));
 sky130_fd_sc_hd__diode_2 ANTENNA_c614_A1 (.DIODE(clknet_1_1__leaf_net352));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A2 (.DIODE(clknet_1_1__leaf_net352));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_A0 (.DIODE(clknet_1_1__leaf_net352));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_A2 (.DIODE(clknet_1_1__leaf_net352));
 sky130_fd_sc_hd__diode_2 ANTENNA_c745_A3 (.DIODE(clknet_1_1__leaf_net352));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net352_X (.DIODE(clknet_1_1__leaf_net352));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_A3 (.DIODE(clknet_1_0__leaf_net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_c610_A1 (.DIODE(clknet_1_0__leaf_net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_c611_A1 (.DIODE(clknet_1_0__leaf_net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_c614_A3 (.DIODE(clknet_1_0__leaf_net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_A1 (.DIODE(clknet_1_0__leaf_net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net877_X (.DIODE(clknet_1_0__leaf_net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_A0 (.DIODE(clknet_1_1__leaf_net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_output127_A (.DIODE(clknet_1_1__leaf_net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net877_X (.DIODE(clknet_1_1__leaf_net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_c536_A2 (.DIODE(clknet_1_0__leaf_net342));
 sky130_fd_sc_hd__diode_2 ANTENNA_c537_A1 (.DIODE(clknet_1_0__leaf_net342));
 sky130_fd_sc_hd__diode_2 ANTENNA_c538_RESET_B (.DIODE(clknet_1_0__leaf_net342));
 sky130_fd_sc_hd__diode_2 ANTENNA_c539_A1 (.DIODE(clknet_1_0__leaf_net342));
 sky130_fd_sc_hd__diode_2 ANTENNA_c661_A3 (.DIODE(clknet_1_0__leaf_net342));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net342_X (.DIODE(clknet_1_0__leaf_net342));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_A1 (.DIODE(clknet_1_1__leaf_net342));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_A0 (.DIODE(clknet_1_1__leaf_net342));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_A1 (.DIODE(clknet_1_1__leaf_net342));
 sky130_fd_sc_hd__diode_2 ANTENNA_c764_A0 (.DIODE(clknet_1_1__leaf_net342));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net342_X (.DIODE(clknet_1_1__leaf_net342));
 sky130_fd_sc_hd__diode_2 ANTENNA_c757_A0 (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer4_A (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_S0 (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer3_X (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_c685_S0 (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer5_X (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_c745_A1 (.DIODE(net1033));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer8_A (.DIODE(net1033));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_A2 (.DIODE(net1033));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_A1 (.DIODE(net1033));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer7_X (.DIODE(net1033));
 sky130_fd_sc_hd__diode_2 ANTENNA_c428_A4 (.DIODE(net1039));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_A0 (.DIODE(net1039));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer12_A (.DIODE(net1039));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_A3 (.DIODE(net1039));
 sky130_fd_sc_hd__diode_2 ANTENNA_c406_RESET_B (.DIODE(net1039));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone13_X (.DIODE(net1039));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer15_A (.DIODE(net1040));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_A2 (.DIODE(net1040));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer14_X (.DIODE(net1040));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_A2 (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_c558_A1 (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer15_X (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer19_A (.DIODE(net1043));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer18_A (.DIODE(net1043));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_A3 (.DIODE(net1043));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer17_X (.DIODE(net1043));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_A0 (.DIODE(net1050));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_A1 (.DIODE(net1050));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer24_X (.DIODE(net1050));
 sky130_fd_sc_hd__diode_2 ANTENNA_c271_A4 (.DIODE(net1052));
 sky130_fd_sc_hd__diode_2 ANTENNA_c541_A0 (.DIODE(net1052));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone13_A2 (.DIODE(net1052));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer25_A (.DIODE(net1052));
 sky130_fd_sc_hd__diode_2 ANTENNA_c532_RESET_B (.DIODE(net1052));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone26_X (.DIODE(net1052));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer30_A (.DIODE(net1055));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_A1 (.DIODE(net1055));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer29_X (.DIODE(net1055));
 sky130_fd_sc_hd__diode_2 ANTENNA_c613_A0 (.DIODE(net1057));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_A2 (.DIODE(net1057));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer31_X (.DIODE(net1057));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout206_A (.DIODE(net1059));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer33_X (.DIODE(net1059));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_A1 (.DIODE(net1060));
 sky130_fd_sc_hd__diode_2 ANTENNA_c739_A3 (.DIODE(net1060));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_A0 (.DIODE(net1060));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer35_A (.DIODE(net1060));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer34_X (.DIODE(net1060));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout209_A (.DIODE(net1064));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer38_X (.DIODE(net1064));
 sky130_fd_sc_hd__diode_2 ANTENNA_c563_A1 (.DIODE(net1068));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer43_A (.DIODE(net1068));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_A0 (.DIODE(net1068));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_S0 (.DIODE(net1068));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer42_X (.DIODE(net1068));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer53_A (.DIODE(net1077));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_A1 (.DIODE(net1077));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer52_A (.DIODE(net1077));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_A2 (.DIODE(net1077));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer51_X (.DIODE(net1077));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_A1 (.DIODE(net1080));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer54_X (.DIODE(net1080));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone26_A0 (.DIODE(net1081));
 sky130_fd_sc_hd__diode_2 ANTENNA_c269_A2 (.DIODE(net1081));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_A3 (.DIODE(net1081));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_A0 (.DIODE(net1081));
 sky130_fd_sc_hd__diode_2 ANTENNA_c212_A3 (.DIODE(net1081));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone55_X (.DIODE(net1081));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer57_A (.DIODE(net1082));
 sky130_fd_sc_hd__diode_2 ANTENNA_c665_A3 (.DIODE(net1082));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer56_X (.DIODE(net1082));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_S0 (.DIODE(net1085));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_A2 (.DIODE(net1085));
 sky130_fd_sc_hd__diode_2 ANTENNA_c286_S0 (.DIODE(net1085));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_S0 (.DIODE(net1085));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_A2 (.DIODE(net1085));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone59_X (.DIODE(net1085));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_A2 (.DIODE(net1086));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_A3 (.DIODE(net1086));
 sky130_fd_sc_hd__diode_2 ANTENNA_c528_D (.DIODE(net1086));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_A3 (.DIODE(net1086));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_A2 (.DIODE(net1086));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone60_X (.DIODE(net1086));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_A1 (.DIODE(net1087));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer62_A (.DIODE(net1087));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_A3 (.DIODE(net1087));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer61_X (.DIODE(net1087));
 sky130_fd_sc_hd__diode_2 ANTENNA_c536_S0 (.DIODE(net1098));
 sky130_fd_sc_hd__diode_2 ANTENNA_c537_A3 (.DIODE(net1098));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_B1 (.DIODE(net1098));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_A2 (.DIODE(net1098));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_A2 (.DIODE(net1098));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone72_X (.DIODE(net1098));
 sky130_fd_sc_hd__diode_2 ANTENNA_c723_A3 (.DIODE(net1101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c747_S0 (.DIODE(net1101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_A3 (.DIODE(net1101));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer75_X (.DIODE(net1101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_A0 (.DIODE(net1104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c446_A3 (.DIODE(net1104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c372_A1 (.DIODE(net1104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_A1 (.DIODE(net1104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_S1 (.DIODE(net1104));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone78_X (.DIODE(net1104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_A2 (.DIODE(net1105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c406_SCE (.DIODE(net1105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c222_A2 (.DIODE(net1105));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer76_A (.DIODE(net1105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_S0 (.DIODE(net1105));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone79_X (.DIODE(net1105));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer81_A (.DIODE(net1106));
 sky130_fd_sc_hd__diode_2 ANTENNA_output172_A (.DIODE(net1106));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer80_X (.DIODE(net1106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_S0 (.DIODE(net1108));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_A1 (.DIODE(net1108));
 sky130_fd_sc_hd__diode_2 ANTENNA_c762_A2 (.DIODE(net1108));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_A3 (.DIODE(net1108));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_A3 (.DIODE(net1108));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone82_X (.DIODE(net1108));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_A2 (.DIODE(net1109));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer84_A (.DIODE(net1109));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer83_X (.DIODE(net1109));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_S1 (.DIODE(net1112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_A1 (.DIODE(net1112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_A1 (.DIODE(net1112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_A3 (.DIODE(net1112));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer85_A (.DIODE(net1112));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone86_X (.DIODE(net1112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_A1 (.DIODE(net1113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_A2 (.DIODE(net1113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_S0 (.DIODE(net1113));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer87_X (.DIODE(net1113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_A3 (.DIODE(net1114));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_A3 (.DIODE(net1114));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_A1 (.DIODE(net1114));
 sky130_fd_sc_hd__diode_2 ANTENNA_output148_A (.DIODE(net1114));
 sky130_fd_sc_hd__diode_2 ANTENNA_c184_A2 (.DIODE(net1114));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone88_X (.DIODE(net1114));
 sky130_fd_sc_hd__diode_2 ANTENNA_c346_A3 (.DIODE(net1115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c230_A1 (.DIODE(net1115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c229_S0 (.DIODE(net1115));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer89_X (.DIODE(net1115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c543_A3 (.DIODE(net1118));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone13_A0 (.DIODE(net1118));
 sky130_fd_sc_hd__diode_2 ANTENNA_c665_A2 (.DIODE(net1118));
 sky130_fd_sc_hd__diode_2 ANTENNA_output101_A (.DIODE(net1118));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_A3 (.DIODE(net1118));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_A1 (.DIODE(net1118));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone92_X (.DIODE(net1118));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_S1 (.DIODE(net1120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_S0 (.DIODE(net1120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c402_SCE (.DIODE(net1120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_S1 (.DIODE(net1120));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone94_X (.DIODE(net1120));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1_X (.DIODE(net1161));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone26_A2 (.DIODE(net1153));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone13_A3 (.DIODE(net1153));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_A3 (.DIODE(net1153));
 sky130_fd_sc_hd__diode_2 ANTENNA_c529_A4 (.DIODE(net1153));
 sky130_fd_sc_hd__diode_2 ANTENNA_c430_D (.DIODE(net1153));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_A1 (.DIODE(net1153));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_A3 (.DIODE(net1153));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_A2 (.DIODE(net1153));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_A3 (.DIODE(net1153));
 sky130_fd_sc_hd__diode_2 ANTENNA_c140_A3 (.DIODE(net1153));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout2_X (.DIODE(net1133));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_A1 (.DIODE(net1133));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_A3 (.DIODE(net1133));
 sky130_fd_sc_hd__diode_2 ANTENNA_c661_A2 (.DIODE(net1133));
 sky130_fd_sc_hd__diode_2 ANTENNA_c547_A2 (.DIODE(net1133));
 sky130_fd_sc_hd__diode_2 ANTENNA_c533_A1 (.DIODE(net1133));
 sky130_fd_sc_hd__diode_2 ANTENNA_c437_A1 (.DIODE(net1133));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_A2 (.DIODE(net1133));
 sky130_fd_sc_hd__diode_2 ANTENNA_c190_A3 (.DIODE(net1133));
 sky130_fd_sc_hd__diode_2 ANTENNA_c180_B1 (.DIODE(net1133));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_S0 (.DIODE(net1133));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout4_X (.DIODE(net1135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_A0 (.DIODE(net1135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_A3 (.DIODE(net1135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_A1 (.DIODE(net1135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c286_S1 (.DIODE(net1135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c159_A2 (.DIODE(net1135));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone13_A1 (.DIODE(net1135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c413_S0 (.DIODE(net1135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_A1 (.DIODE(net1135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c134_A3 (.DIODE(net1135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_A2 (.DIODE(net1135));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer13 (.A(net45),
    .X(net1136));
 sky130_fd_sc_hd__mux4_1 clone14 (.A0(net22),
    .A1(net753),
    .A2(net993),
    .A3(net1160),
    .S0(net1148),
    .S1(net972),
    .X(net1137));
 sky130_fd_sc_hd__a41o_1 clone15 (.A1(net26),
    .A2(net18),
    .A3(net993),
    .A4(net1121),
    .B1(net25),
    .X(net1138));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer26 (.A(net295),
    .X(net1139));
 sky130_fd_sc_hd__mux4_1 clone27 (.A0(net823),
    .A1(net237),
    .A2(net958),
    .A3(net635),
    .S0(net668),
    .S1(net687),
    .X(net1140));
 sky130_fd_sc_hd__a41o_1 clone28 (.A1(net991),
    .A2(net994),
    .A3(net756),
    .A4(net1024),
    .B1(net996),
    .X(net1141));
 sky130_fd_sc_hd__a41o_1 clone29 (.A1(net998),
    .A2(net1024),
    .A3(net1007),
    .A4(net994),
    .B1(net1011),
    .X(net1142));
 sky130_fd_sc_hd__a41o_1 clone30 (.A1(net128),
    .A2(net944),
    .A3(net994),
    .A4(net125),
    .B1(net949),
    .X(net1143));
 sky130_fd_sc_hd__mux4_1 clone31 (.A0(net954),
    .A1(net911),
    .A2(net953),
    .A3(net753),
    .S0(net966),
    .S1(net1003),
    .X(net1144));
 sky130_fd_sc_hd__clkbuf_1 clone32 (.A(net30),
    .X(net1145));
 sky130_fd_sc_hd__clkbuf_1 clone33 (.A(net31),
    .X(net1146));
 sky130_fd_sc_hd__clkbuf_1 clone34 (.A(net32),
    .X(net1147));
 sky130_fd_sc_hd__a41o_1 clone35 (.A1(net991),
    .A2(net994),
    .A3(net756),
    .A4(net1024),
    .B1(net996),
    .X(net1148));
 sky130_fd_sc_hd__clkbuf_1 clone36 (.A(net123),
    .X(net1149));
 sky130_fd_sc_hd__clkbuf_1 clone37 (.A(net851),
    .X(net1150));
 sky130_fd_sc_hd__clkbuf_1 clone38 (.A(net21),
    .X(net1151));
 sky130_fd_sc_hd__clkbuf_1 clone39 (.A(net922),
    .X(net1152));
 sky130_fd_sc_hd__clkbuf_1 clone40 (.A(net975),
    .X(net1153));
 sky130_fd_sc_hd__clkbuf_1 clone41 (.A(net774),
    .X(net1154));
 sky130_fd_sc_hd__clkbuf_1 clone42 (.A(net21),
    .X(net1155));
 sky130_fd_sc_hd__a41o_1 clone43 (.A1(net1161),
    .A2(net1011),
    .A3(net1160),
    .A4(net998),
    .B1(net18),
    .X(net1156));
 sky130_fd_sc_hd__clkbuf_1 clone44 (.A(net27),
    .X(net1157));
 sky130_fd_sc_hd__clkbuf_1 clone45 (.A(net947),
    .X(net1158));
 sky130_fd_sc_hd__clkbuf_1 clone46 (.A(net1162),
    .X(net1159));
 sky130_fd_sc_hd__clkbuf_1 clone47 (.A(net978),
    .X(net1160));
 sky130_fd_sc_hd__clkbuf_1 clone48 (.A(net975),
    .X(net1161));
 sky130_fd_sc_hd__clkbuf_1 clone49 (.A(net851),
    .X(net1162));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_186 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_282 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_440 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_283 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_400 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_412 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_198 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_340 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_451 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_168 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_168 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_114 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_191 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_17 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_171 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_478 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_114 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_351 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_442 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_469 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_242 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_412 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_13 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_31 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_357 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_488 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_102 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_339 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_88 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_254 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_283 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_118 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_256 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_84 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_60 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_392 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_412 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_339 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_8 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_20 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_271 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_115 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_311 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_450 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_544 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_95 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_144 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_219 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_336 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_47 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_219 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_423 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_242 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_13 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_423 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_400 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_507 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_368 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_87 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_128 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_143 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_490 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_476 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_10 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_5 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_310 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_479 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_24 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_451 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_107 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_14 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_379 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_87 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_135 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_303 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_227 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_282 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_123 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_135 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_58 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_5 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_12 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_133 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_214 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_617 ();
endmodule
