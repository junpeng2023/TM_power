module netlist_0 (clk,
    in0,
    in1,
    in10,
    in11,
    in12,
    in13,
    in14,
    in15,
    in16,
    in17,
    in18,
    in19,
    in2,
    in20,
    in21,
    in22,
    in23,
    in24,
    in3,
    in4,
    in5,
    in6,
    in7,
    in8,
    in9,
    out0,
    out1,
    out10,
    out11,
    out12,
    out13,
    out14,
    out15,
    out16,
    out17,
    out18,
    out19,
    out2,
    out20,
    out21,
    out22,
    out23,
    out24,
    out3,
    out4,
    out5,
    out6,
    out7,
    out8,
    out9,
    rst);
 input clk;
 input in0;
 input in1;
 input in10;
 input in11;
 input in12;
 input in13;
 input in14;
 input in15;
 input in16;
 input in17;
 input in18;
 input in19;
 input in2;
 input in20;
 input in21;
 input in22;
 input in23;
 input in24;
 input in3;
 input in4;
 input in5;
 input in6;
 input in7;
 input in8;
 input in9;
 output out0;
 output out1;
 output out10;
 output out11;
 output out12;
 output out13;
 output out14;
 output out15;
 output out16;
 output out17;
 output out18;
 output out19;
 output out2;
 output out20;
 output out21;
 output out22;
 output out23;
 output out24;
 output out3;
 output out4;
 output out5;
 output out6;
 output out7;
 output out8;
 output out9;
 input rst;

 wire net0;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net63;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net64;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net65;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net66;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net67;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net68;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net69;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net7;
 wire net70;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net71;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net72;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net73;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net74;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net747;
 wire net748;
 wire net749;
 wire net75;
 wire net750;
 wire net751;
 wire net752;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net76;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net77;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net78;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net79;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net746;
 wire net753;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire clknet_leaf_0_clk;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire clknet_0_net721;
 wire clknet_1_0__leaf_net721;
 wire clknet_1_1__leaf_net721;
 wire clknet_0_net730;
 wire clknet_1_0__leaf_net730;
 wire clknet_1_1__leaf_net730;
 wire clknet_0_net733;
 wire clknet_1_0__leaf_net733;
 wire clknet_1_1__leaf_net733;
 wire clknet_0_net794;
 wire clknet_1_0__leaf_net794;
 wire clknet_1_1__leaf_net794;
 wire clknet_0_net714;
 wire clknet_1_0__leaf_net714;
 wire clknet_1_1__leaf_net714;
 wire clknet_0_net779;
 wire clknet_1_0__leaf_net779;
 wire clknet_1_1__leaf_net779;
 wire clknet_0_net278;
 wire clknet_1_0__leaf_net278;
 wire clknet_1_1__leaf_net278;
 wire clknet_0_net285;
 wire clknet_1_0__leaf_net285;
 wire clknet_1_1__leaf_net285;
 wire clknet_0_net284;
 wire clknet_1_0__leaf_net284;
 wire clknet_1_1__leaf_net284;
 wire clknet_0_net287;
 wire clknet_1_0__leaf_net287;
 wire clknet_1_1__leaf_net287;
 wire clknet_0_net248;
 wire clknet_1_0__leaf_net248;
 wire clknet_1_1__leaf_net248;
 wire clknet_0_net255;
 wire clknet_1_0__leaf_net255;
 wire clknet_1_1__leaf_net255;
 wire clknet_0_net256;
 wire clknet_1_0__leaf_net256;
 wire clknet_1_1__leaf_net256;
 wire clknet_0_net520;
 wire clknet_1_0__leaf_net520;
 wire clknet_1_1__leaf_net520;
 wire clknet_0_net523;
 wire clknet_1_0__leaf_net523;
 wire clknet_1_1__leaf_net523;
 wire clknet_0_net525;
 wire clknet_1_0__leaf_net525;
 wire clknet_1_1__leaf_net525;
 wire clknet_0_net530;
 wire clknet_1_0__leaf_net530;
 wire clknet_1_1__leaf_net530;
 wire clknet_0_net527;
 wire clknet_1_0__leaf_net527;
 wire clknet_1_1__leaf_net527;
 wire clknet_0_net521;
 wire clknet_1_0__leaf_net521;
 wire clknet_1_1__leaf_net521;
 wire clknet_0_net640;
 wire clknet_1_0__leaf_net640;
 wire clknet_1_1__leaf_net640;
 wire clknet_0_net566;
 wire clknet_1_0__leaf_net566;
 wire clknet_1_1__leaf_net566;
 wire clknet_0_net524;
 wire clknet_1_0__leaf_net524;
 wire clknet_1_1__leaf_net524;
 wire clknet_0_net251;
 wire clknet_1_0__leaf_net251;
 wire clknet_1_1__leaf_net251;
 wire clknet_0_net264;
 wire clknet_1_0__leaf_net264;
 wire clknet_1_1__leaf_net264;
 wire clknet_0_net252;
 wire clknet_1_0__leaf_net252;
 wire clknet_1_1__leaf_net252;
 wire clknet_0_net761;
 wire clknet_1_0__leaf_net761;
 wire clknet_1_1__leaf_net761;
 wire clknet_0_net96;
 wire clknet_1_0__leaf_net96;
 wire clknet_1_1__leaf_net96;
 wire clknet_0_net95;
 wire clknet_1_0__leaf_net95;
 wire clknet_1_1__leaf_net95;
 wire clknet_0_net97;
 wire clknet_1_0__leaf_net97;
 wire clknet_1_1__leaf_net97;
 wire clknet_0_net724;
 wire clknet_1_0__leaf_net724;
 wire clknet_1_1__leaf_net724;
 wire clknet_0_net725;
 wire clknet_1_0__leaf_net725;
 wire clknet_1_1__leaf_net725;
 wire clknet_0_net727;
 wire clknet_1_0__leaf_net727;
 wire clknet_1_1__leaf_net727;
 wire clknet_0_net726;
 wire clknet_1_0__leaf_net726;
 wire clknet_1_1__leaf_net726;
 wire clknet_0_net709;
 wire clknet_1_0__leaf_net709;
 wire clknet_1_1__leaf_net709;
 wire clknet_0_net710;
 wire clknet_1_0__leaf_net710;
 wire clknet_1_1__leaf_net710;
 wire clknet_0_net519;
 wire clknet_1_0__leaf_net519;
 wire clknet_1_1__leaf_net519;
 wire clknet_0_net518;
 wire clknet_1_0__leaf_net518;
 wire clknet_1_1__leaf_net518;
 wire clknet_0_net308;
 wire clknet_1_0__leaf_net308;
 wire clknet_1_1__leaf_net308;
 wire clknet_0_net306;
 wire clknet_1_0__leaf_net306;
 wire clknet_1_1__leaf_net306;
 wire clknet_0_net318;
 wire clknet_1_0__leaf_net318;
 wire clknet_1_1__leaf_net318;
 wire clknet_0_net303;
 wire clknet_1_0__leaf_net303;
 wire clknet_1_1__leaf_net303;
 wire clknet_0_net190;
 wire clknet_1_0__leaf_net190;
 wire clknet_1_1__leaf_net190;
 wire clknet_0_net187;
 wire clknet_1_0__leaf_net187;
 wire clknet_1_1__leaf_net187;
 wire clknet_0_net188;
 wire clknet_1_0__leaf_net188;
 wire clknet_1_1__leaf_net188;
 wire clknet_0_net183;
 wire clknet_1_0__leaf_net183;
 wire clknet_1_1__leaf_net183;
 wire clknet_0_net191;
 wire clknet_1_0__leaf_net191;
 wire clknet_1_1__leaf_net191;
 wire clknet_0_net194;
 wire clknet_1_0__leaf_net194;
 wire clknet_1_1__leaf_net194;
 wire clknet_0_net321;
 wire clknet_1_0__leaf_net321;
 wire clknet_1_1__leaf_net321;
 wire clknet_0_net319;
 wire clknet_1_0__leaf_net319;
 wire clknet_1_1__leaf_net319;
 wire clknet_0_net186;
 wire clknet_1_0__leaf_net186;
 wire clknet_1_1__leaf_net186;
 wire clknet_0_net185;
 wire clknet_1_0__leaf_net185;
 wire clknet_1_1__leaf_net185;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;

 sky130_fd_sc_hd__and3_1 c100 (.A(net79),
    .B(net78),
    .C(net84),
    .X(net85));
 sky130_fd_sc_hd__and3_1 c101 (.A(net67),
    .B(net79),
    .C(net75),
    .X(net86));
 sky130_fd_sc_hd__and3_1 c102 (.A(net86),
    .B(net84),
    .C(net80),
    .X(net87));
 sky130_fd_sc_hd__sdfrbp_1 c103 (.CLK(clknet_leaf_32_clk),
    .D(net85),
    .RESET_B(net72),
    .SCD(net87),
    .SCE(net82),
    .Q(net88));
 sky130_fd_sc_hd__sdfxbp_1 c104 (.CLK(clknet_leaf_32_clk),
    .D(net75),
    .SCD(net87),
    .SCE(net959),
    .Q(net90),
    .Q_N(net89));
 sky130_fd_sc_hd__clkbuf_1 c105 (.A(net90),
    .X(net91));
 sky130_fd_sc_hd__clkbuf_1 c106 (.A(net59),
    .X(net92));
 sky130_fd_sc_hd__clkbuf_2 c107 (.A(net91),
    .X(net93));
 sky130_fd_sc_hd__and2_0 c108 (.A(net93),
    .B(net92),
    .X(net94));
 sky130_fd_sc_hd__buf_1 c109 (.A(clknet_1_0__leaf_net761),
    .X(net95));
 sky130_fd_sc_hd__buf_1 c110 (.A(clknet_1_1__leaf_net761),
    .X(net96));
 sky130_fd_sc_hd__and2_0 c111 (.A(clknet_1_0__leaf_net95),
    .B(net93),
    .X(net97));
 sky130_fd_sc_hd__and2_2 c112 (.A(net91),
    .B(net93),
    .X(net98));
 sky130_fd_sc_hd__and2_0 c113 (.A(net92),
    .B(clknet_1_1__leaf_net95),
    .X(net99));
 sky130_fd_sc_hd__dfstp_1 c114 (.CLK(clknet_leaf_32_clk),
    .D(net93),
    .SET_B(net908),
    .Q(net100));
 sky130_fd_sc_hd__sdfxbp_1 c115 (.CLK(clknet_leaf_33_clk),
    .D(clknet_1_0__leaf_net97),
    .SCD(net98),
    .SCE(clknet_1_0__leaf_net95),
    .Q(net101));
 sky130_fd_sc_hd__sdfxtp_1 c116 (.CLK(clknet_leaf_32_clk),
    .D(net98),
    .SCD(clknet_1_0__leaf_net96),
    .SCE(clknet_1_1__leaf_net95),
    .Q(net102));
 sky130_fd_sc_hd__and2_0 c117 (.A(net102),
    .B(net90),
    .X(net103));
 sky130_fd_sc_hd__dfstp_1 c118 (.CLK(clknet_leaf_32_clk),
    .D(net864),
    .SET_B(clknet_1_1__leaf_net97),
    .Q(net104));
 sky130_fd_sc_hd__dlrbn_1 c119 (.D(net99),
    .GATE_N(clknet_leaf_32_clk),
    .RESET_B(net950),
    .Q(net105));
 sky130_fd_sc_hd__and2_0 c120 (.A(net103),
    .B(net104),
    .X(net106));
 sky130_fd_sc_hd__or4bb_1 c121 (.A(net100),
    .B(net106),
    .C_N(net104),
    .D_N(net93),
    .X(net107));
 sky130_fd_sc_hd__sdfxtp_1 c122 (.CLK(clknet_leaf_32_clk),
    .D(clknet_1_1__leaf_net96),
    .SCD(net104),
    .SCE(net107),
    .Q(net108));
 sky130_fd_sc_hd__sdfxtp_1 c123 (.CLK(clknet_leaf_32_clk),
    .D(net106),
    .SCD(net107),
    .SCE(net980),
    .Q(net109));
 sky130_fd_sc_hd__mux4_1 c124 (.A0(net105),
    .A1(net108),
    .A2(net109),
    .A3(net104),
    .S0(net98),
    .S1(net93),
    .X(net110));
 sky130_fd_sc_hd__dfbbn_1 c125 (.CLK_N(clknet_leaf_27_clk),
    .D(net109),
    .RESET_B(net908),
    .SET_B(net778),
    .Q(net111));
 sky130_fd_sc_hd__and2_0 c126 (.A(net753),
    .B(net806),
    .X(net112));
 sky130_fd_sc_hd__and2_0 c127 (.A(net112),
    .B(net819),
    .X(net113));
 sky130_fd_sc_hd__and2_0 c128 (.A(net113),
    .B(net801),
    .X(net114));
 sky130_fd_sc_hd__and2_2 c129 (.A(net800),
    .B(net799),
    .X(net115));
 sky130_fd_sc_hd__and2_0 c130 (.A(net115),
    .B(net815),
    .X(net116));
 sky130_fd_sc_hd__and2_1 c131 (.A(net802),
    .B(net115),
    .X(net117));
 sky130_fd_sc_hd__and2_0 c132 (.A(net116),
    .B(net808),
    .X(net118));
 sky130_fd_sc_hd__and2_0 c133 (.A(net813),
    .B(net117),
    .X(net119));
 sky130_fd_sc_hd__dlrbn_1 c134 (.D(net119),
    .GATE_N(clknet_leaf_4_clk),
    .RESET_B(net115),
    .Q(net120));
 sky130_fd_sc_hd__and2_0 c135 (.A(net115),
    .B(net746),
    .X(net121));
 sky130_fd_sc_hd__and2_1 c136 (.A(net117),
    .B(net805),
    .X(net122));
 sky130_fd_sc_hd__dlrbp_1 c137 (.D(net114),
    .GATE(clknet_leaf_4_clk),
    .RESET_B(net122),
    .Q(net123));
 sky130_fd_sc_hd__dlrbp_1 c138 (.D(net865),
    .GATE(clknet_leaf_4_clk),
    .RESET_B(net122),
    .Q(net125),
    .Q_N(net124));
 sky130_fd_sc_hd__dlrtn_1 c139 (.D(net122),
    .GATE_N(clknet_leaf_4_clk),
    .RESET_B(net862),
    .Q(net126));
 sky130_fd_sc_hd__and3_2 c140 (.A(net126),
    .B(net124),
    .C(net115),
    .X(net127));
 sky130_fd_sc_hd__and3_1 c141 (.A(net964),
    .B(net903),
    .C(net117),
    .X(net128));
 sky130_fd_sc_hd__dfbbn_1 c142 (.CLK_N(clknet_leaf_4_clk),
    .D(net121),
    .RESET_B(net122),
    .SET_B(net124),
    .Q(net130),
    .Q_N(net129));
 sky130_fd_sc_hd__dfbbp_1 c143 (.CLK(clknet_leaf_4_clk),
    .D(net862),
    .RESET_B(net128),
    .SET_B(net130),
    .Q(net131));
 sky130_fd_sc_hd__sdfbbp_1 c144 (.CLK(clknet_leaf_4_clk),
    .D(net118),
    .RESET_B(net130),
    .SCD(net127),
    .SCE(net128),
    .SET_B(net115),
    .Q(net132));
 sky130_fd_sc_hd__a2111o_1 c145 (.A1(net131),
    .A2(net117),
    .B1(net129),
    .C1(net124),
    .D1(net115),
    .X(net133));
 sky130_fd_sc_hd__mux4_1 c146 (.A0(net132),
    .A1(net133),
    .A2(net122),
    .A3(net129),
    .S0(net115),
    .S1(net127),
    .X(net134));
 sky130_fd_sc_hd__buf_1 c147 (.A(net127),
    .X(net135));
 sky130_fd_sc_hd__buf_1 c148 (.A(net747),
    .X(net136));
 sky130_fd_sc_hd__clkbuf_1 c149 (.A(net136),
    .X(net137));
 sky130_fd_sc_hd__dlrtn_1 c150 (.D(net18),
    .GATE_N(clknet_leaf_3_clk),
    .RESET_B(net135),
    .Q(net138));
 sky130_fd_sc_hd__buf_1 c151 (.A(net747),
    .X(net139));
 sky130_fd_sc_hd__dlrtn_1 c152 (.D(net135),
    .GATE_N(clknet_leaf_3_clk),
    .RESET_B(net893),
    .Q(net140));
 sky130_fd_sc_hd__and3_1 c153 (.A(net975),
    .B(net818),
    .C(net139),
    .X(net141));
 sky130_fd_sc_hd__and2_0 c154 (.A(net139),
    .B(net16),
    .X(net142));
 sky130_fd_sc_hd__and2_0 c155 (.A(net136),
    .B(net139),
    .X(net143));
 sky130_fd_sc_hd__and2_2 c156 (.A(net143),
    .B(net139),
    .X(net144));
 sky130_fd_sc_hd__and2_1 c157 (.A(net2),
    .B(net143),
    .X(net145));
 sky130_fd_sc_hd__dlrtp_1 c158 (.D(net142),
    .GATE(clknet_leaf_3_clk),
    .RESET_B(net145),
    .Q(net146));
 sky130_fd_sc_hd__and3_1 c159 (.A(net141),
    .B(net146),
    .C(net145),
    .X(net147));
 sky130_fd_sc_hd__and2_1 c160 (.A(net145),
    .B(net146),
    .X(net148));
 sky130_fd_sc_hd__dlrtp_1 c161 (.D(net147),
    .GATE(clknet_leaf_3_clk),
    .RESET_B(net148),
    .Q(net149));
 sky130_fd_sc_hd__mux4_1 c162 (.A0(net140),
    .A1(net148),
    .A2(net145),
    .A3(net144),
    .S0(net146),
    .S1(clknet_1_0__leaf_net779),
    .X(net150));
 sky130_fd_sc_hd__and3_1 c163 (.A(net136),
    .B(net145),
    .C(net144),
    .X(net151));
 sky130_fd_sc_hd__and2_0 c164 (.A(net149),
    .B(net780),
    .X(net152));
 sky130_fd_sc_hd__dlrtp_1 c165 (.D(net148),
    .GATE(clknet_leaf_3_clk),
    .RESET_B(net152),
    .Q(net153));
 sky130_fd_sc_hd__and2_0 c166 (.A(net137),
    .B(net153),
    .X(net154));
 sky130_fd_sc_hd__and2_0 c167 (.A(net154),
    .B(net146),
    .X(net155));
 sky130_fd_sc_hd__buf_1 c168 (.A(net30),
    .X(net156));
 sky130_fd_sc_hd__buf_1 c169 (.A(net156),
    .X(net157));
 sky130_fd_sc_hd__and2_0 c170 (.A(net156),
    .B(net157),
    .X(net158));
 sky130_fd_sc_hd__buf_1 c171 (.A(net157),
    .X(net159));
 sky130_fd_sc_hd__buf_1 c172 (.A(net156),
    .X(net160));
 sky130_fd_sc_hd__dlymetal6s2s_1 c173 (.A(net156),
    .X(net161));
 sky130_fd_sc_hd__buf_1 c174 (.A(net760),
    .X(net162));
 sky130_fd_sc_hd__and2_1 c175 (.A(net161),
    .B(net162),
    .X(net163));
 sky130_fd_sc_hd__sdfxbp_1 c176 (.CLK(clknet_leaf_37_clk),
    .D(net157),
    .SCD(net163),
    .SCE(net161),
    .Q(net164));
 sky130_fd_sc_hd__and2_2 c177 (.A(net161),
    .B(net162),
    .X(net165));
 sky130_fd_sc_hd__sdfrtn_1 c178 (.CLK_N(clknet_leaf_0_clk),
    .D(net157),
    .RESET_B(net165),
    .SCD(net162),
    .SCE(net163),
    .Q(net166));
 sky130_fd_sc_hd__sdfrtp_2 c179 (.CLK(clknet_leaf_37_clk),
    .D(net163),
    .RESET_B(net161),
    .SCD(net144),
    .SCE(net165),
    .Q(net167));
 sky130_fd_sc_hd__and2_0 c180 (.A(net160),
    .B(net167),
    .X(net168));
 sky130_fd_sc_hd__sdfxbp_1 c181 (.CLK(clknet_leaf_37_clk),
    .D(net887),
    .SCD(net165),
    .SCE(net161),
    .Q(net170),
    .Q_N(net169));
 sky130_fd_sc_hd__sdfxtp_1 c182 (.CLK(clknet_leaf_0_clk),
    .D(net162),
    .SCD(net165),
    .SCE(net860),
    .Q(net171));
 sky130_fd_sc_hd__and2_0 c183 (.A(net166),
    .B(net171),
    .X(net172));
 sky130_fd_sc_hd__sdfxtp_1 c184 (.CLK(clknet_leaf_37_clk),
    .D(net158),
    .SCD(net159),
    .SCE(net927),
    .Q(net173));
 sky130_fd_sc_hd__clkbuf_1 c185 (.A(net760),
    .X(net174));
 sky130_fd_sc_hd__sdfrtp_1 c186 (.CLK(clknet_leaf_0_clk),
    .D(net165),
    .RESET_B(net844),
    .SCD(net174),
    .SCE(net159),
    .Q(net175));
 sky130_fd_sc_hd__and3_1 c187 (.A(net175),
    .B(net160),
    .C(net173),
    .X(net176));
 sky130_fd_sc_hd__mux4_1 c188 (.A0(net174),
    .A1(net176),
    .A2(net171),
    .A3(net173),
    .S0(net165),
    .S1(net167),
    .X(net177));
 sky130_fd_sc_hd__and2_1 c189 (.A(net170),
    .B(net167),
    .X(net178));
 sky130_fd_sc_hd__and2_1 c190 (.A(net178),
    .B(net48),
    .X(net179));
 sky130_fd_sc_hd__edfxbp_1 c191 (.CLK(clknet_leaf_0_clk),
    .D(net178),
    .DE(net179),
    .Q(net181),
    .Q_N(net180));
 sky130_fd_sc_hd__edfxtp_1 c192 (.CLK(clknet_leaf_30_clk),
    .D(net179),
    .DE(net958),
    .Q(net182));
 sky130_fd_sc_hd__sdlclkp_1 c193 (.CLK(clknet_leaf_0_clk),
    .GATE(net178),
    .SCE(net179),
    .GCLK(net183));
 sky130_fd_sc_hd__and2_0 c194 (.A(net182),
    .B(net178),
    .X(net184));
 sky130_fd_sc_hd__and2_0 c195 (.A(net184),
    .B(clknet_1_0__leaf_net183),
    .X(net185));
 sky130_fd_sc_hd__and2_0 c196 (.A(net184),
    .B(clknet_1_0__leaf_net183),
    .X(net186));
 sky130_fd_sc_hd__sdlclkp_2 c197 (.CLK(clknet_leaf_30_clk),
    .GATE(clknet_1_0__leaf_net185),
    .SCE(clknet_1_0__leaf_net186),
    .GCLK(net187));
 sky130_fd_sc_hd__and3_1 c198 (.A(clknet_1_0__leaf_net183),
    .B(net184),
    .C(clknet_1_1__leaf_net187),
    .X(net188));
 sky130_fd_sc_hd__and2_0 c199 (.A(clknet_1_0__leaf_net187),
    .B(net180),
    .X(net189));
 sky130_fd_sc_hd__sdlclkp_4 c200 (.CLK(clknet_leaf_29_clk),
    .GATE(clknet_1_0__leaf_net188),
    .SCE(clknet_1_1__leaf_net185),
    .GCLK(net190));
 sky130_fd_sc_hd__and2_0 c201 (.A(net958),
    .B(clknet_1_1__leaf_net183),
    .X(net191));
 sky130_fd_sc_hd__sdfbbn_1 c202 (.CLK_N(clknet_leaf_30_clk),
    .D(clknet_1_1__leaf_net190),
    .RESET_B(clknet_1_0__leaf_net188),
    .SCD(clknet_1_0__leaf_net191),
    .SCE(net178),
    .SET_B(clknet_1_1__leaf_net187),
    .Q(net193),
    .Q_N(net192));
 sky130_fd_sc_hd__and2_0 c203 (.A(clknet_1_1__leaf_net191),
    .B(net193),
    .X(net194));
 sky130_fd_sc_hd__or4bb_1 c204 (.A(clknet_1_0__leaf_net187),
    .B(net192),
    .C_N(clknet_1_0__leaf_net183),
    .D_N(net866),
    .X(net195));
 sky130_fd_sc_hd__sdfxtp_1 c205 (.CLK(clknet_leaf_30_clk),
    .D(net193),
    .SCD(clknet_1_0__leaf_net186),
    .SCE(clknet_1_1__leaf_net183),
    .Q(net196));
 sky130_fd_sc_hd__sdfbbn_1 c206 (.CLK_N(clknet_leaf_30_clk),
    .D(net182),
    .RESET_B(clknet_1_0__leaf_net191),
    .SCD(clknet_1_0__leaf_net186),
    .SCE(net180),
    .SET_B(clknet_1_0__leaf_net183),
    .Q(net198),
    .Q_N(net197));
 sky130_fd_sc_hd__sdfrtp_1 c207 (.CLK(clknet_leaf_30_clk),
    .D(net195),
    .RESET_B(clknet_1_0__leaf_net190),
    .SCD(net197),
    .SCE(clknet_1_0__leaf_net186),
    .Q(net199));
 sky130_fd_sc_hd__a2111o_1 c208 (.A1(net196),
    .A2(net198),
    .B1(net878),
    .C1(clknet_1_1__leaf_net191),
    .D1(net192),
    .X(net200));
 sky130_fd_sc_hd__sdfsbp_1 c209 (.CLK(clknet_leaf_30_clk),
    .D(clknet_1_1__leaf_net188),
    .SCD(net200),
    .SCE(net958),
    .SET_B(clknet_1_0__leaf_net194),
    .Q(net201));
 sky130_fd_sc_hd__dfrbp_1 c210 (.CLK(clknet_leaf_31_clk),
    .D(net954),
    .RESET_B(net73),
    .Q(net203),
    .Q_N(net202));
 sky130_fd_sc_hd__and2_1 c211 (.A(net878),
    .B(net202),
    .X(net204));
 sky130_fd_sc_hd__clkbuf_1 c212 (.A(net204),
    .X(net205));
 sky130_fd_sc_hd__and2_1 c213 (.A(net870),
    .B(net204),
    .X(net206));
 sky130_fd_sc_hd__and2_0 c214 (.A(net205),
    .B(net206),
    .X(net207));
 sky130_fd_sc_hd__and2_1 c215 (.A(net206),
    .B(net204),
    .X(net208));
 sky130_fd_sc_hd__dfrbp_1 c216 (.CLK(clknet_leaf_28_clk),
    .D(net204),
    .RESET_B(net871),
    .Q(net209));
 sky130_fd_sc_hd__dfrtn_1 c217 (.CLK_N(clknet_leaf_30_clk),
    .D(net207),
    .RESET_B(net206),
    .Q(net210));
 sky130_fd_sc_hd__and2_0 c218 (.A(net83),
    .B(net203),
    .X(net211));
 sky130_fd_sc_hd__dfrtp_1 c219 (.CLK(clknet_leaf_30_clk),
    .D(clknet_1_0__leaf_net194),
    .RESET_B(net871),
    .Q(net212));
 sky130_fd_sc_hd__and2_1 c220 (.A(net210),
    .B(net204),
    .X(net213));
 sky130_fd_sc_hd__and2_1 c221 (.A(net209),
    .B(net974),
    .X(net214));
 sky130_fd_sc_hd__dfrtp_1 c222 (.CLK(clknet_leaf_32_clk),
    .D(net73),
    .RESET_B(net213),
    .Q(net215));
 sky130_fd_sc_hd__and2_0 c223 (.A(net213),
    .B(net215),
    .X(net216));
 sky130_fd_sc_hd__dfbbn_1 c224 (.CLK_N(clknet_leaf_27_clk),
    .D(net216),
    .RESET_B(net913),
    .SET_B(net202),
    .Q(net217));
 sky130_fd_sc_hd__and2_1 c225 (.A(net211),
    .B(net928),
    .X(net218));
 sky130_fd_sc_hd__and3_1 c226 (.A(net214),
    .B(net217),
    .C(net218),
    .X(net219));
 sky130_fd_sc_hd__dfbbn_1 c227 (.CLK_N(clknet_leaf_28_clk),
    .D(net219),
    .RESET_B(net218),
    .SET_B(net214),
    .Q(net220));
 sky130_fd_sc_hd__dfbbp_1 c228 (.CLK(clknet_leaf_28_clk),
    .D(net208),
    .RESET_B(net220),
    .SET_B(net218),
    .Q(net221));
 sky130_fd_sc_hd__mux4_1 c229 (.A0(net189),
    .A1(net221),
    .A2(net214),
    .A3(net210),
    .S0(net82),
    .S1(net213),
    .X(net222));
 sky130_fd_sc_hd__sdfxbp_1 c230 (.CLK(clknet_leaf_27_clk),
    .D(net222),
    .SCD(net219),
    .SCE(net204),
    .Q(net224),
    .Q_N(net223));
 sky130_fd_sc_hd__buf_1 c231 (.A(net218),
    .X(net225));
 sky130_fd_sc_hd__clkbuf_1 c232 (.A(net111),
    .X(net226));
 sky130_fd_sc_hd__clkbuf_1 c233 (.A(net770),
    .X(net837));
 sky130_fd_sc_hd__buf_1 c234 (.A(net770),
    .X(net227));
 sky130_fd_sc_hd__dfrtp_1 c235 (.CLK(clknet_leaf_27_clk),
    .D(net225),
    .RESET_B(net846),
    .Q(net228));
 sky130_fd_sc_hd__and2_0 c236 (.A(net227),
    .B(net228),
    .X(net229));
 sky130_fd_sc_hd__and2_0 c237 (.A(net229),
    .B(net228),
    .X(net230));
 sky130_fd_sc_hd__and2_1 c238 (.A(net227),
    .B(net953),
    .X(net231));
 sky130_fd_sc_hd__dfsbp_1 c239 (.CLK(clknet_leaf_27_clk),
    .D(net230),
    .SET_B(net225),
    .Q(net233),
    .Q_N(net232));
 sky130_fd_sc_hd__and2_0 c240 (.A(net231),
    .B(net232),
    .X(net234));
 sky130_fd_sc_hd__and3_1 c241 (.A(net226),
    .B(net233),
    .C(net227),
    .X(net235));
 sky130_fd_sc_hd__a2111o_1 c242 (.A1(net228),
    .A2(net235),
    .B1(net231),
    .C1(net939),
    .D1(net227),
    .X(net236));
 sky130_fd_sc_hd__and2_0 c243 (.A(net234),
    .B(net231),
    .X(net237));
 sky130_fd_sc_hd__dfsbp_1 c244 (.CLK(clknet_leaf_27_clk),
    .D(net236),
    .SET_B(net231),
    .Q(net238));
 sky130_fd_sc_hd__sdfxbp_1 c245 (.CLK(clknet_leaf_26_clk),
    .D(net237),
    .SCD(net235),
    .SCE(net231),
    .Q(net239));
 sky130_fd_sc_hd__and3_1 c246 (.A(net965),
    .B(net227),
    .C(net235),
    .X(net240));
 sky130_fd_sc_hd__dfstp_1 c247 (.CLK(clknet_leaf_27_clk),
    .D(net240),
    .SET_B(net858),
    .Q(net241));
 sky130_fd_sc_hd__and3_1 c248 (.A(net235),
    .B(net227),
    .C(net231),
    .X(net242));
 sky130_fd_sc_hd__sdfxtp_1 c249 (.CLK(clknet_leaf_27_clk),
    .D(net935),
    .SCD(net953),
    .SCE(net242),
    .Q(net243));
 sky130_fd_sc_hd__and2_0 c25 (.A(net804),
    .B(net810),
    .X(net0));
 sky130_fd_sc_hd__dfstp_1 c250 (.CLK(clknet_leaf_26_clk),
    .D(net910),
    .SET_B(net242),
    .Q(net244));
 sky130_fd_sc_hd__sdfxtp_1 c251 (.CLK(clknet_leaf_26_clk),
    .D(net932),
    .SCD(net242),
    .SCE(net235),
    .Q(net245));
 sky130_fd_sc_hd__buf_1 c252 (.A(net127),
    .X(net246));
 sky130_fd_sc_hd__clkbuf_2 c253 (.X(net247));
 sky130_fd_sc_hd__and2_0 c254 (.A(net247),
    .B(clknet_1_0__leaf_net779),
    .X(net248));
 sky130_fd_sc_hd__buf_1 c255 (.A(net873),
    .X(net249));
 sky130_fd_sc_hd__dfstp_1 c256 (.CLK(clknet_leaf_4_clk),
    .D(net246),
    .SET_B(net249),
    .Q(net250));
 sky130_fd_sc_hd__and2_0 c257 (.A(net247),
    .B(clknet_1_0__leaf_net248),
    .X(net251));
 sky130_fd_sc_hd__and2_0 c258 (.A(clknet_1_0__leaf_net251),
    .B(net247),
    .X(net252));
 sky130_fd_sc_hd__dlrbn_1 c259 (.D(clknet_1_1__leaf_net252),
    .GATE_N(clknet_leaf_4_clk),
    .RESET_B(net246),
    .Q(net254),
    .Q_N(net253));
 sky130_fd_sc_hd__and2_0 c26 (.A(net809),
    .B(net810),
    .X(net1));
 sky130_fd_sc_hd__and2_0 c260 (.A(clknet_1_1__leaf_net248),
    .B(net253),
    .X(net255));
 sky130_fd_sc_hd__and2_0 c261 (.A(net254),
    .B(clknet_1_0__leaf_net255),
    .X(net256));
 sky130_fd_sc_hd__dlrbn_1 c262 (.D(clknet_1_0__leaf_net252),
    .GATE_N(clknet_leaf_2_clk),
    .RESET_B(clknet_1_0__leaf_net248),
    .Q(net258),
    .Q_N(net257));
 sky130_fd_sc_hd__dlrbp_1 c263 (.D(clknet_1_1__leaf_net255),
    .GATE(clknet_leaf_5_clk),
    .RESET_B(clknet_1_0__leaf_net256),
    .Q(net260),
    .Q_N(net259));
 sky130_fd_sc_hd__or4bb_1 c264 (.A(net249),
    .B(net260),
    .C_N(net250),
    .D_N(net247),
    .X(net261));
 sky130_fd_sc_hd__and3_1 c265 (.A(net127),
    .B(net261),
    .C(net249),
    .X(net262));
 sky130_fd_sc_hd__or4bb_1 c266 (.A(net250),
    .B(net258),
    .C_N(net253),
    .D_N(net247),
    .X(net263));
 sky130_fd_sc_hd__and2_0 c267 (.A(clknet_1_0__leaf_net251),
    .B(net257),
    .X(net264));
 sky130_fd_sc_hd__sdfsbp_1 c268 (.CLK(clknet_leaf_5_clk),
    .D(net254),
    .SCD(net262),
    .SCE(net957),
    .SET_B(net901),
    .Q(net266),
    .Q_N(net265));
 sky130_fd_sc_hd__sdfxtp_1 c269 (.CLK(clknet_leaf_2_clk),
    .D(clknet_1_0__leaf_net264),
    .SCD(net929),
    .SCE(clknet_1_1__leaf_net251),
    .Q(net267));
 sky130_fd_sc_hd__and3_1 c27 (.A(net811),
    .B(net814),
    .C(net809),
    .X(net2));
 sky130_fd_sc_hd__sdfbbp_1 c270 (.CLK(clknet_leaf_2_clk),
    .D(net262),
    .RESET_B(net267),
    .SCD(net250),
    .SCE(net926),
    .SET_B(clknet_1_0__leaf_net256),
    .Q(net269),
    .Q_N(net268));
 sky130_fd_sc_hd__mux4_1 c271 (.A0(net263),
    .A1(net261),
    .A2(clknet_1_1__leaf_net264),
    .A3(net268),
    .S0(net247),
    .S1(net267),
    .X(net270));
 sky130_fd_sc_hd__and3_1 c272 (.A(net269),
    .B(net265),
    .C(net782),
    .X(net271));
 sky130_fd_sc_hd__and2_1 c273 (.A(net271),
    .B(net144),
    .X(net272));
 sky130_fd_sc_hd__dlrbp_1 c274 (.D(net155),
    .GATE(clknet_leaf_2_clk),
    .RESET_B(net144),
    .Q(net274),
    .Q_N(net273));
 sky130_fd_sc_hd__dlrtn_1 c275 (.D(net272),
    .GATE_N(clknet_leaf_2_clk),
    .RESET_B(net863),
    .Q(net275));
 sky130_fd_sc_hd__dlrtn_1 c276 (.D(net275),
    .GATE_N(clknet_leaf_2_clk),
    .RESET_B(net272),
    .Q(net276));
 sky130_fd_sc_hd__dlrtn_1 c277 (.D(net144),
    .GATE_N(clknet_leaf_1_clk),
    .RESET_B(net272),
    .Q(net277));
 sky130_fd_sc_hd__and2_0 c278 (.A(net259),
    .B(clknet_1_1__leaf_net779),
    .X(net278));
 sky130_fd_sc_hd__dfbbn_1 c279 (.CLK_N(clknet_leaf_2_clk),
    .D(net869),
    .RESET_B(net272),
    .SET_B(net273),
    .Q(net279));
 sky130_fd_sc_hd__and2_0 c28 (.A(net1),
    .B(net810),
    .X(net3));
 sky130_fd_sc_hd__dlrtp_1 c280 (.D(net151),
    .GATE(clknet_leaf_2_clk),
    .RESET_B(net272),
    .Q(net280));
 sky130_fd_sc_hd__and2_0 c281 (.A(net280),
    .B(net144),
    .X(net281));
 sky130_fd_sc_hd__dlrtp_1 c282 (.D(net281),
    .GATE(clknet_leaf_2_clk),
    .RESET_B(net874),
    .Q(net282));
 sky130_fd_sc_hd__dlrtp_1 c283 (.D(net272),
    .GATE(clknet_leaf_2_clk),
    .RESET_B(clknet_1_0__leaf_net278),
    .Q(net283));
 sky130_fd_sc_hd__and2_0 c284 (.A(clknet_1_1__leaf_net278),
    .B(net282),
    .X(net284));
 sky130_fd_sc_hd__and3_1 c285 (.A(net277),
    .B(clknet_1_0__leaf_net278),
    .C(clknet_1_0__leaf_net284),
    .X(net285));
 sky130_fd_sc_hd__and3_1 c286 (.A(net282),
    .B(clknet_1_0__leaf_net284),
    .C(net273),
    .X(net286));
 sky130_fd_sc_hd__and2_0 c287 (.A(clknet_1_1__leaf_net284),
    .B(net274),
    .X(net287));
 sky130_fd_sc_hd__sdfstp_1 c288 (.CLK(clknet_leaf_1_clk),
    .D(net286),
    .SCD(clknet_1_1__leaf_net284),
    .SCE(clknet_1_0__leaf_net285),
    .SET_B(net277),
    .Q(net288));
 sky130_fd_sc_hd__dfbbn_1 c289 (.CLK_N(clknet_leaf_1_clk),
    .D(clknet_1_0__leaf_net287),
    .RESET_B(net282),
    .SET_B(clknet_1_1__leaf_net284),
    .Q(net290),
    .Q_N(net289));
 sky130_fd_sc_hd__and2_0 c29 (.A(net810),
    .B(net809),
    .X(net4));
 sky130_fd_sc_hd__sdfbbn_1 c290 (.CLK_N(clknet_leaf_2_clk),
    .D(net283),
    .RESET_B(clknet_1_0__leaf_net287),
    .SCD(net949),
    .SCE(clknet_1_0__leaf_net284),
    .SET_B(net273),
    .Q(net291));
 sky130_fd_sc_hd__edfxbp_1 c291 (.CLK(clknet_leaf_2_clk),
    .D(net863),
    .DE(clknet_1_1__leaf_net287),
    .Q(net293),
    .Q_N(net292));
 sky130_fd_sc_hd__mux4_1 c292 (.A0(net293),
    .A1(net283),
    .A2(net288),
    .A3(net282),
    .S0(net289),
    .S1(clknet_1_1__leaf_net287),
    .X(net294));
 sky130_fd_sc_hd__or4bb_1 c293 (.A(net291),
    .B(net290),
    .C_N(net282),
    .D_N(net292),
    .X(net295));
 sky130_fd_sc_hd__clkbuf_1 c294 (.A(net167),
    .X(net296));
 sky130_fd_sc_hd__clkbuf_1 c295 (.A(net781),
    .X(net297));
 sky130_fd_sc_hd__edfxtp_1 c296 (.CLK(clknet_leaf_1_clk),
    .D(clknet_1_1__leaf_net285),
    .DE(net297),
    .Q(net298));
 sky130_fd_sc_hd__buf_1 c297 (.A(net784),
    .X(net299));
 sky130_fd_sc_hd__and2_0 c298 (.A(net298),
    .B(net299),
    .X(net300));
 sky130_fd_sc_hd__and2_1 c299 (.A(net296),
    .B(net299),
    .X(net301));
 sky130_fd_sc_hd__and2_0 c30 (.A(net812),
    .B(net809),
    .X(net5));
 sky130_fd_sc_hd__and2_1 c300 (.A(net299),
    .B(net301),
    .X(net302));
 sky130_fd_sc_hd__sdlclkp_1 c301 (.CLK(clknet_leaf_1_clk),
    .GATE(net302),
    .SCE(net973),
    .GCLK(net303));
 sky130_fd_sc_hd__and2_0 c302 (.A(net297),
    .B(net296),
    .X(net304));
 sky130_fd_sc_hd__and2_0 c303 (.A(net304),
    .B(net300),
    .X(net305));
 sky130_fd_sc_hd__sdlclkp_2 c304 (.CLK(clknet_leaf_1_clk),
    .GATE(clknet_1_1__leaf_net303),
    .SCE(net305),
    .GCLK(net306));
 sky130_fd_sc_hd__and2_1 c305 (.A(net300),
    .B(net860),
    .X(net307));
 sky130_fd_sc_hd__sdlclkp_4 c306 (.CLK(clknet_leaf_1_clk),
    .GATE(net307),
    .SCE(net301),
    .GCLK(net308));
 sky130_fd_sc_hd__and2_0 c307 (.A(net172),
    .B(clknet_1_0__leaf_net306),
    .X(net309));
 sky130_fd_sc_hd__dfrbp_1 c308 (.CLK(clknet_leaf_1_clk),
    .D(net305),
    .RESET_B(clknet_1_0__leaf_net308),
    .Q(net311),
    .Q_N(net310));
 sky130_fd_sc_hd__dfrbp_1 c309 (.CLK(clknet_leaf_29_clk),
    .D(net900),
    .RESET_B(net861),
    .Q(net313),
    .Q_N(net312));
 sky130_fd_sc_hd__and2_0 c31 (.A(net8),
    .B(net809),
    .X(net6));
 sky130_fd_sc_hd__dfrtn_1 c310 (.CLK_N(clknet_leaf_1_clk),
    .D(net298),
    .RESET_B(net302),
    .Q(net314));
 sky130_fd_sc_hd__and2_0 c311 (.A(net314),
    .B(net313),
    .X(net315));
 sky130_fd_sc_hd__sdfbbn_1 c312 (.CLK_N(clknet_leaf_1_clk),
    .D(clknet_1_0__leaf_net303),
    .RESET_B(net310),
    .SCD(clknet_1_1__leaf_net308),
    .SCE(net302),
    .SET_B(net298),
    .Q(net316));
 sky130_fd_sc_hd__and3_1 c313 (.A(net315),
    .B(net314),
    .C(net312),
    .X(net317));
 sky130_fd_sc_hd__and3_1 c314 (.A(net316),
    .B(net309),
    .C(clknet_1_1__leaf_net306),
    .X(net318));
 sky130_fd_sc_hd__and2_0 c315 (.A(net317),
    .B(clknet_1_1__leaf_net194),
    .X(net319));
 sky130_fd_sc_hd__dfrtp_2 c316 (.CLK(clknet_leaf_30_clk),
    .D(clknet_1_0__leaf_net319),
    .RESET_B(clknet_1_1__leaf_net186),
    .Q(net320));
 sky130_fd_sc_hd__and2_0 c317 (.A(net48),
    .B(clknet_1_1__leaf_net194),
    .X(net321));
 sky130_fd_sc_hd__dfrtp_1 c318 (.CLK(clknet_leaf_29_clk),
    .D(clknet_1_1__leaf_net319),
    .RESET_B(net847),
    .Q(net322));
 sky130_fd_sc_hd__dfrtp_1 c319 (.CLK(clknet_leaf_29_clk),
    .D(clknet_1_0__leaf_net321),
    .RESET_B(clknet_1_0__leaf_net319),
    .Q(net323));
 sky130_fd_sc_hd__and2_1 c32 (.A(net3),
    .B(net6),
    .X(net7));
 sky130_fd_sc_hd__and2_2 c320 (.A(net841),
    .B(net847),
    .X(net324));
 sky130_fd_sc_hd__dfbbp_1 c321 (.CLK(clknet_leaf_29_clk),
    .D(clknet_1_1__leaf_net319),
    .RESET_B(clknet_1_1__leaf_net321),
    .SET_B(net324),
    .Q(net326),
    .Q_N(net325));
 sky130_fd_sc_hd__and3_1 c322 (.A(net324),
    .B(net320),
    .C(net323),
    .X(net327));
 sky130_fd_sc_hd__dfsbp_1 c323 (.CLK(clknet_leaf_29_clk),
    .D(net317),
    .SET_B(clknet_1_0__leaf_net321),
    .Q(net328));
 sky130_fd_sc_hd__and3_1 c324 (.A(net320),
    .B(net324),
    .C(net327),
    .X(net329));
 sky130_fd_sc_hd__and3_1 c325 (.A(net322),
    .B(net320),
    .C(net325),
    .X(net330));
 sky130_fd_sc_hd__and2_0 c326 (.A(net841),
    .B(net326),
    .X(net331));
 sky130_fd_sc_hd__sdfxbp_1 c327 (.CLK(clknet_leaf_29_clk),
    .D(clknet_1_1__leaf_net321),
    .SCD(net330),
    .SCE(net324),
    .Q(net333),
    .Q_N(net332));
 sky130_fd_sc_hd__and2_0 c328 (.A(net330),
    .B(net327),
    .X(net334));
 sky130_fd_sc_hd__sdfxbp_1 c329 (.CLK(clknet_leaf_29_clk),
    .D(net331),
    .SCD(net330),
    .SCE(clknet_1_0__leaf_net321),
    .Q(net336),
    .Q_N(net335));
 sky130_fd_sc_hd__and3_1 c33 (.A(net816),
    .B(net817),
    .C(net807),
    .X(net8));
 sky130_fd_sc_hd__sdfxtp_1 c330 (.CLK(clknet_leaf_20_clk),
    .D(net334),
    .SCD(net324),
    .SCE(net940),
    .Q(net337));
 sky130_fd_sc_hd__sdfxtp_1 c331 (.CLK(clknet_leaf_20_clk),
    .D(clknet_1_1__leaf_net186),
    .SCD(net894),
    .SCE(net330),
    .Q(net338));
 sky130_fd_sc_hd__mux4_1 c332 (.A0(net327),
    .A1(net336),
    .A2(net338),
    .A3(net330),
    .S0(net324),
    .S1(net301),
    .X(net339));
 sky130_fd_sc_hd__mux4_1 c333 (.A0(net333),
    .A1(net339),
    .A2(net334),
    .A3(clknet_1_1__leaf_net321),
    .S0(clknet_1_1__leaf_net186),
    .S1(net320),
    .X(net340));
 sky130_fd_sc_hd__mux4_1 c334 (.A0(net329),
    .A1(net334),
    .A2(net332),
    .A3(net330),
    .S0(clknet_1_1__leaf_net321),
    .S1(net785),
    .X(net341));
 sky130_fd_sc_hd__mux4_1 c335 (.A0(net963),
    .A1(net336),
    .A2(net320),
    .A3(net327),
    .S0(net785),
    .S1(net786),
    .X(net342));
 sky130_fd_sc_hd__and2_1 c336 (.A(net215),
    .B(net223),
    .X(net343));
 sky130_fd_sc_hd__dlymetal6s2s_1 c337 (.A(net343),
    .X(net344));
 sky130_fd_sc_hd__and2_2 c338 (.A(net344),
    .B(net343),
    .X(net345));
 sky130_fd_sc_hd__dfsbp_1 c339 (.CLK(clknet_leaf_28_clk),
    .D(net345),
    .SET_B(net344),
    .Q(net347),
    .Q_N(net346));
 sky130_fd_sc_hd__and2_0 c34 (.A(net4),
    .B(net6),
    .X(net9));
 sky130_fd_sc_hd__sdfxtp_1 c340 (.CLK(clknet_leaf_28_clk),
    .D(net976),
    .SCD(net858),
    .SCE(net345),
    .Q(net348));
 sky130_fd_sc_hd__and2_0 c341 (.A(net347),
    .B(net325),
    .X(net349));
 sky130_fd_sc_hd__and2_1 c342 (.A(net347),
    .B(net83),
    .X(net350));
 sky130_fd_sc_hd__and2_0 c343 (.A(net350),
    .B(net343),
    .X(net351));
 sky130_fd_sc_hd__and2_0 c344 (.A(net349),
    .B(net343),
    .X(net352));
 sky130_fd_sc_hd__dfstp_1 c345 (.CLK(clknet_leaf_28_clk),
    .D(net343),
    .SET_B(net345),
    .Q(net353));
 sky130_fd_sc_hd__and2_1 c346 (.A(net969),
    .B(net351),
    .X(net354));
 sky130_fd_sc_hd__dfstp_1 c347 (.CLK(clknet_leaf_28_clk),
    .D(net345),
    .SET_B(net354),
    .Q(net355));
 sky130_fd_sc_hd__sdfstp_1 c348 (.CLK(clknet_leaf_21_clk),
    .D(net349),
    .SCD(net355),
    .SCE(net345),
    .SET_B(net855),
    .Q(net356));
 sky130_fd_sc_hd__dfbbn_1 c349 (.CLK_N(clknet_leaf_28_clk),
    .D(net350),
    .RESET_B(net354),
    .SET_B(net353),
    .Q(net357));
 sky130_fd_sc_hd__dfbbn_1 c35 (.CLK_N(clknet_leaf_3_clk),
    .D(net5),
    .RESET_B(net809),
    .SET_B(net7),
    .Q(net11),
    .Q_N(net10));
 sky130_fd_sc_hd__and3_1 c350 (.A(net356),
    .B(net355),
    .C(net350),
    .X(net358));
 sky130_fd_sc_hd__and2_0 c351 (.A(net922),
    .B(net355),
    .X(net359));
 sky130_fd_sc_hd__and2_0 c352 (.A(net351),
    .B(net344),
    .X(net360));
 sky130_fd_sc_hd__and2_0 c353 (.A(net352),
    .B(net355),
    .X(net361));
 sky130_fd_sc_hd__dfstp_1 c354 (.CLK(clknet_leaf_26_clk),
    .D(net360),
    .SET_B(net354),
    .Q(net362));
 sky130_fd_sc_hd__and2_0 c355 (.A(net358),
    .B(net349),
    .X(net363));
 sky130_fd_sc_hd__dfbbn_1 c356 (.CLK_N(clknet_leaf_21_clk),
    .D(net363),
    .RESET_B(net355),
    .SET_B(net346),
    .Q(net364));
 sky130_fd_sc_hd__buf_1 c357 (.A(net892),
    .X(net365));
 sky130_fd_sc_hd__and2_1 c358 (.A(net228),
    .B(net223),
    .X(net366));
 sky130_fd_sc_hd__and2_1 c359 (.A(net867),
    .B(net365),
    .X(net367));
 sky130_fd_sc_hd__dfbbn_1 c36 (.CLK_N(clknet_leaf_36_clk),
    .D(net9),
    .RESET_B(net904),
    .SET_B(net810),
    .Q(net13),
    .Q_N(net12));
 sky130_fd_sc_hd__and2_0 c360 (.A(net365),
    .B(net344),
    .X(net368));
 sky130_fd_sc_hd__or4bb_2 c361 (.A(net362),
    .B(net367),
    .C_N(net218),
    .D_N(net365),
    .X(net369));
 sky130_fd_sc_hd__dfbbp_1 c362 (.CLK(clknet_leaf_26_clk),
    .D(net368),
    .RESET_B(net369),
    .SET_B(net365),
    .Q(net371),
    .Q_N(net370));
 sky130_fd_sc_hd__clkbuf_1 c363 (.A(net933),
    .X(net372));
 sky130_fd_sc_hd__and2_1 c364 (.A(net372),
    .B(net367),
    .X(net373));
 sky130_fd_sc_hd__sdfxbp_1 c365 (.CLK(clknet_leaf_21_clk),
    .D(net359),
    .SCD(net373),
    .SCE(net371),
    .Q(net375),
    .Q_N(net374));
 sky130_fd_sc_hd__sdfxbp_1 c366 (.CLK(clknet_leaf_24_clk),
    .D(net367),
    .SCD(net369),
    .SCE(net955),
    .Q(net377),
    .Q_N(net376));
 sky130_fd_sc_hd__and2_1 c367 (.A(net357),
    .B(net377),
    .X(net378));
 sky130_fd_sc_hd__and3_1 c368 (.A(net239),
    .B(net371),
    .C(net375),
    .X(net379));
 sky130_fd_sc_hd__and2_0 c369 (.A(net378),
    .B(net371),
    .X(net380));
 sky130_fd_sc_hd__and2_0 c37 (.A(net13),
    .B(net10),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 c370 (.A(net754),
    .X(net381));
 sky130_fd_sc_hd__sdfstp_1 c371 (.CLK(clknet_leaf_26_clk),
    .D(net380),
    .SCD(net371),
    .SCE(net373),
    .SET_B(net367),
    .Q(net382));
 sky130_fd_sc_hd__sedfxbp_1 c372 (.CLK(clknet_leaf_26_clk),
    .D(net977),
    .DE(net382),
    .SCD(net373),
    .SCE(net370),
    .Q(net383));
 sky130_fd_sc_hd__mux4_1 c373 (.A0(net381),
    .A1(net367),
    .A2(net378),
    .A3(net365),
    .S0(net369),
    .S1(net370),
    .X(net384));
 sky130_fd_sc_hd__and2_0 c374 (.A(net962),
    .B(net378),
    .X(net385));
 sky130_fd_sc_hd__and3_1 c375 (.A(net378),
    .B(net380),
    .C(net787),
    .X(net386));
 sky130_fd_sc_hd__sdfxtp_1 c376 (.CLK(clknet_leaf_25_clk),
    .D(net385),
    .SCD(net386),
    .SCE(net787),
    .Q(net387));
 sky130_fd_sc_hd__sedfxbp_1 c377 (.CLK(clknet_leaf_24_clk),
    .D(net379),
    .DE(net387),
    .SCD(net381),
    .SCE(net369),
    .Q(net388));
 sky130_fd_sc_hd__clkbuf_1 c378 (.A(net775),
    .X(net389));
 sky130_fd_sc_hd__clkbuf_1 c379 (.A(net389),
    .X(net390));
 sky130_fd_sc_hd__dfbbp_1 c38 (.CLK(clknet_leaf_36_clk),
    .D(net14),
    .RESET_B(net11),
    .SET_B(net7),
    .Q(net15));
 sky130_fd_sc_hd__clkbuf_1 c380 (.A(net390),
    .X(net391));
 sky130_fd_sc_hd__and2_1 c381 (.A(net271),
    .B(net389),
    .X(net392));
 sky130_fd_sc_hd__sdfxtp_1 c382 (.CLK(clknet_leaf_8_clk),
    .D(net391),
    .SCD(net392),
    .SCE(clknet_1_1__leaf_net256),
    .Q(net393));
 sky130_fd_sc_hd__and2_0 c383 (.A(net389),
    .B(net393),
    .X(net394));
 sky130_fd_sc_hd__and2_2 c384 (.A(net914),
    .B(net392),
    .X(net395));
 sky130_fd_sc_hd__and3_1 c385 (.A(net914),
    .B(net392),
    .C(net394),
    .X(net396));
 sky130_fd_sc_hd__sdfxtp_1 c386 (.CLK(clknet_leaf_7_clk),
    .D(net390),
    .SCD(net394),
    .SCE(net395),
    .Q(net397));
 sky130_fd_sc_hd__dfbbn_1 c387 (.CLK_N(clknet_leaf_7_clk),
    .D(net391),
    .RESET_B(net395),
    .SET_B(net392),
    .Q(net399),
    .Q_N(net398));
 sky130_fd_sc_hd__clkbuf_1 c388 (.A(net774),
    .X(net400));
 sky130_fd_sc_hd__and2_0 c389 (.A(net394),
    .B(net398),
    .X(net401));
 sky130_fd_sc_hd__and3_1 c39 (.A(net0),
    .B(net13),
    .C(net809),
    .X(net16));
 sky130_fd_sc_hd__and2_2 c390 (.A(net260),
    .B(net401),
    .X(net402));
 sky130_fd_sc_hd__dlrbn_1 c391 (.D(net401),
    .GATE_N(clknet_leaf_7_clk),
    .RESET_B(net396),
    .Q(net404),
    .Q_N(net403));
 sky130_fd_sc_hd__dfbbn_1 c392 (.CLK_N(clknet_leaf_5_clk),
    .D(net397),
    .RESET_B(net402),
    .SET_B(net395),
    .Q(net406),
    .Q_N(net405));
 sky130_fd_sc_hd__dfbbp_1 c393 (.CLK(clknet_leaf_5_clk),
    .D(net406),
    .RESET_B(net404),
    .SET_B(net395),
    .Q(net408),
    .Q_N(net407));
 sky130_fd_sc_hd__dlrbn_1 c394 (.D(net395),
    .GATE_N(clknet_leaf_8_clk),
    .RESET_B(net399),
    .Q(net410),
    .Q_N(net409));
 sky130_fd_sc_hd__and2_0 c395 (.A(net400),
    .B(net405),
    .X(net411));
 sky130_fd_sc_hd__and3_1 c396 (.A(net392),
    .B(net400),
    .C(net397),
    .X(net412));
 sky130_fd_sc_hd__sdfbbp_1 c397 (.CLK(clknet_leaf_7_clk),
    .D(net404),
    .RESET_B(net412),
    .SCD(net411),
    .SCE(net402),
    .SET_B(net392),
    .Q(net413));
 sky130_fd_sc_hd__mux4_1 c398 (.A0(net413),
    .A1(net411),
    .A2(net403),
    .A3(net395),
    .S0(net412),
    .S1(net402),
    .X(net414));
 sky130_fd_sc_hd__clkbuf_1 c399 (.A(net756),
    .X(net415));
 sky130_fd_sc_hd__a2111o_1 c40 (.A1(net809),
    .A2(net14),
    .B1(net952),
    .C1(net16),
    .D1(net810),
    .X(net17));
 sky130_fd_sc_hd__buf_1 c400 (.A(net756),
    .X(net416));
 sky130_fd_sc_hd__and2_0 c401 (.A(net416),
    .B(net788),
    .X(net417));
 sky130_fd_sc_hd__dlrbp_1 c402 (.D(net415),
    .GATE(clknet_leaf_8_clk),
    .RESET_B(net402),
    .Q(net419),
    .Q_N(net418));
 sky130_fd_sc_hd__and2_1 c403 (.A(net418),
    .B(net788),
    .X(net420));
 sky130_fd_sc_hd__and2_1 c404 (.A(net417),
    .B(net420),
    .X(net421));
 sky130_fd_sc_hd__and2_0 c405 (.A(net415),
    .B(net420),
    .X(net422));
 sky130_fd_sc_hd__dlrbp_1 c406 (.D(net420),
    .GATE(clknet_leaf_8_clk),
    .RESET_B(net402),
    .Q(net424),
    .Q_N(net423));
 sky130_fd_sc_hd__and2_0 c407 (.A(net420),
    .B(net783),
    .X(net425));
 sky130_fd_sc_hd__and2_0 c408 (.A(net422),
    .B(net425),
    .X(net426));
 sky130_fd_sc_hd__and2_1 c409 (.A(net417),
    .B(net422),
    .X(net427));
 sky130_fd_sc_hd__sdfbbn_1 c41 (.CLK_N(clknet_leaf_36_clk),
    .D(net6),
    .RESET_B(net17),
    .SCD(net803),
    .SCE(net810),
    .SET_B(net4),
    .Q(net18));
 sky130_fd_sc_hd__dlrtn_1 c410 (.D(net943),
    .GATE_N(clknet_leaf_9_clk),
    .RESET_B(net427),
    .Q(net428));
 sky130_fd_sc_hd__and3_1 c411 (.A(net425),
    .B(net428),
    .C(net423),
    .X(net429));
 sky130_fd_sc_hd__sdfxbp_1 c412 (.CLK(clknet_leaf_8_clk),
    .D(net427),
    .SCD(net429),
    .SCE(net943),
    .Q(net431),
    .Q_N(net430));
 sky130_fd_sc_hd__sdfxbp_1 c413 (.CLK(clknet_leaf_9_clk),
    .D(net907),
    .SCD(net426),
    .SCE(net428),
    .Q(net433),
    .Q_N(net432));
 sky130_fd_sc_hd__sdfxtp_2 c414 (.CLK(clknet_leaf_9_clk),
    .D(net429),
    .SCD(net943),
    .SCE(net427),
    .Q(net434));
 sky130_fd_sc_hd__a2111o_1 c415 (.A1(net416),
    .A2(net430),
    .B1(net432),
    .C1(net434),
    .D1(net420),
    .X(net435));
 sky130_fd_sc_hd__sdfxtp_1 c416 (.CLK(clknet_leaf_9_clk),
    .D(net426),
    .SCD(net435),
    .SCE(net937),
    .Q(net436));
 sky130_fd_sc_hd__a2111o_1 c417 (.A1(net433),
    .A2(net434),
    .B1(net436),
    .C1(net423),
    .D1(net420),
    .X(net437));
 sky130_fd_sc_hd__mux4_1 c418 (.A0(net436),
    .A1(net433),
    .A2(net437),
    .A3(net423),
    .S0(net435),
    .S1(net938),
    .X(net438));
 sky130_fd_sc_hd__sedfxtp_1 c419 (.CLK(clknet_leaf_9_clk),
    .D(net979),
    .DE(net435),
    .SCD(net438),
    .SCE(net937),
    .Q(net439));
 sky130_fd_sc_hd__buf_1 c42 (.A(in14),
    .X(net19));
 sky130_fd_sc_hd__buf_1 c420 (.A(net888),
    .X(net440));
 sky130_fd_sc_hd__dlymetal6s2s_1 c421 (.A(net301),
    .X(net441));
 sky130_fd_sc_hd__clkbuf_1 c422 (.A(net755),
    .X(net442));
 sky130_fd_sc_hd__dlrtn_1 c423 (.D(net441),
    .GATE_N(clknet_leaf_20_clk),
    .RESET_B(net440),
    .Q(net443));
 sky130_fd_sc_hd__dlrtn_1 c424 (.D(clknet_1_1__leaf_net318),
    .GATE_N(clknet_leaf_9_clk),
    .RESET_B(net428),
    .Q(net444));
 sky130_fd_sc_hd__buf_1 c425 (.A(net439),
    .X(net445));
 sky130_fd_sc_hd__sdfxtp_1 c426 (.CLK(clknet_leaf_20_clk),
    .D(net445),
    .SCD(net443),
    .SCE(net441),
    .Q(net446));
 sky130_fd_sc_hd__and2_1 c427 (.A(net434),
    .B(net444),
    .X(net447));
 sky130_fd_sc_hd__and3_1 c428 (.A(net442),
    .B(net447),
    .C(net446),
    .X(net448));
 sky130_fd_sc_hd__dfbbn_1 c429 (.CLK_N(clknet_leaf_19_clk),
    .D(net445),
    .RESET_B(net448),
    .SET_B(net441),
    .Q(net450),
    .Q_N(net449));
 sky130_fd_sc_hd__clkbuf_2 c43 (.A(net19),
    .X(net20));
 sky130_fd_sc_hd__and2_0 c430 (.A(net446),
    .B(net449),
    .X(net451));
 sky130_fd_sc_hd__and2_0 c431 (.A(net450),
    .B(net447),
    .X(net452));
 sky130_fd_sc_hd__and2_1 c432 (.A(net451),
    .B(net447),
    .X(net453));
 sky130_fd_sc_hd__and2_1 c433 (.A(net453),
    .B(net452),
    .X(net454));
 sky130_fd_sc_hd__and3_1 c434 (.A(net421),
    .B(net453),
    .C(net451),
    .X(net455));
 sky130_fd_sc_hd__dfbbn_1 c435 (.CLK_N(clknet_leaf_19_clk),
    .D(net447),
    .RESET_B(net455),
    .SET_B(net454),
    .Q(net456));
 sky130_fd_sc_hd__dlrtp_1 c436 (.D(net455),
    .GATE(clknet_leaf_19_clk),
    .RESET_B(net454),
    .Q(net457));
 sky130_fd_sc_hd__and3_1 c437 (.A(net452),
    .B(net891),
    .C(net457),
    .X(net458));
 sky130_fd_sc_hd__dfbbp_1 c438 (.CLK(clknet_leaf_19_clk),
    .D(net444),
    .RESET_B(net456),
    .SET_B(net458),
    .Q(net460),
    .Q_N(net459));
 sky130_fd_sc_hd__sdfbbn_1 c439 (.CLK_N(clknet_leaf_19_clk),
    .D(net458),
    .RESET_B(net441),
    .SCD(net460),
    .SCE(net453),
    .SET_B(net445),
    .Q(net461));
 sky130_fd_sc_hd__and2_1 c44 (.A(net16),
    .B(net20),
    .X(net21));
 sky130_fd_sc_hd__and3_1 c440 (.A(net443),
    .B(net447),
    .C(net459),
    .X(net462));
 sky130_fd_sc_hd__clkbuf_1 c441 (.A(net448),
    .X(net463));
 sky130_fd_sc_hd__buf_1 c442 (.A(net765),
    .X(net464));
 sky130_fd_sc_hd__clkbuf_2 c443 (.A(net872),
    .X(net465));
 sky130_fd_sc_hd__buf_1 c444 (.A(net764),
    .X(net466));
 sky130_fd_sc_hd__and2_2 c445 (.A(net462),
    .B(net466),
    .X(net467));
 sky130_fd_sc_hd__sdfxbp_1 c446 (.CLK(clknet_leaf_21_clk),
    .D(net464),
    .SCD(net467),
    .SCE(net465),
    .Q(net469),
    .Q_N(net468));
 sky130_fd_sc_hd__and2_1 c447 (.A(net464),
    .B(net468),
    .X(net470));
 sky130_fd_sc_hd__and2_0 c448 (.A(net328),
    .B(net466),
    .X(net471));
 sky130_fd_sc_hd__and2_1 c449 (.A(net465),
    .B(net470),
    .X(net472));
 sky130_fd_sc_hd__and2_1 c45 (.A(net20),
    .B(net19),
    .X(net22));
 sky130_fd_sc_hd__and3_1 c450 (.A(net469),
    .B(net465),
    .C(net470),
    .X(net473));
 sky130_fd_sc_hd__and3_1 c451 (.A(net471),
    .B(net470),
    .C(net466),
    .X(net474));
 sky130_fd_sc_hd__dlrtp_1 c452 (.D(net470),
    .GATE(clknet_leaf_19_clk),
    .RESET_B(net463),
    .Q(net475));
 sky130_fd_sc_hd__and2_0 c453 (.A(net461),
    .B(net475),
    .X(net476));
 sky130_fd_sc_hd__and2_1 c454 (.A(net476),
    .B(net475),
    .X(net477));
 sky130_fd_sc_hd__and3_1 c455 (.A(net473),
    .B(net474),
    .C(net468),
    .X(net478));
 sky130_fd_sc_hd__mux4_1 c456 (.A0(net469),
    .A1(net477),
    .A2(net476),
    .A3(net459),
    .S0(net467),
    .S1(net470),
    .X(net479));
 sky130_fd_sc_hd__or4bb_1 c457 (.A(net464),
    .B(net471),
    .C_N(net470),
    .D_N(net981),
    .X(net480));
 sky130_fd_sc_hd__and3_1 c458 (.A(net326),
    .B(net472),
    .C(net480),
    .X(net481));
 sky130_fd_sc_hd__sdfxbp_1 c459 (.CLK(clknet_leaf_22_clk),
    .D(net480),
    .SCD(net481),
    .SCE(net473),
    .Q(net482));
 sky130_fd_sc_hd__clkbuf_1 c46 (.X(net23));
 sky130_fd_sc_hd__sdfxtp_1 c460 (.CLK(clknet_leaf_22_clk),
    .D(net478),
    .SCD(net902),
    .SCE(net472),
    .Q(net483));
 sky130_fd_sc_hd__and2_0 c461 (.A(net474),
    .B(net931),
    .X(net484));
 sky130_fd_sc_hd__buf_1 c462 (.A(net771),
    .X(net485));
 sky130_fd_sc_hd__clkbuf_1 c463 (.A(net485),
    .X(net486));
 sky130_fd_sc_hd__dlrtp_1 c464 (.D(net467),
    .GATE(clknet_leaf_21_clk),
    .RESET_B(net477),
    .Q(net487));
 sky130_fd_sc_hd__and2_1 c465 (.A(net486),
    .B(net477),
    .X(net488));
 sky130_fd_sc_hd__and2_0 c466 (.A(net344),
    .B(net850),
    .X(net489));
 sky130_fd_sc_hd__sdfxtp_1 c467 (.CLK(clknet_leaf_21_clk),
    .D(net850),
    .SCD(net488),
    .SCE(net467),
    .Q(net490));
 sky130_fd_sc_hd__buf_1 c468 (.A(net470),
    .X(net820));
 sky130_fd_sc_hd__and2_0 c469 (.A(net440),
    .B(net485),
    .X(net491));
 sky130_fd_sc_hd__buf_1 c47 (.A(net745),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_1 c470 (.A(net771),
    .X(net492));
 sky130_fd_sc_hd__clkbuf_1 c471 (.A(net485),
    .X(net493));
 sky130_fd_sc_hd__edfxbp_1 c472 (.CLK(clknet_leaf_21_clk),
    .D(net361),
    .DE(net488),
    .Q(net495),
    .Q_N(net494));
 sky130_fd_sc_hd__and2_0 c473 (.A(net490),
    .B(net495),
    .X(net496));
 sky130_fd_sc_hd__and3_1 c474 (.A(net486),
    .B(net495),
    .C(net477),
    .X(net497));
 sky130_fd_sc_hd__sdfxtp_1 c475 (.CLK(clknet_leaf_22_clk),
    .D(net497),
    .SCD(net488),
    .SCE(net494),
    .Q(net498));
 sky130_fd_sc_hd__and3_1 c476 (.A(net466),
    .B(net492),
    .C(net495),
    .X(net499));
 sky130_fd_sc_hd__and3_1 c477 (.A(net956),
    .B(net495),
    .C(net820),
    .X(net500));
 sky130_fd_sc_hd__dfbbn_1 c478 (.CLK_N(clknet_leaf_21_clk),
    .D(net500),
    .RESET_B(net493),
    .SET_B(net495),
    .Q(net502),
    .Q_N(net501));
 sky130_fd_sc_hd__or4bb_1 c479 (.A(net491),
    .B(net499),
    .C_N(net501),
    .D_N(net494),
    .X(net503));
 sky130_fd_sc_hd__and2_0 c48 (.A(net15),
    .B(net23),
    .X(net25));
 sky130_fd_sc_hd__a2111o_1 c480 (.A1(net503),
    .A2(net496),
    .B1(net499),
    .C1(net501),
    .D1(net494),
    .X(net504));
 sky130_fd_sc_hd__sdfbbn_1 c481 (.CLK_N(clknet_leaf_21_clk),
    .D(net496),
    .RESET_B(net490),
    .SCD(net917),
    .SCE(net494),
    .SET_B(net467),
    .Q(net505));
 sky130_fd_sc_hd__dfbbn_1 c482 (.CLK_N(clknet_leaf_22_clk),
    .D(net917),
    .RESET_B(net504),
    .SET_B(net905),
    .Q(net829));
 sky130_fd_sc_hd__dfxbp_1 c487 (.CLK(clknet_leaf_24_clk),
    .D(net484),
    .Q(net836),
    .Q_N(net827));
 sky130_fd_sc_hd__and2_1 c488 (.A(net388),
    .B(net827),
    .X(net506));
 sky130_fd_sc_hd__and2_1 c489 (.A(net366),
    .B(net506),
    .X(net507));
 sky130_fd_sc_hd__dfrbp_1 c49 (.CLK(clknet_leaf_35_clk),
    .D(net22),
    .RESET_B(net20),
    .Q(net27),
    .Q_N(net26));
 sky130_fd_sc_hd__buf_1 c490 (.A(net507),
    .X(net508));
 sky130_fd_sc_hd__and2_0 c491 (.A(net836),
    .B(net506),
    .X(net509));
 sky130_fd_sc_hd__dfxbp_1 c492 (.CLK(clknet_leaf_24_clk),
    .D(net508),
    .Q(net511),
    .Q_N(net510));
 sky130_fd_sc_hd__and3_1 c493 (.A(net506),
    .B(net509),
    .C(net510),
    .X(net512));
 sky130_fd_sc_hd__edfxtp_1 c494 (.CLK(clknet_leaf_24_clk),
    .D(net508),
    .DE(net967),
    .Q(net513));
 sky130_fd_sc_hd__dfbbp_1 c495 (.CLK(clknet_leaf_24_clk),
    .D(net509),
    .RESET_B(net512),
    .SET_B(net875),
    .Q(net833),
    .Q_N(net514));
 sky130_fd_sc_hd__or4bb_1 c496 (.A(net506),
    .B(net513),
    .C_N(net833),
    .D_N(net510),
    .X(net832));
 sky130_fd_sc_hd__sedfxtp_4 c497 (.CLK(clknet_leaf_24_clk),
    .D(net833),
    .DE(net511),
    .SCD(net508),
    .SCE(net513),
    .Q(net825));
 sky130_fd_sc_hd__a2111o_1 c498 (.A1(net509),
    .A2(net507),
    .B1(net833),
    .C1(net825),
    .D1(net510),
    .X(net834));
 sky130_fd_sc_hd__or4bb_1 c499 (.A(net511),
    .B(net825),
    .C_N(net514),
    .D_N(net513),
    .X(net831));
 sky130_fd_sc_hd__dfrbp_1 c50 (.CLK(clknet_leaf_36_clk),
    .D(net7),
    .RESET_B(net24),
    .Q(net29),
    .Q_N(net28));
 sky130_fd_sc_hd__sdfbbp_1 c500 (.CLK(clknet_leaf_24_clk),
    .D(net513),
    .RESET_B(net512),
    .SCD(net832),
    .SCE(net825),
    .SET_B(net877),
    .Q(net823),
    .Q_N(net826));
 sky130_fd_sc_hd__mux4_1 c501 (.A0(net507),
    .A1(net834),
    .A2(net832),
    .A3(net831),
    .S0(net825),
    .S1(net513),
    .X(net515));
 sky130_fd_sc_hd__mux4_1 c502 (.A0(net513),
    .A1(net831),
    .A2(net511),
    .A3(net514),
    .S0(net825),
    .S1(net835),
    .X(net516));
 sky130_fd_sc_hd__mux4_1 c503 (.A0(net512),
    .A1(net516),
    .A2(net834),
    .A3(net825),
    .S0(net514),
    .S1(net510),
    .X(net517));
 sky130_fd_sc_hd__sdlclkp_1 c504 (.CLK(clknet_leaf_7_clk),
    .GATE(net899),
    .SCE(net402),
    .GCLK(net518));
 sky130_fd_sc_hd__sdlclkp_2 c505 (.CLK(clknet_leaf_7_clk),
    .GATE(clknet_1_0__leaf_net518),
    .SCE(net402),
    .GCLK(net519));
 sky130_fd_sc_hd__sdlclkp_4 c506 (.CLK(clknet_leaf_8_clk),
    .GATE(clknet_1_0__leaf_net519),
    .SCE(clknet_1_1__leaf_net256),
    .GCLK(net520));
 sky130_fd_sc_hd__and2_0 c507 (.A(clknet_1_1__leaf_net520),
    .B(clknet_1_0__leaf_net519),
    .X(net521));
 sky130_fd_sc_hd__and2_0 c508 (.A(clknet_1_1__leaf_net518),
    .B(clknet_1_1__leaf_net519),
    .X(net522));
 sky130_fd_sc_hd__and2_0 c509 (.A(clknet_1_0__leaf_net520),
    .B(net788),
    .X(net523));
 sky130_fd_sc_hd__dfrtn_1 c51 (.CLK_N(clknet_leaf_37_clk),
    .D(net21),
    .RESET_B(net19),
    .Q(net30));
 sky130_fd_sc_hd__and2_0 c510 (.A(clknet_1_1__leaf_net519),
    .B(clknet_1_1__leaf_net521),
    .X(net524));
 sky130_fd_sc_hd__and2_0 c511 (.A(clknet_1_0__leaf_net523),
    .B(clknet_1_0__leaf_net519),
    .X(net525));
 sky130_fd_sc_hd__and2_0 c512 (.A(clknet_1_0__leaf_net524),
    .B(clknet_1_1__leaf_net523),
    .X(net526));
 sky130_fd_sc_hd__and2_0 c513 (.A(clknet_1_1__leaf_net525),
    .B(clknet_1_1__leaf_net519),
    .X(net527));
 sky130_fd_sc_hd__dfrbp_1 c514 (.CLK(clknet_leaf_6_clk),
    .D(net526),
    .RESET_B(clknet_1_1__leaf_net524),
    .Q(net529),
    .Q_N(net528));
 sky130_fd_sc_hd__and2_0 c515 (.A(net522),
    .B(clknet_1_0__leaf_net525),
    .X(net530));
 sky130_fd_sc_hd__dfrbp_1 c516 (.CLK(clknet_leaf_6_clk),
    .D(net882),
    .RESET_B(clknet_1_1__leaf_net530),
    .Q(net532),
    .Q_N(net531));
 sky130_fd_sc_hd__dfrtn_1 c517 (.CLK_N(clknet_leaf_7_clk),
    .D(net868),
    .RESET_B(clknet_1_0__leaf_net530),
    .Q(net533));
 sky130_fd_sc_hd__sdfbbn_1 c518 (.CLK_N(clknet_leaf_6_clk),
    .D(net532),
    .RESET_B(net528),
    .SCD(clknet_1_1__leaf_net530),
    .SCE(clknet_1_1__leaf_net521),
    .SET_B(clknet_1_1__leaf_net519),
    .Q(net534));
 sky130_fd_sc_hd__dfrtp_1 c519 (.CLK(clknet_leaf_6_clk),
    .D(net534),
    .RESET_B(clknet_1_1__leaf_net527),
    .Q(net535));
 sky130_fd_sc_hd__sdfxbp_1 c52 (.CLK(clknet_leaf_35_clk),
    .D(net918),
    .SCD(net22),
    .SCE(net20),
    .Q(net32),
    .Q_N(net31));
 sky130_fd_sc_hd__dfrtp_1 c520 (.CLK(clknet_leaf_7_clk),
    .D(net916),
    .RESET_B(clknet_1_0__leaf_net530),
    .Q(net536));
 sky130_fd_sc_hd__and3_1 c521 (.A(net536),
    .B(net535),
    .C(net533),
    .X(net537));
 sky130_fd_sc_hd__sdfbbn_1 c522 (.CLK_N(clknet_leaf_7_clk),
    .D(net880),
    .RESET_B(clknet_1_0__leaf_net527),
    .SCD(net537),
    .SCE(clknet_1_0__leaf_net530),
    .SET_B(clknet_1_0__leaf_net521),
    .Q(net538));
 sky130_fd_sc_hd__and2_0 c523 (.A(net538),
    .B(net531),
    .X(net539));
 sky130_fd_sc_hd__and2_1 c524 (.A(net539),
    .B(net537),
    .X(net540));
 sky130_fd_sc_hd__dfrtp_1 c525 (.CLK(clknet_leaf_8_clk),
    .D(net438),
    .RESET_B(net843),
    .Q(net541));
 sky130_fd_sc_hd__clkbuf_1 c526 (.A(net920),
    .X(net542));
 sky130_fd_sc_hd__and2_2 c527 (.A(net920),
    .B(net144),
    .X(net543));
 sky130_fd_sc_hd__dfsbp_1 c528 (.CLK(clknet_leaf_8_clk),
    .D(net540),
    .SET_B(net543),
    .Q(net545),
    .Q_N(net544));
 sky130_fd_sc_hd__and2_1 c529 (.A(net545),
    .B(net920),
    .X(net546));
 sky130_fd_sc_hd__and3_1 c53 (.A(net29),
    .B(net24),
    .C(net31),
    .X(net33));
 sky130_fd_sc_hd__and2_1 c530 (.A(net923),
    .B(net545),
    .X(net547));
 sky130_fd_sc_hd__dfsbp_1 c531 (.CLK(clknet_leaf_8_clk),
    .D(net920),
    .SET_B(net543),
    .Q(net548));
 sky130_fd_sc_hd__dfstp_1 c532 (.CLK(clknet_leaf_8_clk),
    .D(net543),
    .SET_B(net547),
    .Q(net549));
 sky130_fd_sc_hd__and2_0 c533 (.A(net279),
    .B(net547),
    .X(net550));
 sky130_fd_sc_hd__and2_0 c534 (.A(net547),
    .B(net546),
    .X(net551));
 sky130_fd_sc_hd__and3_1 c535 (.A(net549),
    .B(clknet_1_0__leaf_net521),
    .C(net546),
    .X(net552));
 sky130_fd_sc_hd__and2_2 c536 (.A(net542),
    .B(net546),
    .X(net553));
 sky130_fd_sc_hd__and2_0 c537 (.A(net545),
    .B(net553),
    .X(net554));
 sky130_fd_sc_hd__sdfxbp_1 c538 (.CLK(clknet_leaf_8_clk),
    .D(net550),
    .SCD(net553),
    .SCE(net543),
    .Q(net555));
 sky130_fd_sc_hd__sdfxbp_1 c539 (.CLK(clknet_leaf_10_clk),
    .D(net552),
    .SCD(net554),
    .SCE(net937),
    .Q(net556));
 sky130_fd_sc_hd__sdfxbp_1 c54 (.CLK(clknet_leaf_36_clk),
    .D(net22),
    .SCD(net918),
    .SCE(net24),
    .Q(net35),
    .Q_N(net34));
 sky130_fd_sc_hd__and3_1 c540 (.A(net555),
    .B(net541),
    .C(net547),
    .X(net557));
 sky130_fd_sc_hd__and3_1 c541 (.A(net428),
    .B(net553),
    .C(net546),
    .X(net558));
 sky130_fd_sc_hd__sedfxtp_1 c542 (.CLK(clknet_leaf_6_clk),
    .D(net548),
    .DE(net558),
    .SCD(net945),
    .SCE(net553),
    .Q(net559));
 sky130_fd_sc_hd__sdfrbp_1 c543 (.CLK(clknet_leaf_11_clk),
    .D(net546),
    .RESET_B(net845),
    .SCD(net558),
    .SCE(net544),
    .Q(net560));
 sky130_fd_sc_hd__sdfrbp_1 c544 (.CLK(clknet_leaf_10_clk),
    .D(net890),
    .RESET_B(net558),
    .SCD(net547),
    .SCE(net543),
    .Q(net561));
 sky130_fd_sc_hd__sdfrtn_1 c545 (.CLK_N(clknet_leaf_10_clk),
    .D(net561),
    .RESET_B(net557),
    .SCD(net421),
    .SCE(net558),
    .Q(net562));
 sky130_fd_sc_hd__dlymetal6s2s_1 c546 (.A(net460),
    .X(net563));
 sky130_fd_sc_hd__clkbuf_2 c547 (.A(net563),
    .X(net564));
 sky130_fd_sc_hd__and2_0 c548 (.A(net564),
    .B(net563),
    .X(net565));
 sky130_fd_sc_hd__and2_0 c549 (.A(net437),
    .B(clknet_1_0__leaf_net521),
    .X(net566));
 sky130_fd_sc_hd__and2_0 c55 (.A(net33),
    .B(net798),
    .X(net36));
 sky130_fd_sc_hd__sdfxtp_1 c550 (.CLK(clknet_leaf_10_clk),
    .D(net563),
    .SCD(clknet_1_0__leaf_net566),
    .SCE(net564),
    .Q(net567));
 sky130_fd_sc_hd__and2_0 c551 (.A(net564),
    .B(net563),
    .X(net568));
 sky130_fd_sc_hd__and2_1 c552 (.A(net941),
    .B(net564),
    .X(net569));
 sky130_fd_sc_hd__sdfxtp_1 c553 (.CLK(clknet_leaf_10_clk),
    .D(net565),
    .SCD(net569),
    .SCE(net941),
    .Q(net570));
 sky130_fd_sc_hd__clkbuf_1 c554 (.A(net749),
    .X(net571));
 sky130_fd_sc_hd__clkbuf_1 c555 (.A(net970),
    .X(net572));
 sky130_fd_sc_hd__and2_0 c556 (.A(net570),
    .B(net567),
    .X(net573));
 sky130_fd_sc_hd__sdfxtp_1 c557 (.CLK(clknet_leaf_10_clk),
    .D(net572),
    .SCD(clknet_1_0__leaf_net566),
    .SCE(net564),
    .Q(net574));
 sky130_fd_sc_hd__mux4_1 c558 (.A0(net906),
    .A1(clknet_1_1__leaf_net566),
    .A2(net457),
    .A3(net567),
    .S0(net553),
    .S1(net563),
    .X(net575));
 sky130_fd_sc_hd__and3_2 c559 (.A(net551),
    .B(net924),
    .C(net564),
    .X(net576));
 sky130_fd_sc_hd__and3_1 c56 (.A(net25),
    .B(net966),
    .C(net28),
    .X(net37));
 sky130_fd_sc_hd__dfbbn_1 c560 (.CLK_N(clknet_leaf_10_clk),
    .D(net571),
    .RESET_B(net569),
    .SET_B(net576),
    .Q(net577));
 sky130_fd_sc_hd__dfbbn_1 c561 (.CLK_N(clknet_leaf_18_clk),
    .D(net897),
    .RESET_B(net576),
    .SET_B(net439),
    .Q(net579),
    .Q_N(net578));
 sky130_fd_sc_hd__dfbbp_1 c562 (.CLK(clknet_leaf_18_clk),
    .D(clknet_1_1__leaf_net566),
    .RESET_B(net578),
    .SET_B(net576),
    .Q(net580));
 sky130_fd_sc_hd__sdfxbp_1 c563 (.CLK(clknet_leaf_10_clk),
    .D(net579),
    .SCD(net906),
    .SCE(net576),
    .Q(net582),
    .Q_N(net581));
 sky130_fd_sc_hd__sdfxbp_1 c564 (.CLK(clknet_leaf_10_clk),
    .D(net842),
    .SCD(net563),
    .SCE(net569),
    .Q(net583));
 sky130_fd_sc_hd__and3_1 c565 (.A(net553),
    .B(net842),
    .C(net579),
    .X(net584));
 sky130_fd_sc_hd__sdfbbp_1 c566 (.CLK(clknet_leaf_10_clk),
    .D(net898),
    .RESET_B(net584),
    .SCD(net947),
    .SCE(net941),
    .SET_B(clknet_1_1__leaf_net566),
    .Q(net586),
    .Q_N(net585));
 sky130_fd_sc_hd__clkbuf_1 c567 (.A(net477),
    .X(net587));
 sky130_fd_sc_hd__buf_1 c568 (.A(net759),
    .X(net588));
 sky130_fd_sc_hd__and2_0 c569 (.A(net573),
    .B(net466),
    .X(net589));
 sky130_fd_sc_hd__sdfxtp_1 c57 (.CLK(clknet_leaf_36_clk),
    .D(net37),
    .SCD(net919),
    .SCE(net21),
    .Q(net38));
 sky130_fd_sc_hd__and2_0 c570 (.A(net589),
    .B(net553),
    .X(net590));
 sky130_fd_sc_hd__and2_0 c571 (.A(net588),
    .B(net465),
    .X(net591));
 sky130_fd_sc_hd__and2_1 c572 (.A(net591),
    .B(net588),
    .X(net592));
 sky130_fd_sc_hd__and2_0 c573 (.A(net465),
    .B(net589),
    .X(net593));
 sky130_fd_sc_hd__clkbuf_1 c574 (.A(net758),
    .X(net594));
 sky130_fd_sc_hd__dfstp_1 c575 (.CLK(clknet_leaf_17_clk),
    .D(net594),
    .SET_B(net592),
    .Q(net595));
 sky130_fd_sc_hd__dfstp_1 c576 (.CLK(clknet_leaf_17_clk),
    .D(net859),
    .SET_B(net592),
    .Q(net838));
 sky130_fd_sc_hd__dlrbn_1 c577 (.D(net587),
    .GATE_N(clknet_leaf_17_clk),
    .RESET_B(net859),
    .Q(net597),
    .Q_N(net596));
 sky130_fd_sc_hd__dlrbn_1 c578 (.D(net590),
    .GATE_N(clknet_leaf_18_clk),
    .RESET_B(net588),
    .Q(net598));
 sky130_fd_sc_hd__sdfxtp_1 c579 (.CLK(clknet_leaf_18_clk),
    .D(net598),
    .SCD(net596),
    .SCE(net576),
    .Q(net599));
 sky130_fd_sc_hd__and3_1 c58 (.A(net24),
    .B(net26),
    .C(net29),
    .X(net39));
 sky130_fd_sc_hd__and2_0 c580 (.A(net457),
    .B(net599),
    .X(net600));
 sky130_fd_sc_hd__sdfrtp_1 c581 (.CLK(clknet_leaf_18_clk),
    .D(net597),
    .RESET_B(net592),
    .SCD(net594),
    .SCE(net599),
    .Q(net601));
 sky130_fd_sc_hd__and2_2 c582 (.A(net589),
    .B(net909),
    .X(net602));
 sky130_fd_sc_hd__sdfxtp_1 c583 (.CLK(clknet_leaf_18_clk),
    .D(net564),
    .SCD(net944),
    .SCE(net602),
    .Q(net603));
 sky130_fd_sc_hd__sdfrtp_1 c584 (.CLK(clknet_leaf_18_clk),
    .D(net883),
    .RESET_B(net597),
    .SCD(net600),
    .SCE(net602),
    .Q(net828));
 sky130_fd_sc_hd__sdfrtp_1 c585 (.CLK(clknet_leaf_18_clk),
    .D(net600),
    .RESET_B(net859),
    .SCD(net602),
    .SCE(net592),
    .Q(net604));
 sky130_fd_sc_hd__and2_0 c586 (.A(net599),
    .B(net604),
    .X(net605));
 sky130_fd_sc_hd__and2_0 c587 (.A(net968),
    .B(net605),
    .X(net606));
 sky130_fd_sc_hd__buf_1 c588 (.A(net763),
    .X(net607));
 sky130_fd_sc_hd__buf_1 c589 (.A(net498),
    .X(net608));
 sky130_fd_sc_hd__and3_1 c59 (.A(net38),
    .B(net36),
    .C(net39),
    .X(net40));
 sky130_fd_sc_hd__buf_1 c590 (.A(net607),
    .X(net609));
 sky130_fd_sc_hd__clkbuf_1 c591 (.A(net762),
    .X(net610));
 sky130_fd_sc_hd__and2_1 c592 (.A(net608),
    .B(net610),
    .X(net611));
 sky130_fd_sc_hd__and2_0 c593 (.A(net611),
    .B(net609),
    .X(net612));
 sky130_fd_sc_hd__and2_0 c594 (.A(net580),
    .B(net609),
    .X(net613));
 sky130_fd_sc_hd__and2_1 c595 (.A(net611),
    .B(net613),
    .X(net614));
 sky130_fd_sc_hd__and2_0 c596 (.A(net613),
    .B(net608),
    .X(net615));
 sky130_fd_sc_hd__sdfxtp_1 c597 (.CLK(clknet_leaf_22_clk),
    .D(net612),
    .SCD(net609),
    .SCE(net614),
    .Q(net616));
 sky130_fd_sc_hd__dlrbp_1 c598 (.D(net614),
    .GATE(clknet_leaf_22_clk),
    .RESET_B(net616),
    .Q(net618),
    .Q_N(net617));
 sky130_fd_sc_hd__and2_1 c599 (.A(net608),
    .B(net611),
    .X(net821));
 sky130_fd_sc_hd__mux4_1 c60 (.A0(net36),
    .A1(net39),
    .A2(net33),
    .A3(net20),
    .S0(net31),
    .S1(net22),
    .X(net41));
 sky130_fd_sc_hd__dlrbp_1 c600 (.D(net615),
    .GATE(clknet_leaf_17_clk),
    .RESET_B(net607),
    .Q(net620),
    .Q_N(net619));
 sky130_fd_sc_hd__dfbbn_1 c601 (.CLK_N(clknet_leaf_22_clk),
    .D(net610),
    .RESET_B(net614),
    .SET_B(net616),
    .Q(net622),
    .Q_N(net621));
 sky130_fd_sc_hd__dfbbn_1 c602 (.CLK_N(clknet_leaf_23_clk),
    .D(net616),
    .RESET_B(net921),
    .SET_B(net840),
    .Q(net623));
 sky130_fd_sc_hd__dfbbp_1 c603 (.CLK(clknet_leaf_23_clk),
    .D(net885),
    .RESET_B(net623),
    .SET_B(net840),
    .Q(net625),
    .Q_N(net624));
 sky130_fd_sc_hd__sdfxbp_1 c604 (.CLK(clknet_leaf_22_clk),
    .D(net879),
    .SCD(net625),
    .SCE(net840),
    .Q(net626));
 sky130_fd_sc_hd__and3_1 c605 (.A(net609),
    .B(net626),
    .C(net624),
    .X(net627));
 sky130_fd_sc_hd__mux4_1 c606 (.A0(net627),
    .A1(net617),
    .A2(net625),
    .A3(net611),
    .S0(net607),
    .S1(net840),
    .X(net628));
 sky130_fd_sc_hd__sdfbbn_1 c607 (.CLK_N(clknet_leaf_22_clk),
    .D(net911),
    .RESET_B(net616),
    .SCD(net624),
    .SCE(net840),
    .SET_B(net791),
    .Q(net629));
 sky130_fd_sc_hd__sdfsbp_1 c608 (.CLK(clknet_leaf_16_clk),
    .D(net607),
    .SCD(net629),
    .SCE(net942),
    .SET_B(net840),
    .Q(net630),
    .Q_N(net822));
 sky130_fd_sc_hd__and3_1 c61 (.A(net32),
    .B(net34),
    .C(net776),
    .X(net42));
 sky130_fd_sc_hd__sdfbbn_1 c62 (.CLK_N(clknet_leaf_37_clk),
    .D(net42),
    .RESET_B(net35),
    .SCD(net33),
    .SCE(net39),
    .SET_B(net22),
    .Q(net43));
 sky130_fd_sc_hd__buf_1 c63 (.A(net46),
    .X(net44));
 sky130_fd_sc_hd__buf_1 c630 (.A(net540),
    .X(net631));
 sky130_fd_sc_hd__buf_1 c631 (.X(net632));
 sky130_fd_sc_hd__clkbuf_1 c632 (.A(net757),
    .X(net633));
 sky130_fd_sc_hd__and2_0 c633 (.A(net633),
    .B(net540),
    .X(net634));
 sky130_fd_sc_hd__dlrtn_1 c634 (.D(net634),
    .GATE_N(clknet_leaf_6_clk),
    .RESET_B(net633),
    .Q(net635));
 sky130_fd_sc_hd__and2_0 c635 (.A(net633),
    .B(net632),
    .X(net636));
 sky130_fd_sc_hd__and2_1 c636 (.A(net912),
    .B(net635),
    .X(net637));
 sky130_fd_sc_hd__dlrtn_1 c637 (.D(net631),
    .GATE_N(clknet_leaf_12_clk),
    .RESET_B(net540),
    .Q(net638));
 sky130_fd_sc_hd__and2_0 c638 (.A(clknet_1_1__leaf_net521),
    .B(net632),
    .X(net639));
 sky130_fd_sc_hd__and2_0 c639 (.A(net639),
    .B(net635),
    .X(net640));
 sky130_fd_sc_hd__clkbuf_1 c64 (.A(net46),
    .X(net45));
 sky130_fd_sc_hd__sdfxbp_1 c640 (.CLK(clknet_leaf_6_clk),
    .D(net637),
    .SCD(net631),
    .SCE(clknet_1_0__leaf_net640),
    .Q(net642),
    .Q_N(net641));
 sky130_fd_sc_hd__dlrtn_1 c641 (.D(net915),
    .GATE_N(clknet_leaf_11_clk),
    .RESET_B(clknet_1_0__leaf_net640),
    .Q(net643));
 sky130_fd_sc_hd__and3_1 c642 (.A(net635),
    .B(net636),
    .C(net643),
    .X(net644));
 sky130_fd_sc_hd__sdfxtp_1 c643 (.CLK(clknet_leaf_6_clk),
    .D(net634),
    .SCD(net637),
    .SCE(clknet_1_1__leaf_net521),
    .Q(net645));
 sky130_fd_sc_hd__or4bb_1 c644 (.A(net636),
    .B(net644),
    .C_N(net540),
    .D_N(net889),
    .X(net646));
 sky130_fd_sc_hd__sdfbbn_1 c645 (.CLK_N(clknet_leaf_12_clk),
    .D(net644),
    .RESET_B(net646),
    .SCD(net638),
    .SCE(net641),
    .SET_B(net637),
    .Q(net647));
 sky130_fd_sc_hd__and3_1 c646 (.A(net632),
    .B(net643),
    .C(net641),
    .X(net648));
 sky130_fd_sc_hd__and3_1 c647 (.A(net648),
    .B(net644),
    .C(net642),
    .X(net649));
 sky130_fd_sc_hd__sdfxtp_1 c648 (.CLK(clknet_leaf_12_clk),
    .D(net876),
    .SCD(net649),
    .SCE(net644),
    .Q(net650));
 sky130_fd_sc_hd__sdfbbp_1 c649 (.CLK(clknet_leaf_12_clk),
    .D(net881),
    .RESET_B(net647),
    .SCD(net649),
    .SCE(net648),
    .SET_B(net637),
    .Q(net651));
 sky130_fd_sc_hd__buf_1 c65 (.A(net767),
    .X(net46));
 sky130_fd_sc_hd__sdfbbn_1 c650 (.CLK_N(clknet_leaf_12_clk),
    .D(net651),
    .RESET_B(clknet_1_1__leaf_net640),
    .SCD(net648),
    .SCE(net649),
    .SET_B(net638),
    .Q(net653),
    .Q_N(net652));
 sky130_fd_sc_hd__and2_0 c651 (.A(net653),
    .B(net553),
    .X(net654));
 sky130_fd_sc_hd__buf_2 c652 (.A(net773),
    .X(net655));
 sky130_fd_sc_hd__dlymetal6s2s_1 c653 (.A(net772),
    .X(net656));
 sky130_fd_sc_hd__and2_0 c654 (.A(net655),
    .B(net656),
    .X(net657));
 sky130_fd_sc_hd__and2_0 c655 (.A(net655),
    .B(net978),
    .X(net658));
 sky130_fd_sc_hd__dlrtp_1 c656 (.D(net656),
    .GATE(clknet_leaf_11_clk),
    .RESET_B(net654),
    .Q(net659));
 sky130_fd_sc_hd__and2_1 c657 (.A(net657),
    .B(net655),
    .X(net660));
 sky130_fd_sc_hd__dlrtp_1 c658 (.D(net649),
    .GATE(clknet_leaf_12_clk),
    .RESET_B(net656),
    .Q(net661));
 sky130_fd_sc_hd__and2_1 c659 (.A(net661),
    .B(net660),
    .X(net662));
 sky130_fd_sc_hd__clkbuf_1 c66 (.A(net46),
    .X(net47));
 sky130_fd_sc_hd__sdfxtp_1 c660 (.CLK(clknet_leaf_11_clk),
    .D(net662),
    .SCD(net657),
    .SCE(net655),
    .Q(net663));
 sky130_fd_sc_hd__dfbbn_1 c661 (.CLK_N(clknet_leaf_11_clk),
    .D(net556),
    .RESET_B(net662),
    .SET_B(net660),
    .Q(net664));
 sky130_fd_sc_hd__and3_1 c662 (.A(net660),
    .B(net655),
    .C(net663),
    .X(net665));
 sky130_fd_sc_hd__dfbbn_1 c663 (.CLK_N(clknet_leaf_11_clk),
    .D(net658),
    .RESET_B(net665),
    .SET_B(net662),
    .Q(net667),
    .Q_N(net666));
 sky130_fd_sc_hd__dfbbp_1 c664 (.CLK(clknet_leaf_11_clk),
    .D(net562),
    .RESET_B(net665),
    .SET_B(net666),
    .Q(net669),
    .Q_N(net668));
 sky130_fd_sc_hd__and3_1 c665 (.A(net669),
    .B(net667),
    .C(net663),
    .X(net670));
 sky130_fd_sc_hd__a2111o_1 c666 (.A1(net659),
    .A2(net669),
    .B1(net652),
    .C1(net670),
    .D1(net655),
    .X(net671));
 sky130_fd_sc_hd__and3_1 c667 (.A(net638),
    .B(net667),
    .C(net668),
    .X(net672));
 sky130_fd_sc_hd__and3_1 c668 (.A(net663),
    .B(net671),
    .C(net661),
    .X(net673));
 sky130_fd_sc_hd__sdfbbn_1 c669 (.CLK_N(clknet_leaf_12_clk),
    .D(net673),
    .RESET_B(net961),
    .SCD(net661),
    .SCE(net656),
    .SET_B(net655),
    .Q(net674));
 sky130_fd_sc_hd__buf_2 c67 (.A(net47),
    .X(net48));
 sky130_fd_sc_hd__mux4_1 c670 (.A0(net664),
    .A1(net670),
    .A2(net665),
    .A3(net659),
    .S0(net655),
    .S1(net668),
    .X(net675));
 sky130_fd_sc_hd__sdfbbp_1 c671 (.CLK(clknet_leaf_13_clk),
    .D(net674),
    .RESET_B(net666),
    .SCD(net673),
    .SCE(net655),
    .SET_B(net856),
    .Q(net676));
 sky130_fd_sc_hd__clkbuf_1 c672 (.A(net586),
    .X(net677));
 sky130_fd_sc_hd__buf_1 c673 (.A(net677),
    .X(net678));
 sky130_fd_sc_hd__and2_0 c674 (.A(net676),
    .B(net585),
    .X(net679));
 sky130_fd_sc_hd__clkbuf_1 c675 (.A(net656),
    .X(net680));
 sky130_fd_sc_hd__buf_1 c676 (.A(net680),
    .X(net681));
 sky130_fd_sc_hd__and2_2 c677 (.A(net678),
    .B(net680),
    .X(net682));
 sky130_fd_sc_hd__buf_1 c678 (.A(net769),
    .X(net683));
 sky130_fd_sc_hd__buf_1 c679 (.A(net768),
    .X(net684));
 sky130_fd_sc_hd__clkbuf_1 c68 (.A(net48),
    .X(net49));
 sky130_fd_sc_hd__dlrtp_1 c680 (.D(net681),
    .GATE(clknet_leaf_13_clk),
    .RESET_B(net682),
    .Q(net685));
 sky130_fd_sc_hd__and3_1 c681 (.A(net681),
    .B(net684),
    .C(net790),
    .X(net686));
 sky130_fd_sc_hd__edfxbp_1 c682 (.CLK(clknet_leaf_13_clk),
    .D(net682),
    .DE(net686),
    .Q(net687));
 sky130_fd_sc_hd__and2_0 c683 (.A(net677),
    .B(net684),
    .X(net688));
 sky130_fd_sc_hd__sdfxbp_1 c684 (.CLK(clknet_leaf_13_clk),
    .D(net683),
    .SCD(net682),
    .SCE(net684),
    .Q(net690),
    .Q_N(net689));
 sky130_fd_sc_hd__or4bb_1 c685 (.A(net679),
    .B(net681),
    .C_N(net678),
    .D_N(net683),
    .X(net691));
 sky130_fd_sc_hd__sdfxbp_1 c686 (.CLK(clknet_leaf_13_clk),
    .D(net895),
    .SCD(net691),
    .SCE(net586),
    .Q(net692));
 sky130_fd_sc_hd__or4bb_1 c687 (.A(net972),
    .B(net683),
    .C_N(net685),
    .D_N(net678),
    .X(net693));
 sky130_fd_sc_hd__sdfxtp_1 c688 (.CLK(clknet_leaf_13_clk),
    .D(net684),
    .SCD(net693),
    .SCE(net683),
    .Q(net694));
 sky130_fd_sc_hd__edfxtp_1 c689 (.CLK(clknet_leaf_13_clk),
    .D(net693),
    .DE(net682),
    .Q(net695));
 sky130_fd_sc_hd__and2_1 c69 (.A(net43),
    .B(net48),
    .X(net50));
 sky130_fd_sc_hd__sdfxtp_1 c690 (.CLK(clknet_leaf_14_clk),
    .D(net688),
    .SCD(net691),
    .SCE(net925),
    .Q(net696));
 sky130_fd_sc_hd__sdfbbn_1 c691 (.CLK_N(clknet_leaf_13_clk),
    .D(net694),
    .RESET_B(net695),
    .SCD(net689),
    .SCE(net678),
    .SET_B(net682),
    .Q(net697));
 sky130_fd_sc_hd__or4bb_1 c692 (.A(net687),
    .B(net697),
    .C_N(net683),
    .D_N(net694),
    .X(net698));
 sky130_fd_sc_hd__buf_1 c693 (.A(net744),
    .X(net699));
 sky130_fd_sc_hd__clkbuf_1 c694 (.A(net743),
    .X(net700));
 sky130_fd_sc_hd__and2_2 c695 (.A(net828),
    .B(net699),
    .X(net701));
 sky130_fd_sc_hd__and2_0 c696 (.A(net696),
    .B(net701),
    .X(net702));
 sky130_fd_sc_hd__and2_1 c697 (.A(net702),
    .B(net700),
    .X(net703));
 sky130_fd_sc_hd__and2_0 c698 (.A(net460),
    .B(net701),
    .X(net704));
 sky130_fd_sc_hd__and2_1 c699 (.A(net699),
    .B(net701),
    .X(net705));
 sky130_fd_sc_hd__buf_1 c70 (.A(net766),
    .X(net51));
 sky130_fd_sc_hd__sdfxtp_1 c700 (.CLK(clknet_leaf_15_clk),
    .D(net703),
    .SCD(net704),
    .SCE(net701),
    .Q(net706));
 sky130_fd_sc_hd__and2_0 c701 (.A(net706),
    .B(net699),
    .X(net707));
 sky130_fd_sc_hd__and2_4 c702 (.A(net698),
    .B(net705),
    .X(net708));
 sky130_fd_sc_hd__sdlclkp_1 c703 (.CLK(clknet_leaf_14_clk),
    .GATE(net686),
    .SCE(net708),
    .GCLK(net709));
 sky130_fd_sc_hd__a2111o_1 c704 (.A1(net702),
    .A2(net699),
    .B1(net707),
    .C1(clknet_1_0__leaf_net709),
    .D1(net701),
    .X(net710));
 sky130_fd_sc_hd__dfbbn_1 c705 (.CLK_N(clknet_leaf_14_clk),
    .D(net701),
    .RESET_B(clknet_1_1__leaf_net709),
    .SET_B(net708),
    .Q(net712),
    .Q_N(net711));
 sky130_fd_sc_hd__mux4_1 c706 (.A0(net712),
    .A1(clknet_1_1__leaf_net709),
    .A2(net705),
    .A3(net703),
    .S0(clknet_1_1__leaf_net710),
    .S1(net701),
    .X(net713));
 sky130_fd_sc_hd__and3_1 c707 (.A(net712),
    .B(clknet_1_1__leaf_net709),
    .C(net793),
    .X(net714));
 sky130_fd_sc_hd__dfbbn_1 c708 (.CLK_N(clknet_leaf_15_clk),
    .D(net708),
    .RESET_B(clknet_1_0__leaf_net709),
    .SET_B(net706),
    .Q(net716),
    .Q_N(net715));
 sky130_fd_sc_hd__and3_1 c709 (.A(net704),
    .B(net707),
    .C(net715),
    .X(net717));
 sky130_fd_sc_hd__and3_1 c71 (.A(net51),
    .B(net48),
    .C(net47),
    .X(net52));
 sky130_fd_sc_hd__dfbbp_1 c710 (.CLK(clknet_leaf_14_clk),
    .D(clknet_1_1__leaf_net714),
    .RESET_B(clknet_1_0__leaf_net710),
    .SET_B(clknet_1_1__leaf_net709),
    .Q(net718));
 sky130_fd_sc_hd__mux4_1 c711 (.A0(net692),
    .A1(net718),
    .A2(clknet_1_0__leaf_net710),
    .A3(net711),
    .S0(net701),
    .S1(net703),
    .X(net719));
 sky130_fd_sc_hd__mux4_1 c712 (.A0(net700),
    .A1(net717),
    .A2(clknet_1_0__leaf_net714),
    .A3(net705),
    .S0(net701),
    .S1(clknet_1_0__leaf_net794),
    .X(net720));
 sky130_fd_sc_hd__and3_1 c713 (.A(net716),
    .B(clknet_1_1__leaf_net794),
    .C(net795),
    .X(net721));
 sky130_fd_sc_hd__sdfxbp_1 c714 (.CLK(clknet_leaf_16_clk),
    .D(net934),
    .SCD(clknet_1_1__leaf_net721),
    .SCE(net840),
    .Q(net723),
    .Q_N(net722));
 sky130_fd_sc_hd__sdlclkp_2 c715 (.CLK(clknet_leaf_15_clk),
    .GATE(net896),
    .SCE(net703),
    .GCLK(net724));
 sky130_fd_sc_hd__and2_0 c716 (.A(clknet_1_0__leaf_net724),
    .B(net722),
    .X(net725));
 sky130_fd_sc_hd__and3_1 c717 (.A(clknet_1_0__leaf_net709),
    .B(net896),
    .C(clknet_1_0__leaf_net725),
    .X(net726));
 sky130_fd_sc_hd__and2_0 c718 (.A(clknet_1_0__leaf_net725),
    .B(clknet_1_1__leaf_net726),
    .X(net727));
 sky130_fd_sc_hd__sdfxbp_1 c719 (.CLK(clknet_leaf_16_clk),
    .D(clknet_1_1__leaf_net724),
    .SCD(clknet_1_1__leaf_net727),
    .SCE(clknet_1_1__leaf_net725),
    .Q(net729),
    .Q_N(net728));
 sky130_fd_sc_hd__sdfxtp_1 c72 (.CLK(clknet_leaf_0_clk),
    .D(net52),
    .SCD(net51),
    .SCE(net48),
    .Q(net53));
 sky130_fd_sc_hd__and3_1 c720 (.A(net896),
    .B(clknet_1_0__leaf_net721),
    .C(net728),
    .X(net730));
 sky130_fd_sc_hd__sdfxtp_1 c721 (.CLK(clknet_leaf_15_clk),
    .D(net703),
    .SCD(net886),
    .SCE(clknet_1_0__leaf_net727),
    .Q(net731));
 sky130_fd_sc_hd__sdfxtp_1 c722 (.CLK(clknet_leaf_15_clk),
    .D(net886),
    .SCD(clknet_1_1__leaf_net730),
    .SCE(net840),
    .Q(net732));
 sky130_fd_sc_hd__and3_1 c723 (.A(clknet_1_0__leaf_net730),
    .B(net732),
    .C(clknet_1_0__leaf_net726),
    .X(net733));
 sky130_fd_sc_hd__mux4_1 c724 (.A0(clknet_1_0__leaf_net724),
    .A1(net731),
    .A2(clknet_1_1__leaf_net727),
    .A3(net722),
    .S0(clknet_1_0__leaf_net733),
    .S1(clknet_1_0__leaf_net709),
    .X(net734));
 sky130_fd_sc_hd__sdfxtp_1 c725 (.CLK(clknet_leaf_17_clk),
    .D(clknet_1_0__leaf_net726),
    .SCD(net946),
    .SCE(net840),
    .Q(net735));
 sky130_fd_sc_hd__dfbbn_1 c726 (.CLK_N(clknet_leaf_17_clk),
    .D(clknet_1_0__leaf_net733),
    .RESET_B(clknet_1_0__leaf_net727),
    .SET_B(clknet_1_0__leaf_net730),
    .Q(net737),
    .Q_N(net736));
 sky130_fd_sc_hd__and3_1 c727 (.A(net735),
    .B(net736),
    .C(net796),
    .X(net738));
 sky130_fd_sc_hd__and3_1 c728 (.A(net732),
    .B(net737),
    .C(net738),
    .X(net739));
 sky130_fd_sc_hd__and3_1 c729 (.A(net737),
    .B(net738),
    .C(net739),
    .X(net740));
 sky130_fd_sc_hd__dfrtp_1 c73 (.CLK(clknet_leaf_35_clk),
    .D(net45),
    .RESET_B(net50),
    .Q(net54));
 sky130_fd_sc_hd__mux4_1 c730 (.A0(clknet_1_0__leaf_net727),
    .A1(net739),
    .A2(net735),
    .A3(net821),
    .S0(net732),
    .S1(net740),
    .X(net741));
 sky130_fd_sc_hd__mux4_1 c731 (.A0(net740),
    .A1(net738),
    .A2(net739),
    .A3(clknet_1_1__leaf_net733),
    .S0(net821),
    .S1(net797),
    .X(net742));
 sky130_fd_sc_hd__dfrtp_1 c74 (.CLK(clknet_leaf_35_clk),
    .D(net49),
    .RESET_B(net45),
    .Q(net55));
 sky130_fd_sc_hd__and2_0 c75 (.A(net851),
    .B(net951),
    .X(net56));
 sky130_fd_sc_hd__or4bb_2 c76 (.A(net47),
    .B(net851),
    .C_N(net54),
    .D_N(net48),
    .X(net57));
 sky130_fd_sc_hd__dfrtp_1 c77 (.CLK(clknet_leaf_31_clk),
    .D(net56),
    .RESET_B(net852),
    .Q(net58));
 sky130_fd_sc_hd__sdfxtp_1 c78 (.CLK(clknet_leaf_34_clk),
    .D(net57),
    .SCD(net50),
    .SCE(net51),
    .Q(net59));
 sky130_fd_sc_hd__dfsbp_1 c79 (.CLK(clknet_leaf_34_clk),
    .D(net50),
    .SET_B(net854),
    .Q(net61),
    .Q_N(net60));
 sky130_fd_sc_hd__and3_1 c80 (.A(net51),
    .B(net60),
    .C(net48),
    .X(net62));
 sky130_fd_sc_hd__dfbbn_1 c81 (.CLK_N(clknet_leaf_37_clk),
    .D(net54),
    .RESET_B(net53),
    .SET_B(net52),
    .Q(net64),
    .Q_N(net63));
 sky130_fd_sc_hd__mux4_1 c82 (.A0(net44),
    .A1(net61),
    .A2(net56),
    .A3(net63),
    .S0(net48),
    .S1(net30),
    .X(net65));
 sky130_fd_sc_hd__mux4_1 c83 (.A0(net971),
    .A1(net62),
    .A2(net64),
    .A3(net65),
    .S0(net48),
    .S1(net57),
    .X(net66));
 sky130_fd_sc_hd__buf_1 c84 (.A(net866),
    .X(net67));
 sky130_fd_sc_hd__buf_1 c85 (.A(net67),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_1 c86 (.A(net68),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_1 c87 (.A(net68),
    .X(net70));
 sky130_fd_sc_hd__buf_1 c88 (.A(net857),
    .X(net71));
 sky130_fd_sc_hd__clkbuf_2 c89 (.A(net849),
    .X(net72));
 sky130_fd_sc_hd__and2_1 c90 (.A(net68),
    .B(net72),
    .X(net73));
 sky130_fd_sc_hd__and2_1 c91 (.A(net68),
    .B(net72),
    .X(net74));
 sky130_fd_sc_hd__and2_1 c92 (.A(net71),
    .B(net72),
    .X(net75));
 sky130_fd_sc_hd__sdfrbp_1 c93 (.CLK(clknet_leaf_31_clk),
    .D(net73),
    .RESET_B(net71),
    .SCD(net74),
    .SCE(net72),
    .Q(net76));
 sky130_fd_sc_hd__dfsbp_1 c94 (.CLK(clknet_leaf_33_clk),
    .D(net69),
    .SET_B(net74),
    .Q(net77));
 sky130_fd_sc_hd__and2_0 c95 (.A(net77),
    .B(net71),
    .X(net78));
 sky130_fd_sc_hd__dfstp_1 c96 (.CLK(clknet_leaf_32_clk),
    .D(net74),
    .SET_B(net75),
    .Q(net79));
 sky130_fd_sc_hd__dfbbn_1 c97 (.CLK_N(clknet_leaf_31_clk),
    .D(net72),
    .RESET_B(net70),
    .SET_B(net74),
    .Q(net81),
    .Q_N(net80));
 sky130_fd_sc_hd__dfbbp_1 c98 (.CLK(clknet_leaf_31_clk),
    .D(net81),
    .RESET_B(net79),
    .SET_B(net74),
    .Q(net83),
    .Q_N(net82));
 sky130_fd_sc_hd__and3_1 c99 (.A(net76),
    .B(net72),
    .C(net71),
    .X(net84));
 sky130_fd_sc_hd__sdfsbp_1 merge732 (.CLK(clknet_leaf_15_clk),
    .D(net606),
    .SCD(net686),
    .SCE(net472),
    .SET_B(net602),
    .Q(net744),
    .Q_N(net743));
 sky130_fd_sc_hd__dfbbn_1 merge733 (.CLK_N(clknet_leaf_36_clk),
    .D(net20),
    .RESET_B(net22),
    .Q(net23),
    .Q_N(net745));
 sky130_fd_sc_hd__dfxtp_1 merge734 (.CLK(clknet_leaf_3_clk),
    .D(net135),
    .Q(net747));
 sky130_fd_sc_hd__dfbbp_1 merge735 (.CLK(clknet_leaf_10_clk),
    .D(clknet_1_0__leaf_net566),
    .RESET_B(net941),
    .SET_B(net569),
    .Q(net749),
    .Q_N(net748));
 sky130_fd_sc_hd__sdfxbp_1 merge736 (.CLK(clknet_leaf_34_clk),
    .D(net69),
    .SCD(net70),
    .SCE(net67),
    .Q(net751),
    .Q_N(net750));
 sky130_fd_sc_hd__sdfxbp_1 merge737 (.CLK(clknet_leaf_4_clk),
    .D(net246),
    .SCD(net127),
    .Q(net247),
    .Q_N(net752));
 sky130_fd_sc_hd__sdfstp_1 merge738 (.CLK(clknet_leaf_24_clk),
    .D(net369),
    .SCD(net370),
    .SCE(net948),
    .SET_B(net373),
    .Q(net754));
 sky130_fd_sc_hd__sdfxtp_1 merge739 (.CLK(clknet_leaf_20_clk),
    .D(net441),
    .SCD(clknet_1_0__leaf_net318),
    .SCE(net301),
    .Q(net755));
 sky130_fd_sc_hd__sdfxtp_1 merge740 (.CLK(clknet_leaf_8_clk),
    .D(net295),
    .SCD(net402),
    .SCE(net409),
    .Q(net756));
 sky130_fd_sc_hd__sdfxtp_1 merge741 (.CLK(clknet_leaf_6_clk),
    .D(net631),
    .SCD(net540),
    .Q(net632));
 sky130_fd_sc_hd__dfbbn_1 merge742 (.CLK_N(clknet_leaf_18_clk),
    .D(net576),
    .RESET_B(net564),
    .SET_B(net593),
    .Q(net759),
    .Q_N(net758));
 sky130_fd_sc_hd__sdfstp_1 merge743 (.CLK(clknet_leaf_0_clk),
    .D(net159),
    .SCD(net160),
    .SCE(net168),
    .SET_B(net853),
    .Q(net760));
 sky130_fd_sc_hd__sdlclkp_4 merge744 (.CLK(clknet_leaf_33_clk),
    .GATE(net94),
    .SCE(net93),
    .GCLK(net761));
 sky130_fd_sc_hd__dfrbp_1 merge745 (.CLK(clknet_leaf_17_clk),
    .D(net602),
    .RESET_B(net848),
    .Q(net763),
    .Q_N(net762));
 sky130_fd_sc_hd__dfrbp_1 merge746 (.CLK(clknet_leaf_18_clk),
    .D(net463),
    .RESET_B(net465),
    .Q(net765),
    .Q_N(net764));
 sky130_fd_sc_hd__dfbbn_1 merge747 (.CLK_N(clknet_leaf_35_clk),
    .D(net40),
    .RESET_B(net49),
    .SET_B(net44),
    .Q(net767),
    .Q_N(net766));
 sky130_fd_sc_hd__dfbbp_1 merge748 (.CLK(clknet_leaf_13_clk),
    .D(net568),
    .RESET_B(net682),
    .SET_B(net681),
    .Q(net769),
    .Q_N(net768));
 sky130_fd_sc_hd__dfrtn_1 merge749 (.CLK_N(clknet_leaf_32_clk),
    .D(net225),
    .RESET_B(net201),
    .Q(net770));
 sky130_fd_sc_hd__dfrtp_1 merge750 (.CLK(clknet_leaf_21_clk),
    .D(net342),
    .RESET_B(net489),
    .Q(net771));
 sky130_fd_sc_hd__sdfxbp_1 merge751 (.CLK(clknet_leaf_11_clk),
    .D(net654),
    .SCD(net553),
    .SCE(net643),
    .Q(net773),
    .Q_N(net772));
 sky130_fd_sc_hd__sdfxbp_1 merge752 (.CLK(clknet_leaf_7_clk),
    .D(clknet_1_0__leaf_net256),
    .SCD(net396),
    .SCE(net936),
    .Q(net775),
    .Q_N(net774));
 sky130_fd_sc_hd__dfxtp_1 s753 (.CLK(clknet_leaf_37_clk),
    .D(net41),
    .Q(net776));
 sky130_fd_sc_hd__dfxtp_1 s754 (.CLK(clknet_leaf_31_clk),
    .D(net66),
    .Q(net777));
 sky130_fd_sc_hd__dlclkp_1 s755 (.CLK(clknet_leaf_27_clk),
    .GATE(net110),
    .GCLK(net778));
 sky130_fd_sc_hd__dlclkp_2 s756 (.CLK(clknet_leaf_4_clk),
    .GATE(net134),
    .GCLK(net779));
 sky130_fd_sc_hd__dlclkp_4 s757 (.CLK(clknet_leaf_3_clk),
    .GATE(net150),
    .GCLK(net780));
 sky130_fd_sc_hd__dlxbn_1 s758 (.D(net177),
    .GATE_N(clknet_leaf_1_clk),
    .Q(net781));
 sky130_fd_sc_hd__dlxbn_1 s759 (.D(net270),
    .GATE_N(clknet_leaf_2_clk),
    .Q(net782));
 sky130_fd_sc_hd__dlxbp_1 s760 (.D(net294),
    .GATE(clknet_leaf_1_clk),
    .Q(net784),
    .Q_N(net783));
 sky130_fd_sc_hd__dlxtn_1 s761 (.D(net340),
    .GATE_N(clknet_leaf_21_clk),
    .Q(net785));
 sky130_fd_sc_hd__dlxtn_1 s762 (.D(net341),
    .GATE_N(clknet_leaf_20_clk),
    .Q(net786));
 sky130_fd_sc_hd__dlxtn_1 s763 (.D(net384),
    .GATE_N(clknet_leaf_24_clk),
    .Q(net787));
 sky130_fd_sc_hd__dlxtp_1 s764 (.D(net414),
    .GATE(clknet_leaf_8_clk),
    .Q(net788));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s765 (.D(net479),
    .SLEEP_B(clknet_leaf_21_clk),
    .Q(net789));
 sky130_fd_sc_hd__dfxbp_1 s766 (.CLK(clknet_leaf_23_clk),
    .D(net515),
    .Q(net824),
    .Q_N(net835));
 sky130_fd_sc_hd__dfxbp_1 s767 (.CLK(clknet_leaf_25_clk),
    .D(net517),
    .Q(net839),
    .Q_N(net830));
 sky130_fd_sc_hd__dfxtp_1 s768 (.CLK(clknet_leaf_18_clk),
    .D(net575),
    .Q(net790));
 sky130_fd_sc_hd__dfxtp_1 s769 (.CLK(clknet_leaf_23_clk),
    .D(net628),
    .Q(net791));
 sky130_fd_sc_hd__dfxtp_1 s770 (.CLK(clknet_leaf_13_clk),
    .D(net675),
    .Q(net792));
 sky130_fd_sc_hd__dlclkp_1 s771 (.CLK(clknet_leaf_14_clk),
    .GATE(net713),
    .GCLK(net793));
 sky130_fd_sc_hd__dlclkp_2 s772 (.CLK(clknet_leaf_14_clk),
    .GATE(net719),
    .GCLK(net794));
 sky130_fd_sc_hd__dlclkp_4 s773 (.CLK(clknet_leaf_15_clk),
    .GATE(net720),
    .GCLK(net795));
 sky130_fd_sc_hd__dlxbn_1 s774 (.D(net734),
    .GATE_N(clknet_leaf_16_clk),
    .Q(net796));
 sky130_fd_sc_hd__dlxbn_1 s775 (.D(net741),
    .GATE_N(clknet_leaf_16_clk),
    .Q(net797));
 sky130_fd_sc_hd__dlxbp_1 s776 (.D(net742),
    .GATE(clknet_leaf_16_clk));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Right_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Right_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Right_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Right_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Right_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Right_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Right_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Right_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Right_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Right_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Right_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Right_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Right_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Right_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Right_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Right_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Right_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Right_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Right_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Right_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Right_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_161 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_162 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_163 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_164 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_165 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_166 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_167 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_168 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_169 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_170 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_171 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_172 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_173 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_174 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_175 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_176 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_177 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_178 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_179 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_180 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_181 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_182 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Left_183 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Left_184 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Left_185 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Left_186 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Left_187 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Left_188 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Left_189 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Left_190 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Left_191 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Left_192 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Left_193 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Left_194 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Left_195 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Left_196 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Left_197 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Left_198 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Left_199 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Left_200 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Left_201 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Left_202 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Left_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1347 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(in0),
    .X(net746));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(in1),
    .X(net753));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(in10),
    .X(net798));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(in11),
    .X(net799));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(in12),
    .X(net800));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(in13),
    .X(net801));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(in15),
    .X(net802));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(in16),
    .X(net803));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(in17),
    .X(net804));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(in18),
    .X(net805));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(in19),
    .X(net806));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(in2),
    .X(net807));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(in20),
    .X(net808));
 sky130_fd_sc_hd__clkbuf_2 input14 (.A(in21),
    .X(net809));
 sky130_fd_sc_hd__clkbuf_2 input15 (.A(in22),
    .X(net810));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(in23),
    .X(net811));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(in24),
    .X(net812));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(in3),
    .X(net813));
 sky130_fd_sc_hd__clkbuf_1 input19 (.A(in4),
    .X(net814));
 sky130_fd_sc_hd__clkbuf_1 input20 (.A(in5),
    .X(net815));
 sky130_fd_sc_hd__clkbuf_1 input21 (.A(in6),
    .X(net816));
 sky130_fd_sc_hd__clkbuf_1 input22 (.A(in7),
    .X(net817));
 sky130_fd_sc_hd__clkbuf_1 input23 (.A(in8),
    .X(net818));
 sky130_fd_sc_hd__clkbuf_1 input24 (.A(in9),
    .X(net819));
 sky130_fd_sc_hd__buf_2 output25 (.A(net820),
    .X(out1));
 sky130_fd_sc_hd__buf_2 output26 (.A(net840),
    .X(out10));
 sky130_fd_sc_hd__buf_2 output27 (.A(net822),
    .X(out11));
 sky130_fd_sc_hd__buf_2 output28 (.A(net823),
    .X(out13));
 sky130_fd_sc_hd__buf_2 output29 (.A(net824),
    .X(out15));
 sky130_fd_sc_hd__buf_2 output30 (.A(net825),
    .X(out16));
 sky130_fd_sc_hd__buf_2 output31 (.A(net826),
    .X(out17));
 sky130_fd_sc_hd__buf_2 output32 (.A(net827),
    .X(out18));
 sky130_fd_sc_hd__buf_2 output33 (.A(net828),
    .X(out19));
 sky130_fd_sc_hd__buf_2 output34 (.A(net829),
    .X(out2));
 sky130_fd_sc_hd__buf_2 output35 (.A(net830),
    .X(out20));
 sky130_fd_sc_hd__buf_2 output36 (.A(net831),
    .X(out21));
 sky130_fd_sc_hd__buf_2 output37 (.A(net832),
    .X(out22));
 sky130_fd_sc_hd__buf_2 output38 (.A(net833),
    .X(out23));
 sky130_fd_sc_hd__buf_2 output39 (.A(net834),
    .X(out24));
 sky130_fd_sc_hd__buf_2 output40 (.A(net835),
    .X(out4));
 sky130_fd_sc_hd__buf_2 output41 (.A(net836),
    .X(out5));
 sky130_fd_sc_hd__buf_2 output42 (.A(net837),
    .X(out6));
 sky130_fd_sc_hd__buf_2 output43 (.A(net838),
    .X(out8));
 sky130_fd_sc_hd__buf_2 output44 (.A(net839),
    .X(out9));
 sky130_fd_sc_hd__clkbuf_4 fanout45 (.A(net821),
    .X(net840));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_0_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_1_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_2_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_3_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_4_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_5_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_6_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_7_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_8_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_9_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_9_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_10_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_11_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_12_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_13_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_14_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_15_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_16_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_17_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_18_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_19_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_20_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_21_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_22_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_22_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_23_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_24_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_24_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_25_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_25_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_26_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_26_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_27_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_27_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_28_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_28_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_29_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_29_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_30_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_30_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_31_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_31_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_32_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_32_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_33_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_33_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_34_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_34_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_35_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_35_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_36_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_36_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_37_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_37_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net721 (.A(net721),
    .X(clknet_0_net721));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net721 (.A(clknet_0_net721),
    .X(clknet_1_0__leaf_net721));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net721 (.A(clknet_0_net721),
    .X(clknet_1_1__leaf_net721));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net730 (.A(net730),
    .X(clknet_0_net730));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net730 (.A(clknet_0_net730),
    .X(clknet_1_0__leaf_net730));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net730 (.A(clknet_0_net730),
    .X(clknet_1_1__leaf_net730));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net733 (.A(net733),
    .X(clknet_0_net733));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net733 (.A(clknet_0_net733),
    .X(clknet_1_0__leaf_net733));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net733 (.A(clknet_0_net733),
    .X(clknet_1_1__leaf_net733));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net794 (.A(net794),
    .X(clknet_0_net794));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net794 (.A(clknet_0_net794),
    .X(clknet_1_0__leaf_net794));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net794 (.A(clknet_0_net794),
    .X(clknet_1_1__leaf_net794));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net714 (.A(net714),
    .X(clknet_0_net714));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net714 (.A(clknet_0_net714),
    .X(clknet_1_0__leaf_net714));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net714 (.A(clknet_0_net714),
    .X(clknet_1_1__leaf_net714));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net779 (.A(net779),
    .X(clknet_0_net779));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net779 (.A(clknet_0_net779),
    .X(clknet_1_0__leaf_net779));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net779 (.A(clknet_0_net779),
    .X(clknet_1_1__leaf_net779));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net278 (.A(net278),
    .X(clknet_0_net278));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net278 (.A(clknet_0_net278),
    .X(clknet_1_0__leaf_net278));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net278 (.A(clknet_0_net278),
    .X(clknet_1_1__leaf_net278));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net285 (.A(net285),
    .X(clknet_0_net285));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net285 (.A(clknet_0_net285),
    .X(clknet_1_0__leaf_net285));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net285 (.A(clknet_0_net285),
    .X(clknet_1_1__leaf_net285));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net284 (.A(net284),
    .X(clknet_0_net284));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net284 (.A(clknet_0_net284),
    .X(clknet_1_0__leaf_net284));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net284 (.A(clknet_0_net284),
    .X(clknet_1_1__leaf_net284));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net287 (.A(net287),
    .X(clknet_0_net287));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net287 (.A(clknet_0_net287),
    .X(clknet_1_0__leaf_net287));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net287 (.A(clknet_0_net287),
    .X(clknet_1_1__leaf_net287));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net248 (.A(net248),
    .X(clknet_0_net248));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net248 (.A(clknet_0_net248),
    .X(clknet_1_0__leaf_net248));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net248 (.A(clknet_0_net248),
    .X(clknet_1_1__leaf_net248));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net255 (.A(net255),
    .X(clknet_0_net255));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net255 (.A(clknet_0_net255),
    .X(clknet_1_0__leaf_net255));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net255 (.A(clknet_0_net255),
    .X(clknet_1_1__leaf_net255));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net256 (.A(net256),
    .X(clknet_0_net256));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net256 (.A(clknet_0_net256),
    .X(clknet_1_0__leaf_net256));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net256 (.A(clknet_0_net256),
    .X(clknet_1_1__leaf_net256));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net520 (.A(net520),
    .X(clknet_0_net520));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net520 (.A(clknet_0_net520),
    .X(clknet_1_0__leaf_net520));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net520 (.A(clknet_0_net520),
    .X(clknet_1_1__leaf_net520));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net523 (.A(net523),
    .X(clknet_0_net523));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net523 (.A(clknet_0_net523),
    .X(clknet_1_0__leaf_net523));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net523 (.A(clknet_0_net523),
    .X(clknet_1_1__leaf_net523));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net525 (.A(net525),
    .X(clknet_0_net525));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net525 (.A(clknet_0_net525),
    .X(clknet_1_0__leaf_net525));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net525 (.A(clknet_0_net525),
    .X(clknet_1_1__leaf_net525));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net530 (.A(net530),
    .X(clknet_0_net530));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net530 (.A(clknet_0_net530),
    .X(clknet_1_0__leaf_net530));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net530 (.A(clknet_0_net530),
    .X(clknet_1_1__leaf_net530));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net527 (.A(net527),
    .X(clknet_0_net527));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net527 (.A(clknet_0_net527),
    .X(clknet_1_0__leaf_net527));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net527 (.A(clknet_0_net527),
    .X(clknet_1_1__leaf_net527));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net521 (.A(net521),
    .X(clknet_0_net521));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net521 (.A(clknet_0_net521),
    .X(clknet_1_0__leaf_net521));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net521 (.A(clknet_0_net521),
    .X(clknet_1_1__leaf_net521));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net640 (.A(net640),
    .X(clknet_0_net640));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net640 (.A(clknet_0_net640),
    .X(clknet_1_0__leaf_net640));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net640 (.A(clknet_0_net640),
    .X(clknet_1_1__leaf_net640));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net566 (.A(net566),
    .X(clknet_0_net566));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net566 (.A(clknet_0_net566),
    .X(clknet_1_0__leaf_net566));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net566 (.A(clknet_0_net566),
    .X(clknet_1_1__leaf_net566));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net524 (.A(net524),
    .X(clknet_0_net524));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net524 (.A(clknet_0_net524),
    .X(clknet_1_0__leaf_net524));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net524 (.A(clknet_0_net524),
    .X(clknet_1_1__leaf_net524));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net251 (.A(net251),
    .X(clknet_0_net251));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net251 (.A(clknet_0_net251),
    .X(clknet_1_0__leaf_net251));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net251 (.A(clknet_0_net251),
    .X(clknet_1_1__leaf_net251));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net264 (.A(net264),
    .X(clknet_0_net264));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net264 (.A(clknet_0_net264),
    .X(clknet_1_0__leaf_net264));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net264 (.A(clknet_0_net264),
    .X(clknet_1_1__leaf_net264));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net252 (.A(net252),
    .X(clknet_0_net252));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net252 (.A(clknet_0_net252),
    .X(clknet_1_0__leaf_net252));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net252 (.A(clknet_0_net252),
    .X(clknet_1_1__leaf_net252));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net761 (.A(net761),
    .X(clknet_0_net761));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net761 (.A(clknet_0_net761),
    .X(clknet_1_0__leaf_net761));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net761 (.A(clknet_0_net761),
    .X(clknet_1_1__leaf_net761));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net96 (.A(net96),
    .X(clknet_0_net96));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net96 (.A(clknet_0_net96),
    .X(clknet_1_0__leaf_net96));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net96 (.A(clknet_0_net96),
    .X(clknet_1_1__leaf_net96));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net95 (.A(net95),
    .X(clknet_0_net95));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net95 (.A(clknet_0_net95),
    .X(clknet_1_0__leaf_net95));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net95 (.A(clknet_0_net95),
    .X(clknet_1_1__leaf_net95));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net97 (.A(net97),
    .X(clknet_0_net97));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net97 (.A(clknet_0_net97),
    .X(clknet_1_0__leaf_net97));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net97 (.A(clknet_0_net97),
    .X(clknet_1_1__leaf_net97));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net724 (.A(net724),
    .X(clknet_0_net724));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net724 (.A(clknet_0_net724),
    .X(clknet_1_0__leaf_net724));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net724 (.A(clknet_0_net724),
    .X(clknet_1_1__leaf_net724));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net725 (.A(net725),
    .X(clknet_0_net725));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net725 (.A(clknet_0_net725),
    .X(clknet_1_0__leaf_net725));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net725 (.A(clknet_0_net725),
    .X(clknet_1_1__leaf_net725));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net727 (.A(net727),
    .X(clknet_0_net727));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net727 (.A(clknet_0_net727),
    .X(clknet_1_0__leaf_net727));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net727 (.A(clknet_0_net727),
    .X(clknet_1_1__leaf_net727));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net726 (.A(net726),
    .X(clknet_0_net726));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net726 (.A(clknet_0_net726),
    .X(clknet_1_0__leaf_net726));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net726 (.A(clknet_0_net726),
    .X(clknet_1_1__leaf_net726));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net709 (.A(net709),
    .X(clknet_0_net709));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net709 (.A(clknet_0_net709),
    .X(clknet_1_0__leaf_net709));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net709 (.A(clknet_0_net709),
    .X(clknet_1_1__leaf_net709));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net710 (.A(net710),
    .X(clknet_0_net710));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net710 (.A(clknet_0_net710),
    .X(clknet_1_0__leaf_net710));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net710 (.A(clknet_0_net710),
    .X(clknet_1_1__leaf_net710));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net519 (.A(net519),
    .X(clknet_0_net519));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net519 (.A(clknet_0_net519),
    .X(clknet_1_0__leaf_net519));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net519 (.A(clknet_0_net519),
    .X(clknet_1_1__leaf_net519));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net518 (.A(net518),
    .X(clknet_0_net518));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net518 (.A(clknet_0_net518),
    .X(clknet_1_0__leaf_net518));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net518 (.A(clknet_0_net518),
    .X(clknet_1_1__leaf_net518));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net308 (.A(net308),
    .X(clknet_0_net308));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net308 (.A(clknet_0_net308),
    .X(clknet_1_0__leaf_net308));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net308 (.A(clknet_0_net308),
    .X(clknet_1_1__leaf_net308));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net306 (.A(net306),
    .X(clknet_0_net306));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net306 (.A(clknet_0_net306),
    .X(clknet_1_0__leaf_net306));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net306 (.A(clknet_0_net306),
    .X(clknet_1_1__leaf_net306));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net318 (.A(net318),
    .X(clknet_0_net318));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net318 (.A(clknet_0_net318),
    .X(clknet_1_0__leaf_net318));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net318 (.A(clknet_0_net318),
    .X(clknet_1_1__leaf_net318));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net303 (.A(net303),
    .X(clknet_0_net303));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net303 (.A(clknet_0_net303),
    .X(clknet_1_0__leaf_net303));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net303 (.A(clknet_0_net303),
    .X(clknet_1_1__leaf_net303));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net190 (.A(net190),
    .X(clknet_0_net190));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net190 (.A(clknet_0_net190),
    .X(clknet_1_0__leaf_net190));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net190 (.A(clknet_0_net190),
    .X(clknet_1_1__leaf_net190));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net187 (.A(net187),
    .X(clknet_0_net187));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net187 (.A(clknet_0_net187),
    .X(clknet_1_0__leaf_net187));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net187 (.A(clknet_0_net187),
    .X(clknet_1_1__leaf_net187));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net188 (.A(net188),
    .X(clknet_0_net188));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net188 (.A(clknet_0_net188),
    .X(clknet_1_0__leaf_net188));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net188 (.A(clknet_0_net188),
    .X(clknet_1_1__leaf_net188));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net183 (.A(net183),
    .X(clknet_0_net183));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net183 (.A(clknet_0_net183),
    .X(clknet_1_0__leaf_net183));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net183 (.A(clknet_0_net183),
    .X(clknet_1_1__leaf_net183));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net191 (.A(net191),
    .X(clknet_0_net191));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net191 (.A(clknet_0_net191),
    .X(clknet_1_0__leaf_net191));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net191 (.A(clknet_0_net191),
    .X(clknet_1_1__leaf_net191));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net194 (.A(net194),
    .X(clknet_0_net194));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net194 (.A(clknet_0_net194),
    .X(clknet_1_0__leaf_net194));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net194 (.A(clknet_0_net194),
    .X(clknet_1_1__leaf_net194));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net321 (.A(net321),
    .X(clknet_0_net321));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net321 (.A(clknet_0_net321),
    .X(clknet_1_0__leaf_net321));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net321 (.A(clknet_0_net321),
    .X(clknet_1_1__leaf_net321));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net319 (.A(net319),
    .X(clknet_0_net319));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net319 (.A(clknet_0_net319),
    .X(clknet_1_0__leaf_net319));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net319 (.A(clknet_0_net319),
    .X(clknet_1_1__leaf_net319));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net186 (.A(net186),
    .X(clknet_0_net186));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net186 (.A(clknet_0_net186),
    .X(clknet_1_0__leaf_net186));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net186 (.A(clknet_0_net186),
    .X(clknet_1_1__leaf_net186));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net185 (.A(net185),
    .X(clknet_0_net185));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net185 (.A(clknet_0_net185),
    .X(clknet_1_0__leaf_net185));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net185 (.A(clknet_0_net185),
    .X(clknet_1_1__leaf_net185));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(net323),
    .X(net841));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(net582),
    .X(net842));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(net788),
    .X(net843));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(net171),
    .X(net844));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(net559),
    .X(net845));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(net89),
    .X(net846));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(net320),
    .X(net847));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(net608),
    .X(net848));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(net751),
    .X(net849));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(net487),
    .X(net850));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(net55),
    .X(net851));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(net57),
    .X(net852));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(net173),
    .X(net853));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(net59),
    .X(net854));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(net346),
    .X(net855));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(net792),
    .X(net856));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(net750),
    .X(net857));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(net224),
    .X(net858));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(net595),
    .X(net859));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(net167),
    .X(net860));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(net307),
    .X(net861));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(net125),
    .X(net862));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(net274),
    .X(net863));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(net101),
    .X(net864));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(net120),
    .X(net865));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(net777),
    .X(net866));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(net245),
    .X(net867));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(net410),
    .X(net868));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(net276),
    .X(net869));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(net203),
    .X(net870));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(net208),
    .X(net871));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(net464),
    .X(net872));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(net752),
    .X(net873));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(net275),
    .X(net874));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(net513),
    .X(net875));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(net645),
    .X(net876));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(net514),
    .X(net877));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(net199),
    .X(net878));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(net620),
    .X(net879));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(net533),
    .X(net880));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(net650),
    .X(net881));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(net529),
    .X(net882));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(net603),
    .X(net883));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(net618),
    .X(net885));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(net729),
    .X(net886));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(net164),
    .X(net887));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(net755),
    .X(net888));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(net643),
    .X(net889));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(net560),
    .X(net890));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(net446),
    .X(net891));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(net243),
    .X(net892));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(net139),
    .X(net893));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(net337),
    .X(net894));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(net685),
    .X(net895));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(net723),
    .X(net896));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(net577),
    .X(net897));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(net583),
    .X(net898));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(net407),
    .X(net899));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(net311),
    .X(net900));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(net250),
    .X(net901));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(net482),
    .X(net902));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(net125),
    .X(net903));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(net11),
    .X(net904));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(net505),
    .X(net905));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(net574),
    .X(net906));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(net431),
    .X(net907));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(net98),
    .X(net908));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(net595),
    .X(net909));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(net233),
    .X(net910));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(net622),
    .X(net911));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(net632),
    .X(net912));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(net213),
    .X(net913));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(net393),
    .X(net914));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(net642),
    .X(net915));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(net408),
    .X(net916));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(net502),
    .X(net917));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(net27),
    .X(net918));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(net35),
    .X(net919));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(net541),
    .X(net920));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(net621),
    .X(net921));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(net348),
    .X(net922));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(net288),
    .X(net923));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(net570),
    .X(net924));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(net695),
    .X(net925));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(net247),
    .X(net926));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(net169),
    .X(net927));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(net212),
    .X(net928));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(net266),
    .X(net929));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(net483),
    .X(net931));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(net244),
    .X(net932));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(net754),
    .X(net933));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(net630),
    .X(net934));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(net241),
    .X(net935));
 sky130_fd_sc_hd__dlygate4sd3_1 hold96 (.A(net397),
    .X(net936));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(net434),
    .X(net937));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(net434),
    .X(net938));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(net232),
    .X(net939));
 sky130_fd_sc_hd__dlygate4sd3_1 hold100 (.A(net335),
    .X(net940));
 sky130_fd_sc_hd__dlygate4sd3_1 hold101 (.A(net567),
    .X(net941));
 sky130_fd_sc_hd__dlygate4sd3_1 hold102 (.A(net619),
    .X(net942));
 sky130_fd_sc_hd__dlygate4sd3_1 hold103 (.A(net424),
    .X(net943));
 sky130_fd_sc_hd__dlygate4sd3_1 hold104 (.A(net599),
    .X(net944));
 sky130_fd_sc_hd__dlygate4sd3_1 hold105 (.A(net544),
    .X(net945));
 sky130_fd_sc_hd__dlygate4sd3_1 hold106 (.A(net732),
    .X(net946));
 sky130_fd_sc_hd__dlygate4sd3_1 hold107 (.A(net581),
    .X(net947));
 sky130_fd_sc_hd__dlygate4sd3_1 hold108 (.A(net376),
    .X(net948));
 sky130_fd_sc_hd__dlygate4sd3_1 hold109 (.A(net290),
    .X(net949));
 sky130_fd_sc_hd__dlygate4sd3_1 hold110 (.A(net98),
    .X(net950));
 sky130_fd_sc_hd__dlygate4sd3_1 hold111 (.A(net53),
    .X(net951));
 sky130_fd_sc_hd__dlygate4sd3_1 hold112 (.A(net12),
    .X(net952));
 sky130_fd_sc_hd__dlygate4sd3_1 hold113 (.A(net228),
    .X(net953));
 sky130_fd_sc_hd__dlygate4sd3_1 hold114 (.A(net83),
    .X(net954));
 sky130_fd_sc_hd__dlygate4sd3_1 hold115 (.A(net374),
    .X(net955));
 sky130_fd_sc_hd__dlygate4sd3_1 hold116 (.A(net364),
    .X(net956));
 sky130_fd_sc_hd__dlygate4sd3_1 hold117 (.A(net259),
    .X(net957));
 sky130_fd_sc_hd__dlygate4sd3_1 hold118 (.A(net181),
    .X(net958));
 sky130_fd_sc_hd__dlygate4sd3_1 hold119 (.A(net88),
    .X(net959));
 sky130_fd_sc_hd__dlygate4sd3_1 hold121 (.A(net672),
    .X(net961));
 sky130_fd_sc_hd__dlygate4sd3_1 hold122 (.A(net383),
    .X(net962));
 sky130_fd_sc_hd__dlygate4sd3_1 hold123 (.A(net338),
    .X(net963));
 sky130_fd_sc_hd__dlygate4sd3_1 hold124 (.A(net123),
    .X(net964));
 sky130_fd_sc_hd__dlygate4sd3_1 hold125 (.A(net238),
    .X(net965));
 sky130_fd_sc_hd__dlygate4sd3_1 hold126 (.A(net32),
    .X(net966));
 sky130_fd_sc_hd__dlygate4sd3_1 hold127 (.A(net511),
    .X(net967));
 sky130_fd_sc_hd__dlygate4sd3_1 hold128 (.A(net601),
    .X(net968));
 sky130_fd_sc_hd__dlygate4sd3_1 hold129 (.A(net353),
    .X(net969));
 sky130_fd_sc_hd__dlygate4sd3_1 hold130 (.A(net748),
    .X(net970));
 sky130_fd_sc_hd__dlygate4sd3_1 hold131 (.A(net58),
    .X(net971));
 sky130_fd_sc_hd__dlygate4sd3_1 hold132 (.A(net690),
    .X(net972));
 sky130_fd_sc_hd__dlygate4sd3_1 hold133 (.A(net299),
    .X(net973));
 sky130_fd_sc_hd__dlygate4sd3_1 hold134 (.A(net210),
    .X(net974));
 sky130_fd_sc_hd__dlygate4sd3_1 hold135 (.A(net138),
    .X(net975));
 sky130_fd_sc_hd__dlygate4sd3_1 hold136 (.A(net347),
    .X(net976));
 sky130_fd_sc_hd__dlygate4sd3_1 hold137 (.A(net375),
    .X(net977));
 sky130_fd_sc_hd__dlygate4sd3_1 hold138 (.A(net653),
    .X(net978));
 sky130_fd_sc_hd__dlygate4sd3_1 hold139 (.A(net419),
    .X(net979));
 sky130_fd_sc_hd__dlygate4sd3_1 hold140 (.A(net104),
    .X(net980));
 sky130_fd_sc_hd__dlygate4sd3_1 hold141 (.A(net789),
    .X(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_A (.DIODE(clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(in0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(in1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(in10));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(in11));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(in12));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(in13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c42_A (.DIODE(in14));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(in15));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(in16));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(in17));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(in18));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(in19));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(in2));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(in20));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(in21));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(in22));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(in23));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(in24));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(in3));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(in4));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(in5));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(in6));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_A (.DIODE(in7));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_A (.DIODE(in8));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_A (.DIODE(in9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c527_B (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_B (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_c277_D (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_c274_RESET_B (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_c273_B (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_SCD (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_C (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_A3 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_X (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_c698_A (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA_c546_A (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_SCD (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_Q (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA_c83_S0 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_c82_S0 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_c80_C (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_c76_D_N (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_c72_SCE (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_c71_B (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_c69_B (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_c68_A (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_c67_X (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_A (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_c190_B (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge751_SCD (.DIODE(net553));
 sky130_fd_sc_hd__diode_2 ANTENNA_c651_B (.DIODE(net553));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_B (.DIODE(net553));
 sky130_fd_sc_hd__diode_2 ANTENNA_c565_A (.DIODE(net553));
 sky130_fd_sc_hd__diode_2 ANTENNA_c558_S0 (.DIODE(net553));
 sky130_fd_sc_hd__diode_2 ANTENNA_c542_SCE (.DIODE(net553));
 sky130_fd_sc_hd__diode_2 ANTENNA_c541_B (.DIODE(net553));
 sky130_fd_sc_hd__diode_2 ANTENNA_c538_SCD (.DIODE(net553));
 sky130_fd_sc_hd__diode_2 ANTENNA_c537_B (.DIODE(net553));
 sky130_fd_sc_hd__diode_2 ANTENNA_c536_X (.DIODE(net553));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout45_X (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_SCE (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_SCE (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_SCE (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_SET_B (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_output26_A (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_SCE (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_S1 (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_SCE (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_SET_B (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_SET_B (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_3__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_2__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_1__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_0__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_X (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_37_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_36_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_35_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_34_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_33_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_32_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_31_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_30_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_29_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_0_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_0__f_clk_X (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_9_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_8_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_7_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_6_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_5_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_4_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_3_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_2_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_1_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_1__f_clk_X (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_28_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_27_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_26_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_25_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_24_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_23_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_22_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_21_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_20_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_2__f_clk_X (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_19_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_18_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_17_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_16_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_15_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_14_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_13_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_12_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_11_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_10_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_3__f_clk_X (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(net366));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_283 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_255 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_338 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_468 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_566 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_595 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_354 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_552 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_84 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_553 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_62 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_407 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_600 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_624 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_133 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_71 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_552 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_17 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_422 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_602 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_10 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_22 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_554 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_608 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_564 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_578 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_5 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_116 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_438 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_588 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_507 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_562 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_245 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_522 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_273 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_22 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_8 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_22 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_542 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_562 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_534 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_356 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_479 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_548 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_494 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_301 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_617 ();
endmodule
