module netlist_1 (clk,
    in0,
    in1,
    in10,
    in11,
    in12,
    in13,
    in14,
    in15,
    in16,
    in17,
    in18,
    in19,
    in2,
    in20,
    in21,
    in22,
    in23,
    in24,
    in25,
    in26,
    in27,
    in28,
    in29,
    in3,
    in30,
    in31,
    in32,
    in33,
    in34,
    in35,
    in36,
    in37,
    in38,
    in39,
    in4,
    in40,
    in41,
    in42,
    in43,
    in44,
    in45,
    in46,
    in47,
    in48,
    in49,
    in5,
    in50,
    in51,
    in52,
    in53,
    in54,
    in55,
    in56,
    in57,
    in58,
    in59,
    in6,
    in60,
    in61,
    in7,
    in8,
    in9,
    out0,
    out1,
    out10,
    out11,
    out12,
    out13,
    out14,
    out15,
    out16,
    out17,
    out18,
    out19,
    out2,
    out20,
    out21,
    out22,
    out23,
    out24,
    out25,
    out26,
    out27,
    out28,
    out29,
    out3,
    out30,
    out31,
    out32,
    out33,
    out34,
    out35,
    out36,
    out37,
    out38,
    out39,
    out4,
    out40,
    out41,
    out42,
    out43,
    out44,
    out45,
    out46,
    out47,
    out48,
    out49,
    out5,
    out50,
    out51,
    out52,
    out53,
    out54,
    out55,
    out56,
    out57,
    out58,
    out59,
    out6,
    out60,
    out61,
    out7,
    out8,
    out9,
    rst);
 input clk;
 input in0;
 input in1;
 input in10;
 input in11;
 input in12;
 input in13;
 input in14;
 input in15;
 input in16;
 input in17;
 input in18;
 input in19;
 input in2;
 input in20;
 input in21;
 input in22;
 input in23;
 input in24;
 input in25;
 input in26;
 input in27;
 input in28;
 input in29;
 input in3;
 input in30;
 input in31;
 input in32;
 input in33;
 input in34;
 input in35;
 input in36;
 input in37;
 input in38;
 input in39;
 input in4;
 input in40;
 input in41;
 input in42;
 input in43;
 input in44;
 input in45;
 input in46;
 input in47;
 input in48;
 input in49;
 input in5;
 input in50;
 input in51;
 input in52;
 input in53;
 input in54;
 input in55;
 input in56;
 input in57;
 input in58;
 input in59;
 input in6;
 input in60;
 input in61;
 input in7;
 input in8;
 input in9;
 output out0;
 output out1;
 output out10;
 output out11;
 output out12;
 output out13;
 output out14;
 output out15;
 output out16;
 output out17;
 output out18;
 output out19;
 output out2;
 output out20;
 output out21;
 output out22;
 output out23;
 output out24;
 output out25;
 output out26;
 output out27;
 output out28;
 output out29;
 output out3;
 output out30;
 output out31;
 output out32;
 output out33;
 output out34;
 output out35;
 output out36;
 output out37;
 output out38;
 output out39;
 output out4;
 output out40;
 output out41;
 output out42;
 output out43;
 output out44;
 output out45;
 output out46;
 output out47;
 output out48;
 output out49;
 output out5;
 output out50;
 output out51;
 output out52;
 output out53;
 output out54;
 output out55;
 output out56;
 output out57;
 output out58;
 output out59;
 output out6;
 output out60;
 output out61;
 output out7;
 output out8;
 output out9;
 input rst;

 wire net0;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net63;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net64;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net65;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net66;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net67;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net617;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_0_net664;
 wire clknet_1_0__leaf_net664;
 wire clknet_1_1__leaf_net664;
 wire clknet_0_net663;
 wire clknet_1_0__leaf_net663;
 wire clknet_1_1__leaf_net663;
 wire clknet_0_net764;
 wire clknet_1_0__leaf_net764;
 wire clknet_1_1__leaf_net764;
 wire clknet_0_net750;
 wire clknet_1_0__leaf_net750;
 wire clknet_1_1__leaf_net750;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;

 sky130_fd_sc_hd__xnor2_4 c100 (.A(net31),
    .B(net35),
    .Y(net37));
 sky130_fd_sc_hd__xnor2_4 c101 (.A(net728),
    .B(net905),
    .Y(net789));
 sky130_fd_sc_hd__a21bo_1 c102 (.A1(net27),
    .A2(net31),
    .B1_N(net25),
    .X(net38));
 sky130_fd_sc_hd__xnor2_2 c103 (.A(net38),
    .B(net789),
    .Y(net39));
 sky130_fd_sc_hd__xnor2_2 c104 (.A(net36),
    .B(net30),
    .Y(net40));
 sky130_fd_sc_hd__a21bo_1 c105 (.A1(net34),
    .A2(net35),
    .B1_N(net39),
    .X(net41));
 sky130_fd_sc_hd__xnor2_4 c106 (.A(net30),
    .B(net34),
    .Y(net42));
 sky130_fd_sc_hd__xnor2_1 c107 (.A(net40),
    .B(net905),
    .Y(net43));
 sky130_fd_sc_hd__a21bo_1 c108 (.A1(net35),
    .A2(net43),
    .B1_N(net38),
    .X(net44));
 sky130_fd_sc_hd__a41o_1 c109 (.A1(net44),
    .A2(net41),
    .A3(net43),
    .A4(net2),
    .B1(net33),
    .X(net45));
 sky130_fd_sc_hd__xnor2_2 c110 (.A(net723),
    .B(net726),
    .Y(net46));
 sky130_fd_sc_hd__xnor2_1 c111 (.A(net46),
    .B(net724),
    .Y(net774));
 sky130_fd_sc_hd__xnor2_2 c112 (.A(net46),
    .B(net726),
    .Y(net47));
 sky130_fd_sc_hd__xnor2_2 c113 (.A(net721),
    .B(net32),
    .Y(net48));
 sky130_fd_sc_hd__xnor2_2 c114 (.A(net808),
    .B(net721),
    .Y(net49));
 sky130_fd_sc_hd__xnor2_1 c115 (.A(net30),
    .B(net46),
    .Y(net50));
 sky130_fd_sc_hd__xnor2_1 c116 (.A(net726),
    .B(net32),
    .Y(net51));
 sky130_fd_sc_hd__xnor2_4 c117 (.A(net49),
    .B(net5),
    .Y(net52));
 sky130_fd_sc_hd__xnor2_4 c118 (.A(net48),
    .B(net52),
    .Y(net768));
 sky130_fd_sc_hd__xnor2_1 c119 (.A(net32),
    .B(net52),
    .Y(net53));
 sky130_fd_sc_hd__xnor2_2 c120 (.A(net7),
    .B(net32),
    .Y(net54));
 sky130_fd_sc_hd__xnor2_1 c121 (.A(net51),
    .B(net54),
    .Y(net55));
 sky130_fd_sc_hd__a21bo_1 c122 (.A1(net47),
    .A2(net54),
    .B1_N(net768),
    .X(net56));
 sky130_fd_sc_hd__xnor2_1 c123 (.A(net50),
    .B(net47),
    .Y(net57));
 sky130_fd_sc_hd__xnor2_1 c124 (.A(net47),
    .B(net768),
    .Y(net751));
 sky130_fd_sc_hd__xnor2_1 c125 (.A(net55),
    .B(net724),
    .Y(net58));
 sky130_fd_sc_hd__xnor2_1 c126 (.A(net54),
    .B(net58),
    .Y(net59));
 sky130_fd_sc_hd__xnor2_1 c127 (.A(net52),
    .B(net53),
    .Y(net60));
 sky130_fd_sc_hd__xnor2_1 c128 (.A(net53),
    .B(net58),
    .Y(net61));
 sky130_fd_sc_hd__a21bo_1 c129 (.A1(net60),
    .A2(net726),
    .B1_N(net718),
    .X(net62));
 sky130_fd_sc_hd__xnor2_1 c130 (.A(net56),
    .B(net52),
    .Y(net63));
 sky130_fd_sc_hd__a21bo_1 c131 (.A1(net61),
    .A2(net60),
    .B1_N(net56),
    .X(net778));
 sky130_fd_sc_hd__xnor2_4 c132 (.A(net676),
    .B(net686),
    .Y(net64));
 sky130_fd_sc_hd__xnor2_4 c133 (.A(net680),
    .B(net675),
    .Y(net65));
 sky130_fd_sc_hd__xnor2_4 c134 (.A(net683),
    .B(net729),
    .Y(net66));
 sky130_fd_sc_hd__xnor2_4 c135 (.A(net813),
    .B(net733),
    .Y(net67));
 sky130_fd_sc_hd__xnor2_4 c136 (.A(net676),
    .B(net680),
    .Y(net68));
 sky130_fd_sc_hd__xnor2_4 c137 (.A(net66),
    .B(net678),
    .Y(net69));
 sky130_fd_sc_hd__xnor2_4 c138 (.A(net732),
    .B(net829),
    .Y(net70));
 sky130_fd_sc_hd__a21bo_4 c139 (.A1(net683),
    .A2(net617),
    .B1_N(net681),
    .X(net71));
 sky130_fd_sc_hd__xnor2_4 c140 (.A(net71),
    .B(net819),
    .Y(net72));
 sky130_fd_sc_hd__a21bo_4 c141 (.A1(net67),
    .A2(net807),
    .B1_N(net71),
    .X(net73));
 sky130_fd_sc_hd__xnor2_4 c142 (.A(net833),
    .B(net73),
    .Y(net74));
 sky130_fd_sc_hd__a21bo_4 c143 (.A1(net72),
    .A2(net70),
    .B1_N(net74),
    .X(net75));
 sky130_fd_sc_hd__xnor2_4 c144 (.A(net68),
    .B(net72),
    .Y(net76));
 sky130_fd_sc_hd__a21bo_4 c145 (.A1(net679),
    .A2(net76),
    .B1_N(net842),
    .X(net77));
 sky130_fd_sc_hd__a21bo_4 c146 (.A1(net66),
    .A2(net75),
    .B1_N(net69),
    .X(net78));
 sky130_fd_sc_hd__a21bo_4 c147 (.A1(net75),
    .A2(net687),
    .B1_N(net71),
    .X(net79));
 sky130_fd_sc_hd__a31o_4 c148 (.A1(net79),
    .A2(net684),
    .A3(net65),
    .B1(net71),
    .X(net80));
 sky130_fd_sc_hd__a21bo_4 c149 (.A1(net73),
    .A2(net78),
    .B1_N(net72),
    .X(net81));
 sky130_fd_sc_hd__xnor2_4 c150 (.A(net827),
    .B(net76),
    .Y(net82));
 sky130_fd_sc_hd__a21bo_4 c151 (.A1(net80),
    .A2(net78),
    .B1_N(net804),
    .X(net83));
 sky130_fd_sc_hd__a21bo_4 c152 (.A1(net80),
    .A2(net66),
    .B1_N(net78),
    .X(net84));
 sky130_fd_sc_hd__a41o_4 c153 (.A1(net83),
    .A2(net70),
    .A3(net82),
    .A4(net81),
    .B1(net828),
    .X(net85));
 sky130_fd_sc_hd__xnor2_4 c154 (.A(net687),
    .B(net81),
    .Y(net86));
 sky130_fd_sc_hd__xnor2_2 c155 (.A(net696),
    .B(net860),
    .Y(net87));
 sky130_fd_sc_hd__xnor2_4 c156 (.A(net698),
    .B(net801),
    .Y(net88));
 sky130_fd_sc_hd__xnor2_2 c157 (.A(net692),
    .B(net617),
    .Y(net89));
 sky130_fd_sc_hd__xnor2_1 c158 (.A(net689),
    .B(net678),
    .Y(net90));
 sky130_fd_sc_hd__xnor2_4 c159 (.A(net703),
    .B(net813),
    .Y(net91));
 sky130_fd_sc_hd__xnor2_1 c160 (.A(net709),
    .B(net68),
    .Y(net92));
 sky130_fd_sc_hd__xnor2_4 c161 (.A(net695),
    .B(net799),
    .Y(net93));
 sky130_fd_sc_hd__xnor2_4 c162 (.A(net697),
    .B(net91),
    .Y(net94));
 sky130_fd_sc_hd__xnor2_4 c163 (.A(net93),
    .B(net701),
    .Y(net95));
 sky130_fd_sc_hd__xnor2_4 c164 (.A(net682),
    .B(net94),
    .Y(net96));
 sky130_fd_sc_hd__xnor2_2 c165 (.A(net86),
    .B(net705),
    .Y(net97));
 sky130_fd_sc_hd__xnor2_4 c166 (.A(net699),
    .B(net96),
    .Y(net98));
 sky130_fd_sc_hd__xnor2_1 c167 (.A(net733),
    .B(net97),
    .Y(net99));
 sky130_fd_sc_hd__a21bo_2 c168 (.A1(net710),
    .A2(net688),
    .B1_N(net906),
    .X(net100));
 sky130_fd_sc_hd__xnor2_4 c169 (.A(net681),
    .B(net88),
    .Y(net101));
 sky130_fd_sc_hd__xnor2_4 c170 (.A(net101),
    .B(net96),
    .Y(net102));
 sky130_fd_sc_hd__xnor2_4 c171 (.A(net95),
    .B(net102),
    .Y(net770));
 sky130_fd_sc_hd__xnor2_1 c172 (.A(net99),
    .B(net100),
    .Y(net103));
 sky130_fd_sc_hd__mux4_2 c173 (.A0(net96),
    .A1(net770),
    .A2(net801),
    .A3(net102),
    .S0(net95),
    .S1(net92),
    .X(net104));
 sky130_fd_sc_hd__a21bo_2 c174 (.A1(net94),
    .A2(net685),
    .B1_N(net104),
    .X(net782));
 sky130_fd_sc_hd__xnor2_1 c175 (.A(net87),
    .B(net102),
    .Y(net105));
 sky130_fd_sc_hd__xnor2_4 c176 (.A(net3),
    .B(net721),
    .Y(net106));
 sky130_fd_sc_hd__xnor2_4 c177 (.A(net855),
    .B(net705),
    .Y(net107));
 sky130_fd_sc_hd__xnor2_1 c178 (.A(net714),
    .B(net97),
    .Y(net108));
 sky130_fd_sc_hd__xnor2_4 c179 (.A(net801),
    .B(net714),
    .Y(net109));
 sky130_fd_sc_hd__xnor2_4 c180 (.A(net727),
    .B(net839),
    .Y(net110));
 sky130_fd_sc_hd__xnor2_4 c181 (.A(net716),
    .B(net722),
    .Y(net767));
 sky130_fd_sc_hd__a21bo_2 c182 (.A1(net730),
    .A2(net110),
    .B1_N(net106),
    .X(net111));
 sky130_fd_sc_hd__xnor2_4 c183 (.A(net111),
    .B(net767),
    .Y(net112));
 sky130_fd_sc_hd__xnor2_2 c184 (.A(net112),
    .B(net3),
    .Y(net113));
 sky130_fd_sc_hd__xnor2_4 c185 (.A(net107),
    .B(net717),
    .Y(net114));
 sky130_fd_sc_hd__a21bo_2 c186 (.A1(net840),
    .A2(net106),
    .B1_N(net713),
    .X(net115));
 sky130_fd_sc_hd__xnor2_1 c187 (.A(net91),
    .B(net113),
    .Y(net116));
 sky130_fd_sc_hd__xnor2_4 c188 (.A(net711),
    .B(net110),
    .Y(net117));
 sky130_fd_sc_hd__a21bo_2 c189 (.A1(net111),
    .A2(net711),
    .B1_N(net727),
    .X(net790));
 sky130_fd_sc_hd__xnor2_1 c190 (.A(net109),
    .B(net115),
    .Y(net118));
 sky130_fd_sc_hd__xnor2_2 c191 (.A(net113),
    .B(net716),
    .Y(net119));
 sky130_fd_sc_hd__xnor2_1 c192 (.A(net118),
    .B(net767),
    .Y(net120));
 sky130_fd_sc_hd__a21bo_1 c193 (.A1(net92),
    .A2(net115),
    .B1_N(net705),
    .X(net121));
 sky130_fd_sc_hd__xnor2_4 c194 (.A(net114),
    .B(net117),
    .Y(net122));
 sky130_fd_sc_hd__a21bo_4 c195 (.A1(net108),
    .A2(net730),
    .B1_N(net118),
    .X(net123));
 sky130_fd_sc_hd__a31o_4 c196 (.A1(net116),
    .A2(net123),
    .A3(net110),
    .B1(net101),
    .X(net124));
 sky130_fd_sc_hd__a41o_4 c197 (.A1(net117),
    .A2(net120),
    .A3(net724),
    .A4(net114),
    .B1(net109),
    .X(net791));
 sky130_fd_sc_hd__xnor2_4 c198 (.A(net688),
    .B(net791),
    .Y(net125));
 sky130_fd_sc_hd__xnor2_4 c199 (.A(net903),
    .B(net107),
    .Y(net126));
 sky130_fd_sc_hd__xnor2_4 c200 (.A(net842),
    .B(net123),
    .Y(net127));
 sky130_fd_sc_hd__xnor2_4 c201 (.A(net126),
    .B(net124),
    .Y(net128));
 sky130_fd_sc_hd__xnor2_4 c202 (.A(net731),
    .B(net127),
    .Y(net129));
 sky130_fd_sc_hd__xnor2_4 c203 (.A(net129),
    .B(net909),
    .Y(net130));
 sky130_fd_sc_hd__xnor2_2 c204 (.A(net119),
    .B(net820),
    .Y(net131));
 sky130_fd_sc_hd__a31o_2 c205 (.A1(net902),
    .A2(net90),
    .A3(net131),
    .B1(net799),
    .X(net132));
 sky130_fd_sc_hd__xnor2_4 c206 (.A(net720),
    .B(net688),
    .Y(net133));
 sky130_fd_sc_hd__xnor2_4 c207 (.A(net799),
    .B(net130),
    .Y(net741));
 sky130_fd_sc_hd__xnor2_4 c208 (.A(net127),
    .B(net128),
    .Y(net763));
 sky130_fd_sc_hd__xnor2_2 c209 (.A(net132),
    .B(net802),
    .Y(net134));
 sky130_fd_sc_hd__xnor2_4 c210 (.A(net24),
    .B(net122),
    .Y(net135));
 sky130_fd_sc_hd__xnor2_2 c211 (.A(net810),
    .B(net854),
    .Y(net775));
 sky130_fd_sc_hd__xnor2_2 c212 (.A(net131),
    .B(net802),
    .Y(net136));
 sky130_fd_sc_hd__sdfbbn_1 c213 (.CLK_N(clknet_4_8_0_clk),
    .D(net133),
    .RESET_B(net132),
    .SCD(net741),
    .SCE(net129),
    .SET_B(net115),
    .Q(net138),
    .Q_N(net137));
 sky130_fd_sc_hd__xnor2_1 c214 (.A(net90),
    .B(net775),
    .Y(net139));
 sky130_fd_sc_hd__a21bo_1 c215 (.A1(net128),
    .A2(net8),
    .B1_N(net137),
    .X(net140));
 sky130_fd_sc_hd__a41o_2 c216 (.A1(net140),
    .A2(net139),
    .A3(net136),
    .A4(net138),
    .B1(net133),
    .X(net141));
 sky130_fd_sc_hd__dfbbn_1 c217 (.CLK_N(clknet_4_8_0_clk),
    .D(net705),
    .RESET_B(net139),
    .SET_B(net141),
    .Q(net143),
    .Q_N(net142));
 sky130_fd_sc_hd__a41o_1 c218 (.A1(net143),
    .A2(net133),
    .A3(net122),
    .A4(net15),
    .B1(net724),
    .X(net144));
 sky130_fd_sc_hd__a21bo_1 c219 (.A1(net144),
    .A2(net140),
    .B1_N(net142),
    .X(net769));
 sky130_fd_sc_hd__xnor2_2 c220 (.A(net134),
    .B(net22),
    .Y(net145));
 sky130_fd_sc_hd__xnor2_1 c221 (.A(net700),
    .B(net145),
    .Y(net146));
 sky130_fd_sc_hd__xnor2_1 c222 (.A(net734),
    .B(net33),
    .Y(net147));
 sky130_fd_sc_hd__clkbuf_1 c223 (.A(net622),
    .X(net148));
 sky130_fd_sc_hd__dfbbn_1 c224 (.CLK_N(clknet_4_8_0_clk),
    .D(net722),
    .RESET_B(net146),
    .SET_B(net42),
    .Q(net149));
 sky130_fd_sc_hd__xnor2_4 c225 (.A(net712),
    .B(net770),
    .Y(net150));
 sky130_fd_sc_hd__xnor2_1 c226 (.A(net145),
    .B(net790),
    .Y(net151));
 sky130_fd_sc_hd__a31o_1 c227 (.A1(net900),
    .A2(net22),
    .A3(net123),
    .B1(net125),
    .X(net152));
 sky130_fd_sc_hd__a31o_2 c228 (.A1(net40),
    .A2(net87),
    .A3(net148),
    .B1(net37),
    .X(net153));
 sky130_fd_sc_hd__a21bo_1 c229 (.A1(net147),
    .A2(net150),
    .B1_N(net39),
    .X(net154));
 sky130_fd_sc_hd__clkbuf_1 c230 (.A(net623),
    .X(net155));
 sky130_fd_sc_hd__a21bo_1 c231 (.A1(net155),
    .A2(net40),
    .B1_N(net153),
    .X(net156));
 sky130_fd_sc_hd__xnor2_4 c232 (.A(net135),
    .B(net802),
    .Y(net157));
 sky130_fd_sc_hd__a21bo_1 c233 (.A1(net22),
    .A2(net138),
    .B1_N(net157),
    .X(net785));
 sky130_fd_sc_hd__a21bo_1 c234 (.A1(net157),
    .A2(net849),
    .B1_N(net153),
    .X(net158));
 sky130_fd_sc_hd__a41o_2 c235 (.A1(net156),
    .A2(net157),
    .A3(net158),
    .A4(net134),
    .B1(net137),
    .X(net159));
 sky130_fd_sc_hd__a31o_1 c236 (.A1(net41),
    .A2(net145),
    .A3(net136),
    .B1(net157),
    .X(net160));
 sky130_fd_sc_hd__dfbbp_1 c237 (.CLK(clknet_4_10_0_clk),
    .D(net151),
    .RESET_B(net157),
    .SET_B(net160),
    .Q(net162),
    .Q_N(net161));
 sky130_fd_sc_hd__sdfxbp_1 c238 (.CLK(clknet_4_10_0_clk),
    .D(net43),
    .SCD(net886),
    .SCE(net769),
    .Q(net163));
 sky130_fd_sc_hd__sdfxbp_1 c239 (.CLK(clknet_4_10_0_clk),
    .D(net162),
    .SCD(net157),
    .SCE(net159),
    .Q(net164));
 sky130_fd_sc_hd__a21bo_1 c240 (.A1(net163),
    .A2(net162),
    .B1_N(net157),
    .X(net788));
 sky130_fd_sc_hd__a21bo_1 c241 (.A1(net887),
    .A2(net791),
    .B1_N(net790),
    .X(net165));
 sky130_fd_sc_hd__xnor2_1 c242 (.A(net63),
    .B(net36),
    .Y(net166));
 sky130_fd_sc_hd__xnor2_1 c243 (.A(net62),
    .B(net37),
    .Y(net167));
 sky130_fd_sc_hd__xnor2_1 c244 (.A(net802),
    .B(net708),
    .Y(net168));
 sky130_fd_sc_hd__xnor2_4 c245 (.A(net123),
    .B(net768),
    .Y(net169));
 sky130_fd_sc_hd__xnor2_4 c246 (.A(net35),
    .B(net169),
    .Y(net777));
 sky130_fd_sc_hd__xnor2_2 c247 (.A(net152),
    .B(net158),
    .Y(net754));
 sky130_fd_sc_hd__xnor2_1 c248 (.A(net37),
    .B(net777),
    .Y(net170));
 sky130_fd_sc_hd__xnor2_1 c249 (.A(net59),
    .B(net36),
    .Y(net773));
 sky130_fd_sc_hd__clkbuf_1 c250 (.A(net627),
    .X(net762));
 sky130_fd_sc_hd__mux4_1 c251 (.A0(net158),
    .A1(net708),
    .A2(net768),
    .A3(net704),
    .S0(net724),
    .S1(net37),
    .X(net171));
 sky130_fd_sc_hd__xnor2_1 c252 (.A(net167),
    .B(net788),
    .Y(net761));
 sky130_fd_sc_hd__mux4_1 c253 (.A0(net702),
    .A1(net36),
    .A2(net777),
    .A3(net37),
    .S0(net768),
    .S1(net154),
    .X(net172));
 sky130_fd_sc_hd__clkbuf_1 c254 (.A(net627),
    .X(net173));
 sky130_fd_sc_hd__xnor2_1 c255 (.A(net138),
    .B(net777),
    .Y(net174));
 sky130_fd_sc_hd__xnor2_1 c256 (.A(net172),
    .B(net37),
    .Y(net783));
 sky130_fd_sc_hd__xnor2_2 c257 (.A(net174),
    .B(net782),
    .Y(net786));
 sky130_fd_sc_hd__xnor2_1 c258 (.A(net168),
    .B(net777),
    .Y(net175));
 sky130_fd_sc_hd__a21bo_1 c259 (.A1(net175),
    .A2(net140),
    .B1_N(net169),
    .X(net176));
 sky130_fd_sc_hd__clkbuf_2 c260 (.A(net641),
    .X(net177));
 sky130_fd_sc_hd__xnor2_1 c261 (.A(net177),
    .B(net52),
    .Y(net757));
 sky130_fd_sc_hd__sdfbbn_1 c262 (.CLK_N(clknet_4_10_0_clk),
    .D(net173),
    .RESET_B(net177),
    .SCD(net757),
    .SCE(net777),
    .SET_B(net786),
    .Q(net780),
    .Q_N(net178));
 sky130_fd_sc_hd__mux4_1 c263 (.A0(net170),
    .A1(net178),
    .A2(net169),
    .A3(net786),
    .S0(net777),
    .S1(net52),
    .X(net179));
 sky130_fd_sc_hd__xnor2_4 c264 (.A(net82),
    .B(net804),
    .Y(net180));
 sky130_fd_sc_hd__xnor2_4 c265 (.A(net84),
    .B(net65),
    .Y(net181));
 sky130_fd_sc_hd__xnor2_4 c266 (.A(net807),
    .B(net82),
    .Y(net182));
 sky130_fd_sc_hd__xnor2_4 c267 (.A(net674),
    .B(net180),
    .Y(net183));
 sky130_fd_sc_hd__xnor2_4 c268 (.A(net853),
    .B(net71),
    .Y(net184));
 sky130_fd_sc_hd__xnor2_4 c269 (.A(net182),
    .B(net184),
    .Y(net185));
 sky130_fd_sc_hd__xnor2_4 c270 (.A(net732),
    .B(net729),
    .Y(net772));
 sky130_fd_sc_hd__xnor2_4 c271 (.A(net181),
    .B(net85),
    .Y(net186));
 sky130_fd_sc_hd__xnor2_2 c272 (.A(net707),
    .B(net71),
    .Y(net187));
 sky130_fd_sc_hd__xnor2_4 c273 (.A(net707),
    .B(net71),
    .Y(net188));
 sky130_fd_sc_hd__xnor2_4 c274 (.A(net186),
    .B(net834),
    .Y(net189));
 sky130_fd_sc_hd__a21bo_4 c275 (.A1(net822),
    .A2(net843),
    .B1_N(net181),
    .X(net190));
 sky130_fd_sc_hd__xnor2_4 c276 (.A(net190),
    .B(net188),
    .Y(net191));
 sky130_fd_sc_hd__a31o_4 c277 (.A1(net188),
    .A2(net617),
    .A3(net806),
    .B1(net811),
    .X(net192));
 sky130_fd_sc_hd__a21bo_4 c278 (.A1(net191),
    .A2(net73),
    .B1_N(net811),
    .X(net193));
 sky130_fd_sc_hd__xnor2_1 c279 (.A(net71),
    .B(net183),
    .Y(net194));
 sky130_fd_sc_hd__xnor2_4 c280 (.A(net189),
    .B(net796),
    .Y(net195));
 sky130_fd_sc_hd__xnor2_2 c281 (.A(net186),
    .B(net190),
    .Y(net196));
 sky130_fd_sc_hd__xnor2_2 c282 (.A(net195),
    .B(net187),
    .Y(net197));
 sky130_fd_sc_hd__a21bo_4 c283 (.A1(net85),
    .A2(net194),
    .B1_N(net192),
    .X(net198));
 sky130_fd_sc_hd__xnor2_4 c284 (.A(net198),
    .B(net862),
    .Y(net199));
 sky130_fd_sc_hd__a31o_4 c285 (.A1(net190),
    .A2(net197),
    .A3(net822),
    .B1(net811),
    .X(net200));
 sky130_fd_sc_hd__xnor2_4 c286 (.A(net617),
    .B(net182),
    .Y(net201));
 sky130_fd_sc_hd__a21bo_1 c287 (.A1(net182),
    .A2(net96),
    .B1_N(net201),
    .X(net202));
 sky130_fd_sc_hd__xnor2_1 c288 (.A(net190),
    .B(net685),
    .Y(net203));
 sky130_fd_sc_hd__xnor2_1 c289 (.A(net68),
    .B(net702),
    .Y(net204));
 sky130_fd_sc_hd__xnor2_1 c290 (.A(net845),
    .B(net907),
    .Y(net205));
 sky130_fd_sc_hd__xnor2_4 c291 (.A(net189),
    .B(net192),
    .Y(net206));
 sky130_fd_sc_hd__a21bo_1 c292 (.A1(net202),
    .A2(net98),
    .B1_N(net205),
    .X(net207));
 sky130_fd_sc_hd__xnor2_1 c293 (.A(net690),
    .B(net199),
    .Y(net744));
 sky130_fd_sc_hd__xnor2_2 c294 (.A(net203),
    .B(net188),
    .Y(net208));
 sky130_fd_sc_hd__clkbuf_4 c295 (.A(net671),
    .X(net746));
 sky130_fd_sc_hd__a21bo_1 c296 (.A1(net199),
    .A2(net78),
    .B1_N(net192),
    .X(net209));
 sky130_fd_sc_hd__a21bo_1 c297 (.A1(net94),
    .A2(net782),
    .B1_N(net206),
    .X(net210));
 sky130_fd_sc_hd__a21bo_2 c298 (.A1(net194),
    .A2(net185),
    .B1_N(net811),
    .X(net211));
 sky130_fd_sc_hd__xnor2_1 c299 (.A(net691),
    .B(net209),
    .Y(net212));
 sky130_fd_sc_hd__xnor2_4 c300 (.A(net676),
    .B(net206),
    .Y(net213));
 sky130_fd_sc_hd__xnor2_4 c301 (.A(net86),
    .B(net816),
    .Y(net214));
 sky130_fd_sc_hd__sdfbbp_1 c302 (.CLK(clknet_4_0_0_clk),
    .D(net211),
    .RESET_B(net204),
    .SCD(net214),
    .SCE(net213),
    .SET_B(net206),
    .Q(net216),
    .Q_N(net215));
 sky130_fd_sc_hd__a21bo_1 c303 (.A1(net813),
    .A2(net216),
    .B1_N(net211),
    .X(net217));
 sky130_fd_sc_hd__clkbuf_2 c304 (.A(net671),
    .X(net218));
 sky130_fd_sc_hd__a21bo_1 c305 (.A1(net675),
    .A2(net217),
    .B1_N(net906),
    .X(net219));
 sky130_fd_sc_hd__a41o_4 c306 (.A1(net204),
    .A2(net94),
    .A3(net206),
    .A4(net219),
    .B1(net813),
    .X(net220));
 sky130_fd_sc_hd__a41o_2 c307 (.A1(net205),
    .A2(net217),
    .A3(net103),
    .A4(net215),
    .B1(net219),
    .X(net221));
 sky130_fd_sc_hd__xnor2_1 c308 (.A(net102),
    .B(net208),
    .Y(net222));
 sky130_fd_sc_hd__xnor2_1 c309 (.A(net105),
    .B(net849),
    .Y(net223));
 sky130_fd_sc_hd__xnor2_2 c310 (.A(net208),
    .B(net124),
    .Y(net224));
 sky130_fd_sc_hd__xnor2_1 c311 (.A(net188),
    .B(net2),
    .Y(net225));
 sky130_fd_sc_hd__xnor2_1 c312 (.A(net686),
    .B(net224),
    .Y(net226));
 sky130_fd_sc_hd__xnor2_4 c313 (.A(net216),
    .B(net220),
    .Y(net227));
 sky130_fd_sc_hd__a21bo_1 c314 (.A1(net685),
    .A2(net734),
    .B1_N(net746),
    .X(net228));
 sky130_fd_sc_hd__a21bo_4 c315 (.A1(net103),
    .A2(net215),
    .B1_N(net89),
    .X(net776));
 sky130_fd_sc_hd__sdfxtp_1 c316 (.CLK(clknet_4_2_0_clk),
    .D(net226),
    .SCD(net678),
    .SCE(net216),
    .Q(net229));
 sky130_fd_sc_hd__xnor2_1 c317 (.A(net228),
    .B(net227),
    .Y(net230));
 sky130_fd_sc_hd__xnor2_1 c318 (.A(net227),
    .B(net817),
    .Y(net231));
 sky130_fd_sc_hd__buf_1 c319 (.A(net613),
    .X(net232));
 sky130_fd_sc_hd__buf_1 c320 (.A(net612),
    .X(net233));
 sky130_fd_sc_hd__sdfxtp_1 c321 (.CLK(clknet_4_2_0_clk),
    .D(net228),
    .SCD(net226),
    .SCE(net223),
    .Q(net234));
 sky130_fd_sc_hd__sdfxtp_1 c322 (.CLK(clknet_4_2_0_clk),
    .D(net230),
    .SCD(net896),
    .SCE(net721),
    .Q(net235));
 sky130_fd_sc_hd__a21bo_2 c323 (.A1(net223),
    .A2(net235),
    .B1_N(net232),
    .X(net236));
 sky130_fd_sc_hd__dfbbn_1 c324 (.CLK_N(clknet_4_2_0_clk),
    .D(net225),
    .RESET_B(net235),
    .SET_B(net231),
    .Q(net238),
    .Q_N(net237));
 sky130_fd_sc_hd__a41o_2 c325 (.A1(net233),
    .A2(net236),
    .A3(net717),
    .A4(net229),
    .B1(net776),
    .X(net239));
 sky130_fd_sc_hd__a21bo_1 c326 (.A1(net235),
    .A2(net239),
    .B1_N(net225),
    .X(net240));
 sky130_fd_sc_hd__a21bo_1 c327 (.A1(net120),
    .A2(net240),
    .B1_N(net105),
    .X(net241));
 sky130_fd_sc_hd__dfbbn_1 c328 (.CLK_N(clknet_4_8_0_clk),
    .D(net241),
    .RESET_B(net239),
    .SET_B(net233),
    .Q(net243),
    .Q_N(net242));
 sky130_fd_sc_hd__mux4_2 c329 (.A0(net232),
    .A1(net240),
    .A2(net236),
    .A3(net242),
    .S0(net241),
    .S1(net124),
    .X(net244));
 sky130_fd_sc_hd__xnor2_1 c330 (.A(net229),
    .B(net227),
    .Y(net245));
 sky130_fd_sc_hd__xnor2_1 c331 (.A(net678),
    .B(net243),
    .Y(net246));
 sky130_fd_sc_hd__a21bo_2 c332 (.A1(net246),
    .A2(net763),
    .B1_N(net115),
    .X(net743));
 sky130_fd_sc_hd__xnor2_1 c333 (.A(net864),
    .B(net240),
    .Y(net247));
 sky130_fd_sc_hd__a41o_1 c334 (.A1(net124),
    .A2(net775),
    .A3(net109),
    .A4(net133),
    .B1(net811),
    .X(net248));
 sky130_fd_sc_hd__xnor2_1 c335 (.A(net144),
    .B(net229),
    .Y(net249));
 sky130_fd_sc_hd__a21bo_1 c336 (.A1(net841),
    .A2(net106),
    .B1_N(net15),
    .X(net250));
 sky130_fd_sc_hd__a21bo_1 c337 (.A1(net249),
    .A2(net239),
    .B1_N(net248),
    .X(net735));
 sky130_fd_sc_hd__dfbbp_1 c338 (.CLK(clknet_4_8_0_clk),
    .D(net245),
    .RESET_B(net106),
    .SET_B(net246),
    .Q(net251));
 sky130_fd_sc_hd__xnor2_4 c339 (.A(net239),
    .B(net78),
    .Y(net252));
 sky130_fd_sc_hd__xnor2_2 c340 (.A(net78),
    .B(net763),
    .Y(net739));
 sky130_fd_sc_hd__buf_1 c341 (.A(net624),
    .X(net253));
 sky130_fd_sc_hd__xnor2_1 c342 (.A(net252),
    .B(net863),
    .Y(net254));
 sky130_fd_sc_hd__a21bo_1 c343 (.A1(net115),
    .A2(net725),
    .B1_N(net229),
    .X(net255));
 sky130_fd_sc_hd__xnor2_1 c344 (.A(net240),
    .B(net248),
    .Y(net256));
 sky130_fd_sc_hd__a21bo_1 c345 (.A1(net250),
    .A2(net678),
    .B1_N(net734),
    .X(net257));
 sky130_fd_sc_hd__xnor2_1 c346 (.A(net255),
    .B(net252),
    .Y(net258));
 sky130_fd_sc_hd__buf_1 c347 (.A(net624),
    .X(net259));
 sky130_fd_sc_hd__xnor2_1 c348 (.A(net257),
    .B(net645),
    .Y(net260));
 sky130_fd_sc_hd__sdfxbp_2 c349 (.CLK(clknet_4_8_0_clk),
    .D(net260),
    .SCD(net227),
    .SCE(net245),
    .Q(net262),
    .Q_N(net261));
 sky130_fd_sc_hd__mux4_1 c350 (.A0(net258),
    .A1(net130),
    .A2(net257),
    .A3(net260),
    .S0(net261),
    .S1(net246),
    .X(net263));
 sky130_fd_sc_hd__sdfxbp_1 c351 (.CLK(clknet_4_12_0_clk),
    .D(net254),
    .SCD(net247),
    .SCE(net262),
    .Q(net265),
    .Q_N(net264));
 sky130_fd_sc_hd__xnor2_4 c352 (.A(net153),
    .B(net261),
    .Y(net266));
 sky130_fd_sc_hd__xnor2_1 c353 (.A(net150),
    .B(net77),
    .Y(net267));
 sky130_fd_sc_hd__xnor2_1 c354 (.A(net851),
    .B(net259),
    .Y(net755));
 sky130_fd_sc_hd__xnor2_1 c355 (.A(net33),
    .B(net721),
    .Y(net268));
 sky130_fd_sc_hd__buf_1 c356 (.A(net629),
    .X(net269));
 sky130_fd_sc_hd__xnor2_1 c357 (.A(net136),
    .B(net849),
    .Y(net270));
 sky130_fd_sc_hd__xnor2_4 c358 (.A(net42),
    .B(net125),
    .Y(net271));
 sky130_fd_sc_hd__xnor2_1 c359 (.A(net268),
    .B(net718),
    .Y(net272));
 sky130_fd_sc_hd__xnor2_1 c360 (.A(net234),
    .B(net270),
    .Y(net273));
 sky130_fd_sc_hd__sdfrbp_1 c361 (.CLK(clknet_4_10_0_clk),
    .D(net165),
    .RESET_B(net734),
    .SCD(net271),
    .SCE(net160),
    .Q(net275),
    .Q_N(net274));
 sky130_fd_sc_hd__xnor2_1 c362 (.A(net272),
    .B(net262),
    .Y(net276));
 sky130_fd_sc_hd__a21bo_1 c363 (.A1(net130),
    .A2(net866),
    .B1_N(net271),
    .X(net765));
 sky130_fd_sc_hd__xnor2_1 c364 (.A(net273),
    .B(net812),
    .Y(net277));
 sky130_fd_sc_hd__buf_1 c365 (.A(net629),
    .X(net278));
 sky130_fd_sc_hd__clkbuf_1 c366 (.A(net641),
    .X(net279));
 sky130_fd_sc_hd__mux4_1 c367 (.A0(net106),
    .A1(net755),
    .A2(net276),
    .A3(net150),
    .S0(net271),
    .S1(net769),
    .X(net280));
 sky130_fd_sc_hd__xnor2_1 c368 (.A(net277),
    .B(net278),
    .Y(net781));
 sky130_fd_sc_hd__a21bo_1 c369 (.A1(net276),
    .A2(net850),
    .B1_N(net812),
    .X(net281));
 sky130_fd_sc_hd__dfrbp_1 c370 (.CLK(clknet_4_11_0_clk),
    .D(net281),
    .RESET_B(net765),
    .Q(net283),
    .Q_N(net282));
 sky130_fd_sc_hd__mux4_1 c371 (.A0(net852),
    .A1(net275),
    .A2(net281),
    .A3(net234),
    .S0(net271),
    .S1(net647),
    .X(net284));
 sky130_fd_sc_hd__xnor2_1 c372 (.A(net284),
    .B(net271),
    .Y(net771));
 sky130_fd_sc_hd__mux4_1 c373 (.A0(net279),
    .A1(net281),
    .A2(net743),
    .A3(net781),
    .S0(net282),
    .S1(net890),
    .X(net285));
 sky130_fd_sc_hd__mux4_1 c392 (.A0(net57),
    .A1(net177),
    .A2(net786),
    .A3(net861),
    .S0(net741),
    .S1(net761),
    .X(net286));
 sky130_fd_sc_hd__mux4_1 c393 (.A0(net154),
    .A1(net77),
    .A2(net765),
    .A3(net767),
    .S0(net177),
    .S1(clknet_1_0__leaf_net750),
    .X(net287));
 sky130_fd_sc_hd__sdfbbn_1 c394 (.CLK_N(clknet_4_10_0_clk),
    .D(net166),
    .RESET_B(net721),
    .SCD(net754),
    .SCE(clknet_1_0__leaf_net750),
    .SET_B(clknet_1_0__leaf_net764),
    .Q(net784),
    .Q_N(net288));
 sky130_fd_sc_hd__mux4_1 c395 (.A0(net267),
    .A1(net791),
    .A2(net288),
    .A3(net757),
    .S0(clknet_1_1__leaf_net750),
    .S1(clknet_1_0__leaf_net764),
    .X(net787));
 sky130_fd_sc_hd__xnor2_4 c396 (.A(net198),
    .B(net856),
    .Y(net289));
 sky130_fd_sc_hd__xnor2_4 c397 (.A(net684),
    .B(net183),
    .Y(net290));
 sky130_fd_sc_hd__xnor2_4 c398 (.A(net289),
    .B(net729),
    .Y(net291));
 sky130_fd_sc_hd__xnor2_4 c399 (.A(net289),
    .B(net70),
    .Y(net292));
 sky130_fd_sc_hd__xnor2_4 c400 (.A(net290),
    .B(net200),
    .Y(net293));
 sky130_fd_sc_hd__xnor2_4 c401 (.A(net292),
    .B(net193),
    .Y(net294));
 sky130_fd_sc_hd__xnor2_2 c402 (.A(net804),
    .B(net294),
    .Y(net295));
 sky130_fd_sc_hd__xnor2_4 c403 (.A(net291),
    .B(net859),
    .Y(net296));
 sky130_fd_sc_hd__xnor2_4 c404 (.A(net806),
    .B(net796),
    .Y(net297));
 sky130_fd_sc_hd__xnor2_4 c405 (.A(net793),
    .B(net844),
    .Y(net298));
 sky130_fd_sc_hd__clkbuf_1 c406 (.A(net611),
    .X(net299));
 sky130_fd_sc_hd__xnor2_4 c407 (.A(net296),
    .B(net298),
    .Y(net300));
 sky130_fd_sc_hd__xnor2_4 c408 (.A(net793),
    .B(net806),
    .Y(net301));
 sky130_fd_sc_hd__xnor2_4 c409 (.A(net294),
    .B(net792),
    .Y(net302));
 sky130_fd_sc_hd__xnor2_4 c410 (.A(net846),
    .B(net795),
    .Y(net303));
 sky130_fd_sc_hd__xnor2_1 c411 (.A(net301),
    .B(net303),
    .Y(net304));
 sky130_fd_sc_hd__buf_4 c412 (.A(net611),
    .X(net305));
 sky130_fd_sc_hd__clkbuf_1 c413 (.A(net639),
    .X(net306));
 sky130_fd_sc_hd__a21bo_4 c414 (.A1(net305),
    .A2(net291),
    .B1_N(net306),
    .X(net307));
 sky130_fd_sc_hd__xnor2_1 c415 (.A(net307),
    .B(net290),
    .Y(net308));
 sky130_fd_sc_hd__xnor2_1 c416 (.A(net290),
    .B(net305),
    .Y(net309));
 sky130_fd_sc_hd__a21bo_1 c417 (.A1(net308),
    .A2(net296),
    .B1_N(net305),
    .X(net310));
 sky130_fd_sc_hd__sdfrbp_1 c418 (.CLK(clknet_4_0_0_clk),
    .D(net309),
    .RESET_B(net303),
    .SCD(net310),
    .SCE(net908),
    .Q(net312),
    .Q_N(net311));
 sky130_fd_sc_hd__xnor2_4 c419 (.A(net218),
    .B(net201),
    .Y(net313));
 sky130_fd_sc_hd__a21bo_1 c420 (.A1(net312),
    .A2(net908),
    .B1_N(net301),
    .X(net314));
 sky130_fd_sc_hd__sdfxtp_1 c421 (.CLK(clknet_4_0_0_clk),
    .D(net310),
    .SCD(net857),
    .SCE(net313),
    .Q(net315));
 sky130_fd_sc_hd__xnor2_1 c422 (.A(net193),
    .B(net815),
    .Y(net316));
 sky130_fd_sc_hd__a31o_1 c423 (.A1(net210),
    .A2(net211),
    .A3(net70),
    .B1(net313),
    .X(net317));
 sky130_fd_sc_hd__a21bo_1 c424 (.A1(net211),
    .A2(net315),
    .B1_N(net863),
    .X(net318));
 sky130_fd_sc_hd__xnor2_2 c425 (.A(net201),
    .B(net312),
    .Y(net319));
 sky130_fd_sc_hd__xnor2_2 c426 (.A(net209),
    .B(net307),
    .Y(net320));
 sky130_fd_sc_hd__xnor2_2 c427 (.A(net320),
    .B(net193),
    .Y(net321));
 sky130_fd_sc_hd__a41o_2 c428 (.A1(net219),
    .A2(net318),
    .A3(net857),
    .A4(net311),
    .B1(net211),
    .X(net322));
 sky130_fd_sc_hd__sdfrtn_1 c429 (.CLK_N(clknet_4_0_0_clk),
    .D(net70),
    .RESET_B(net193),
    .SCD(net310),
    .SCE(net220),
    .Q(net323));
 sky130_fd_sc_hd__a21bo_1 c430 (.A1(net306),
    .A2(net313),
    .B1_N(net210),
    .X(net324));
 sky130_fd_sc_hd__xnor2_1 c431 (.A(net299),
    .B(net324),
    .Y(net325));
 sky130_fd_sc_hd__mux4_1 c432 (.A0(net314),
    .A1(net303),
    .A2(net320),
    .A3(net325),
    .S0(net321),
    .S1(net211),
    .X(net326));
 sky130_fd_sc_hd__xnor2_2 c433 (.A(net104),
    .B(net201),
    .Y(net327));
 sky130_fd_sc_hd__sdfrtp_1 c434 (.CLK(clknet_4_0_0_clk),
    .D(net317),
    .RESET_B(net323),
    .SCD(net302),
    .SCE(net794),
    .Q(net328));
 sky130_fd_sc_hd__buf_1 c435 (.A(net619),
    .X(net329));
 sky130_fd_sc_hd__mux4_1 c436 (.A0(net316),
    .A1(net313),
    .A2(net322),
    .A3(net325),
    .S0(net329),
    .S1(net811),
    .X(net330));
 sky130_fd_sc_hd__clkbuf_1 c437 (.A(net619),
    .X(net331));
 sky130_fd_sc_hd__a21bo_1 c438 (.A1(net331),
    .A2(net313),
    .B1_N(net794),
    .X(net332));
 sky130_fd_sc_hd__mux4_2 c439 (.A0(net323),
    .A1(net794),
    .A2(net332),
    .A3(net313),
    .S0(net811),
    .S1(net649),
    .X(net758));
 sky130_fd_sc_hd__xnor2_1 c440 (.A(net318),
    .B(net224),
    .Y(net333));
 sky130_fd_sc_hd__xnor2_1 c441 (.A(net313),
    .B(net717),
    .Y(net334));
 sky130_fd_sc_hd__a41o_1 c442 (.A1(net674),
    .A2(net322),
    .A3(net222),
    .A4(net725),
    .B1(net794),
    .X(net335));
 sky130_fd_sc_hd__buf_1 c443 (.A(net642),
    .X(net336));
 sky130_fd_sc_hd__xnor2_2 c444 (.A(net329),
    .B(net220),
    .Y(net337));
 sky130_fd_sc_hd__sdfxtp_1 c445 (.CLK(clknet_4_3_0_clk),
    .D(net336),
    .SCD(net236),
    .SCE(net221),
    .Q(net338));
 sky130_fd_sc_hd__clkbuf_1 c446 (.A(net618),
    .X(net339));
 sky130_fd_sc_hd__a21bo_2 c447 (.A1(net110),
    .A2(net236),
    .B1_N(net725),
    .X(net340));
 sky130_fd_sc_hd__a21bo_1 c448 (.A1(net337),
    .A2(net336),
    .B1_N(net798),
    .X(net341));
 sky130_fd_sc_hd__sdfxtp_1 c449 (.CLK(clknet_4_3_0_clk),
    .D(net335),
    .SCD(net212),
    .SCE(net715),
    .Q(net342));
 sky130_fd_sc_hd__a21bo_1 c450 (.A1(net339),
    .A2(net336),
    .B1_N(net222),
    .X(net343));
 sky130_fd_sc_hd__clkbuf_1 c451 (.A(net618),
    .X(net344));
 sky130_fd_sc_hd__xnor2_4 c452 (.A(net815),
    .B(net342),
    .Y(net345));
 sky130_fd_sc_hd__a21bo_4 c453 (.A1(net342),
    .A2(net337),
    .B1_N(net303),
    .X(net346));
 sky130_fd_sc_hd__dfbbn_1 c454 (.CLK_N(clknet_4_9_0_clk),
    .D(net875),
    .RESET_B(net322),
    .SET_B(net345),
    .Q(net348),
    .Q_N(net347));
 sky130_fd_sc_hd__sdfbbn_1 c455 (.CLK_N(clknet_4_12_0_clk),
    .D(net341),
    .RESET_B(net872),
    .SCD(net346),
    .SCE(net776),
    .SET_B(net335),
    .Q(net350),
    .Q_N(net349));
 sky130_fd_sc_hd__buf_1 c456 (.A(net640),
    .X(net351));
 sky130_fd_sc_hd__dfbbn_1 c457 (.CLK_N(clknet_4_3_0_clk),
    .D(net212),
    .RESET_B(net798),
    .SET_B(net346),
    .Q(net353),
    .Q_N(net352));
 sky130_fd_sc_hd__a21bo_1 c458 (.A1(net222),
    .A2(net352),
    .B1_N(net347),
    .X(net354));
 sky130_fd_sc_hd__mux4_1 c459 (.A0(net303),
    .A1(net353),
    .A2(net339),
    .A3(net708),
    .S0(net333),
    .S1(net242),
    .X(net355));
 sky130_fd_sc_hd__mux4_1 c460 (.A0(net89),
    .A1(net353),
    .A2(net345),
    .A3(net236),
    .S0(net350),
    .S1(net650),
    .X(net356));
 sky130_fd_sc_hd__mux4_1 c461 (.A0(net340),
    .A1(net725),
    .A2(net341),
    .A3(net345),
    .S0(net651),
    .S1(net653),
    .X(net357));
 sky130_fd_sc_hd__dlymetal6s2s_1 c462 (.A(net621),
    .X(net358));
 sky130_fd_sc_hd__xnor2_4 c463 (.A(net798),
    .B(net358),
    .Y(net359));
 sky130_fd_sc_hd__dfbbp_1 c464 (.CLK(clknet_4_9_0_clk),
    .D(net826),
    .RESET_B(net9),
    .SET_B(net865),
    .Q(net360));
 sky130_fd_sc_hd__xnor2_1 c465 (.A(net253),
    .B(net351),
    .Y(net361));
 sky130_fd_sc_hd__xnor2_4 c466 (.A(net8),
    .B(net262),
    .Y(net362));
 sky130_fd_sc_hd__a21bo_1 c467 (.A1(net892),
    .A2(net704),
    .B1_N(net674),
    .X(net363));
 sky130_fd_sc_hd__xnor2_4 c468 (.A(net360),
    .B(net133),
    .Y(net364));
 sky130_fd_sc_hd__xnor2_1 c469 (.A(net364),
    .B(net746),
    .Y(net365));
 sky130_fd_sc_hd__a21bo_1 c470 (.A1(net248),
    .A2(net359),
    .B1_N(net708),
    .X(net366));
 sky130_fd_sc_hd__a31o_2 c471 (.A1(net359),
    .A2(net798),
    .A3(net910),
    .B1(net252),
    .X(net748));
 sky130_fd_sc_hd__xnor2_2 c472 (.A(net363),
    .B(net364),
    .Y(net760));
 sky130_fd_sc_hd__xnor2_4 c473 (.A(net23),
    .B(net359),
    .Y(net756));
 sky130_fd_sc_hd__a21bo_1 c474 (.A1(net139),
    .A2(net790),
    .B1_N(net2),
    .X(net367));
 sky130_fd_sc_hd__sdfrtp_1 c475 (.CLK(clknet_4_9_0_clk),
    .D(net367),
    .RESET_B(net760),
    .SCD(net364),
    .SCE(net748),
    .Q(net368));
 sky130_fd_sc_hd__sdfrtp_1 c476 (.CLK(clknet_4_9_0_clk),
    .D(net873),
    .RESET_B(net878),
    .SCD(net756),
    .SCE(net825),
    .Q(net369));
 sky130_fd_sc_hd__a31o_1 c477 (.A1(net369),
    .A2(net344),
    .A3(net756),
    .B1(net109),
    .X(net370));
 sky130_fd_sc_hd__dlymetal6s2s_1 c478 (.A(net894),
    .X(net371));
 sky130_fd_sc_hd__mux4_1 c479 (.A0(net344),
    .A1(net2),
    .A2(net243),
    .A3(net366),
    .S0(net8),
    .S1(net300),
    .X(net372));
 sky130_fd_sc_hd__a31o_1 c480 (.A1(net364),
    .A2(net359),
    .A3(net264),
    .B1(net655),
    .X(net373));
 sky130_fd_sc_hd__sdfxbp_1 c481 (.CLK(clknet_4_9_0_clk),
    .D(net365),
    .SCD(net366),
    .SCE(net791),
    .Q(net375),
    .Q_N(net374));
 sky130_fd_sc_hd__sdfsbp_1 c482 (.CLK(clknet_4_12_0_clk),
    .D(net373),
    .SCD(net361),
    .SCE(net359),
    .SET_B(net256),
    .Q(net376));
 sky130_fd_sc_hd__mux4_1 c483 (.A0(net376),
    .A1(net756),
    .A2(net364),
    .A3(net302),
    .S0(net362),
    .S1(net655),
    .X(net377));
 sky130_fd_sc_hd__buf_2 c484 (.A(net615),
    .X(net378));
 sky130_fd_sc_hd__a21bo_1 c485 (.A1(net375),
    .A2(net266),
    .B1_N(net378),
    .X(net379));
 sky130_fd_sc_hd__clkbuf_1 c486 (.A(net614),
    .X(net752));
 sky130_fd_sc_hd__a21bo_1 c487 (.A1(net897),
    .A2(net300),
    .B1_N(net266),
    .X(net380));
 sky130_fd_sc_hd__sdfxbp_1 c488 (.CLK(clknet_4_9_0_clk),
    .D(net366),
    .SCD(net302),
    .SCE(net269),
    .Q(net382),
    .Q_N(net381));
 sky130_fd_sc_hd__sdfbbp_1 c489 (.CLK(clknet_4_12_0_clk),
    .D(net879),
    .RESET_B(net379),
    .SCD(net340),
    .SCE(net346),
    .SET_B(net371),
    .Q(net384),
    .Q_N(net383));
 sky130_fd_sc_hd__a21bo_1 c490 (.A1(net278),
    .A2(net381),
    .B1_N(net708),
    .X(net385));
 sky130_fd_sc_hd__xnor2_1 c491 (.A(net385),
    .B(net266),
    .Y(net386));
 sky130_fd_sc_hd__sdfxtp_1 c492 (.CLK(clknet_4_11_0_clk),
    .D(net259),
    .SCD(net221),
    .SCE(net2),
    .Q(net766));
 sky130_fd_sc_hd__sdfxtp_1 c493 (.CLK(clknet_4_11_0_clk),
    .D(net39),
    .SCD(net380),
    .SCE(net385),
    .Q(net387));
 sky130_fd_sc_hd__sdfxtp_1 c494 (.CLK(clknet_4_11_0_clk),
    .D(net262),
    .SCD(net748),
    .SCE(net760),
    .Q(net388));
 sky130_fd_sc_hd__a21bo_1 c495 (.A1(net388),
    .A2(net379),
    .B1_N(net745),
    .X(net389));
 sky130_fd_sc_hd__a21bo_1 c496 (.A1(net389),
    .A2(net278),
    .B1_N(net388),
    .X(net753));
 sky130_fd_sc_hd__a21bo_1 c497 (.A1(net9),
    .A2(net262),
    .B1_N(net378),
    .X(net390));
 sky130_fd_sc_hd__a41o_1 c498 (.A1(net270),
    .A2(net388),
    .A3(net269),
    .A4(net385),
    .B1(net812),
    .X(net391));
 sky130_fd_sc_hd__a21bo_1 c499 (.A1(net863),
    .A2(net382),
    .B1_N(net390),
    .X(net392));
 sky130_fd_sc_hd__mux4_1 c500 (.A0(net125),
    .A1(net159),
    .A2(net390),
    .A3(net378),
    .S0(net753),
    .S1(net758),
    .X(net393));
 sky130_fd_sc_hd__a21bo_1 c501 (.A1(net391),
    .A2(net379),
    .B1_N(net383),
    .X(net394));
 sky130_fd_sc_hd__a21bo_1 c502 (.A1(net394),
    .A2(net392),
    .B1_N(net125),
    .X(net395));
 sky130_fd_sc_hd__mux4_1 c503 (.A0(net395),
    .A1(net159),
    .A2(net753),
    .A3(net776),
    .S0(net387),
    .S1(net378),
    .X(net396));
 sky130_fd_sc_hd__a21bo_1 c504 (.A1(net386),
    .A2(net378),
    .B1_N(net387),
    .X(net397));
 sky130_fd_sc_hd__a21bo_1 c505 (.A1(net397),
    .A2(net340),
    .B1_N(net657),
    .X(net398));
 sky130_fd_sc_hd__buf_1 c528 (.A(net633),
    .X(net399));
 sky130_fd_sc_hd__xnor2_2 c529 (.A(net72),
    .B(net795),
    .Y(net400));
 sky130_fd_sc_hd__xnor2_1 c530 (.A(net400),
    .B(net301),
    .Y(net401));
 sky130_fd_sc_hd__xnor2_4 c531 (.A(net297),
    .B(net718),
    .Y(net402));
 sky130_fd_sc_hd__xnor2_2 c532 (.A(net196),
    .B(net300),
    .Y(net403));
 sky130_fd_sc_hd__buf_1 c533 (.A(net869),
    .X(net404));
 sky130_fd_sc_hd__xnor2_1 c534 (.A(net847),
    .B(net404),
    .Y(net405));
 sky130_fd_sc_hd__dfbbn_1 c535 (.CLK_N(clknet_4_1_0_clk),
    .D(net405),
    .RESET_B(net403),
    .SET_B(net196),
    .Q(net406));
 sky130_fd_sc_hd__dfrbp_1 c536 (.CLK(clknet_4_4_0_clk),
    .D(net403),
    .RESET_B(net297),
    .Q(net407));
 sky130_fd_sc_hd__xnor2_1 c537 (.A(net796),
    .B(net830),
    .Y(net408));
 sky130_fd_sc_hd__dfbbn_2 c538 (.CLK_N(clknet_4_1_0_clk),
    .D(net408),
    .RESET_B(net403),
    .SET_B(net297),
    .Q(net409));
 sky130_fd_sc_hd__a21bo_2 c539 (.A1(net294),
    .A2(net399),
    .B1_N(net402),
    .X(net410));
 sky130_fd_sc_hd__dfbbp_1 c540 (.CLK(clknet_4_1_0_clk),
    .D(net406),
    .RESET_B(net304),
    .SET_B(net848),
    .Q(net742),
    .Q_N(net411));
 sky130_fd_sc_hd__sdfxbp_1 c541 (.CLK(clknet_4_4_0_clk),
    .D(net401),
    .SCD(net295),
    .SCE(net411),
    .Q(net413),
    .Q_N(net412));
 sky130_fd_sc_hd__dfrtn_1 c542 (.CLK_N(clknet_4_4_0_clk),
    .D(net407),
    .RESET_B(net403),
    .Q(net414));
 sky130_fd_sc_hd__xnor2_4 c543 (.A(net409),
    .B(net835),
    .Y(net415));
 sky130_fd_sc_hd__dfrtp_1 c544 (.CLK(clknet_4_4_0_clk),
    .D(net410),
    .RESET_B(net405),
    .Q(net416));
 sky130_fd_sc_hd__xnor2_1 c545 (.A(net404),
    .B(net72),
    .Y(net417));
 sky130_fd_sc_hd__xnor2_2 c546 (.A(net416),
    .B(net415),
    .Y(net418));
 sky130_fd_sc_hd__xnor2_2 c547 (.A(net413),
    .B(net418),
    .Y(net419));
 sky130_fd_sc_hd__a21bo_1 c548 (.A1(net412),
    .A2(net400),
    .B1_N(net418),
    .X(net420));
 sky130_fd_sc_hd__sdfxbp_1 c549 (.CLK(clknet_4_4_0_clk),
    .D(net418),
    .SCD(net410),
    .SCE(net400),
    .Q(net422),
    .Q_N(net421));
 sky130_fd_sc_hd__xnor2_1 c550 (.A(net324),
    .B(net307),
    .Y(net423));
 sky130_fd_sc_hd__clkbuf_1 c551 (.A(net637),
    .X(net424));
 sky130_fd_sc_hd__xnor2_4 c552 (.A(net213),
    .B(net307),
    .Y(net425));
 sky130_fd_sc_hd__xnor2_1 c553 (.A(net424),
    .B(net898),
    .Y(net426));
 sky130_fd_sc_hd__xnor2_1 c554 (.A(net417),
    .B(net98),
    .Y(net427));
 sky130_fd_sc_hd__clkbuf_1 c555 (.A(net636),
    .X(net428));
 sky130_fd_sc_hd__a21bo_1 c556 (.A1(net694),
    .A2(net425),
    .B1_N(net427),
    .X(net429));
 sky130_fd_sc_hd__dfrtp_1 c557 (.CLK(clknet_4_6_0_clk),
    .D(net321),
    .RESET_B(net425),
    .Q(net430));
 sky130_fd_sc_hd__xnor2_1 c558 (.A(net425),
    .B(net792),
    .Y(net431));
 sky130_fd_sc_hd__a21bo_1 c559 (.A1(net427),
    .A2(net426),
    .B1_N(net792),
    .X(net432));
 sky130_fd_sc_hd__xnor2_1 c560 (.A(net693),
    .B(net300),
    .Y(net433));
 sky130_fd_sc_hd__sdfxtp_1 c561 (.CLK(clknet_4_6_0_clk),
    .D(net432),
    .SCD(net425),
    .SCE(net794),
    .Q(net434));
 sky130_fd_sc_hd__xnor2_4 c562 (.A(net100),
    .B(net323),
    .Y(net435));
 sky130_fd_sc_hd__dfrtp_1 c563 (.CLK(clknet_4_6_0_clk),
    .D(net429),
    .RESET_B(net425),
    .Q(net436));
 sky130_fd_sc_hd__a21bo_4 c564 (.A1(net434),
    .A2(net435),
    .B1_N(net323),
    .X(net437));
 sky130_fd_sc_hd__xnor2_1 c565 (.A(net414),
    .B(net437),
    .Y(net438));
 sky130_fd_sc_hd__mux4_1 c566 (.A0(net428),
    .A1(net433),
    .A2(net694),
    .A3(net301),
    .S0(net323),
    .S1(net425),
    .X(net439));
 sky130_fd_sc_hd__xnor2_2 c567 (.A(net414),
    .B(net658),
    .Y(net440));
 sky130_fd_sc_hd__a41o_1 c568 (.A1(net426),
    .A2(net437),
    .A3(net425),
    .A4(net746),
    .B1(net322),
    .X(net441));
 sky130_fd_sc_hd__mux4_1 c569 (.A0(net438),
    .A1(net425),
    .A2(net437),
    .A3(net746),
    .S0(net441),
    .S1(net323),
    .X(net442));
 sky130_fd_sc_hd__mux4_1 c570 (.A0(net401),
    .A1(net98),
    .A2(net427),
    .A3(net307),
    .S0(net435),
    .S1(net888),
    .X(net443));
 sky130_fd_sc_hd__dfsbp_1 c571 (.CLK(clknet_4_6_0_clk),
    .D(net431),
    .SET_B(net441),
    .Q(net445),
    .Q_N(net444));
 sky130_fd_sc_hd__xnor2_2 c572 (.A(net718),
    .B(net820),
    .Y(net446));
 sky130_fd_sc_hd__xnor2_1 c573 (.A(net419),
    .B(net338),
    .Y(net447));
 sky130_fd_sc_hd__a41o_1 c574 (.A1(net192),
    .A2(net2),
    .A3(net419),
    .A4(net340),
    .B1(net800),
    .X(net736));
 sky130_fd_sc_hd__a21bo_1 c575 (.A1(net742),
    .A2(net436),
    .B1_N(net653),
    .X(net448));
 sky130_fd_sc_hd__xnor2_1 c576 (.A(net445),
    .B(net654),
    .Y(net449));
 sky130_fd_sc_hd__xnor2_1 c577 (.A(net338),
    .B(net436),
    .Y(net450));
 sky130_fd_sc_hd__xnor2_2 c578 (.A(net800),
    .B(net654),
    .Y(net451));
 sky130_fd_sc_hd__a21bo_1 c579 (.A1(net449),
    .A2(net192),
    .B1_N(net800),
    .X(net452));
 sky130_fd_sc_hd__clkbuf_1 c580 (.A(net631),
    .X(net453));
 sky130_fd_sc_hd__xnor2_1 c581 (.A(net436),
    .B(net445),
    .Y(net454));
 sky130_fd_sc_hd__xnor2_1 c582 (.A(net452),
    .B(net652),
    .Y(net455));
 sky130_fd_sc_hd__buf_1 c583 (.A(net631),
    .X(net456));
 sky130_fd_sc_hd__clkbuf_1 c584 (.A(net643),
    .X(net457));
 sky130_fd_sc_hd__mux4_1 c585 (.A0(net224),
    .A1(net448),
    .A2(net718),
    .A3(net901),
    .S0(net708),
    .S1(net345),
    .X(net458));
 sky130_fd_sc_hd__xnor2_2 c586 (.A(net450),
    .B(net448),
    .Y(net459));
 sky130_fd_sc_hd__a21bo_1 c587 (.A1(net453),
    .A2(net459),
    .B1_N(net454),
    .X(net740));
 sky130_fd_sc_hd__a21bo_1 c588 (.A1(net206),
    .A2(net451),
    .B1_N(net459),
    .X(net460));
 sky130_fd_sc_hd__a21bo_1 c589 (.A1(net220),
    .A2(net459),
    .B1_N(net451),
    .X(net461));
 sky130_fd_sc_hd__a21bo_1 c590 (.A1(net448),
    .A2(net459),
    .B1_N(net740),
    .X(net462));
 sky130_fd_sc_hd__a21bo_1 c591 (.A1(net461),
    .A2(net451),
    .B1_N(net462),
    .X(net463));
 sky130_fd_sc_hd__sdfbbn_1 c592 (.CLK_N(clknet_4_6_0_clk),
    .D(net463),
    .RESET_B(net462),
    .SCD(net800),
    .SCE(net460),
    .SET_B(net660),
    .Q(net464));
 sky130_fd_sc_hd__xnor2_1 c593 (.A(net464),
    .B(net462),
    .Y(net465));
 sky130_fd_sc_hd__clkbuf_1 c594 (.X(net466));
 sky130_fd_sc_hd__clkbuf_1 c595 (.A(net616),
    .X(net467));
 sky130_fd_sc_hd__a21bo_1 c596 (.A1(net370),
    .A2(net460),
    .B1_N(net794),
    .X(net468));
 sky130_fd_sc_hd__a21bo_2 c597 (.A1(net319),
    .A2(net351),
    .B1_N(net740),
    .X(net469));
 sky130_fd_sc_hd__a21bo_1 c598 (.A1(net910),
    .A2(net437),
    .B1_N(net800),
    .X(net470));
 sky130_fd_sc_hd__xnor2_2 c599 (.A(net332),
    .B(net776),
    .Y(net471));
 sky130_fd_sc_hd__sdfbbn_1 c600 (.CLK_N(clknet_4_12_0_clk),
    .D(net468),
    .RESET_B(net265),
    .SCD(net824),
    .SCE(net800),
    .SET_B(net794),
    .Q(net472));
 sky130_fd_sc_hd__a21bo_1 c601 (.A1(net322),
    .A2(net715),
    .B1_N(net471),
    .X(net473));
 sky130_fd_sc_hd__a21bo_1 c602 (.A1(net821),
    .A2(net471),
    .B1_N(net371),
    .X(net474));
 sky130_fd_sc_hd__a21bo_1 c603 (.A1(net351),
    .A2(net109),
    .B1_N(net469),
    .X(net475));
 sky130_fd_sc_hd__a21bo_1 c604 (.A1(net243),
    .A2(net702),
    .B1_N(net471),
    .X(net476));
 sky130_fd_sc_hd__a21bo_2 c605 (.A1(net465),
    .A2(net910),
    .B1_N(net740),
    .X(net477));
 sky130_fd_sc_hd__a21bo_1 c606 (.A1(net467),
    .A2(net471),
    .B1_N(net319),
    .X(net478));
 sky130_fd_sc_hd__xnor2_1 c607 (.A(net371),
    .B(net77),
    .Y(net479));
 sky130_fd_sc_hd__a21bo_1 c608 (.A1(net252),
    .A2(net466),
    .B1_N(net871),
    .X(net480));
 sky130_fd_sc_hd__xnor2_1 c609 (.A(net475),
    .B(net469),
    .Y(net481));
 sky130_fd_sc_hd__a21bo_1 c610 (.A1(net236),
    .A2(net471),
    .B1_N(net469),
    .X(net482));
 sky130_fd_sc_hd__a21bo_1 c611 (.A1(net715),
    .A2(net482),
    .B1_N(net435),
    .X(net483));
 sky130_fd_sc_hd__a31o_1 c612 (.A1(net265),
    .A2(net481),
    .A3(net794),
    .B1(net477),
    .X(net484));
 sky130_fd_sc_hd__a41o_1 c613 (.A1(net708),
    .A2(net482),
    .A3(net794),
    .A4(net800),
    .B1(net477),
    .X(net485));
 sky130_fd_sc_hd__sdfbbp_1 c614 (.CLK(clknet_4_3_0_clk),
    .D(net476),
    .RESET_B(net470),
    .SCD(net322),
    .SCE(net484),
    .SET_B(net302),
    .Q(net486));
 sky130_fd_sc_hd__sdfbbn_1 c615 (.CLK_N(clknet_4_13_0_clk),
    .D(net256),
    .RESET_B(net474),
    .SCD(net481),
    .SCE(net261),
    .SET_B(net362),
    .Q(net487));
 sky130_fd_sc_hd__sdfsbp_1 c616 (.CLK(clknet_4_14_0_clk),
    .D(net340),
    .SCD(net384),
    .SCE(net345),
    .SET_B(net891),
    .Q(net738),
    .Q_N(net488));
 sky130_fd_sc_hd__sdfstp_1 c617 (.CLK(clknet_4_14_0_clk),
    .D(net221),
    .SCD(net385),
    .SCE(net735),
    .SET_B(net867),
    .Q(net489));
 sky130_fd_sc_hd__clkbuf_1 c618 (.A(net672),
    .X(net490));
 sky130_fd_sc_hd__sdfstp_1 c619 (.CLK(clknet_4_11_0_clk),
    .D(net457),
    .SCD(net776),
    .SCE(net390),
    .SET_B(net743),
    .Q(net491));
 sky130_fd_sc_hd__mux4_2 c62 (.A0(net722),
    .A1(net724),
    .A2(net706),
    .A3(net731),
    .S0(net727),
    .S1(net719),
    .X(net0));
 sky130_fd_sc_hd__a21bo_1 c620 (.A1(net2),
    .A2(net45),
    .B1_N(net271),
    .X(net492));
 sky130_fd_sc_hd__clkbuf_1 c621 (.A(net672),
    .X(net493));
 sky130_fd_sc_hd__sdfxtp_1 c622 (.CLK(clknet_4_13_0_clk),
    .D(net473),
    .SCD(net346),
    .SCE(net302),
    .Q(net494));
 sky130_fd_sc_hd__a21bo_1 c623 (.A1(net384),
    .A2(net271),
    .B1_N(net702),
    .X(net495));
 sky130_fd_sc_hd__a21bo_1 c624 (.A1(net493),
    .A2(net489),
    .B1_N(net488),
    .X(net747));
 sky130_fd_sc_hd__mux4_1 c625 (.A0(net495),
    .A1(net789),
    .A2(net790),
    .A3(net791),
    .S0(net437),
    .S1(net812),
    .X(net496));
 sky130_fd_sc_hd__sdfbbn_1 c626 (.CLK_N(clknet_4_12_0_clk),
    .D(net484),
    .RESET_B(net495),
    .SCD(net741),
    .SCE(net437),
    .SET_B(net271),
    .Q(net497));
 sky130_fd_sc_hd__a41o_1 c627 (.A1(net390),
    .A2(net491),
    .A3(net45),
    .A4(net387),
    .B1(net776),
    .X(net498));
 sky130_fd_sc_hd__a31o_1 c628 (.A1(net496),
    .A2(net490),
    .A3(net362),
    .B1(net261),
    .X(net499));
 sky130_fd_sc_hd__sdfxtp_1 c629 (.CLK(clknet_4_11_0_clk),
    .D(net498),
    .SCD(net718),
    .SCE(net765),
    .Q(net737));
 sky130_fd_sc_hd__mux4_2 c63 (.A0(net712),
    .A1(net716),
    .A2(net700),
    .A3(net727),
    .S0(net0),
    .S1(net721),
    .X(net1));
 sky130_fd_sc_hd__mux4_1 c630 (.A0(net269),
    .A1(net702),
    .A2(net221),
    .A3(net485),
    .S0(net390),
    .S1(net109),
    .X(net500));
 sky130_fd_sc_hd__a21bo_1 c631 (.A1(net492),
    .A2(net744),
    .B1_N(net661),
    .X(net501));
 sky130_fd_sc_hd__dfbbn_1 c632 (.CLK_N(clknet_4_14_0_clk),
    .D(net266),
    .RESET_B(net302),
    .SET_B(net812),
    .Q(net502));
 sky130_fd_sc_hd__a21bo_1 c633 (.A1(net437),
    .A2(net398),
    .B1_N(net501),
    .X(net503));
 sky130_fd_sc_hd__dfbbn_1 c634 (.CLK_N(clknet_4_12_0_clk),
    .D(net876),
    .RESET_B(net503),
    .SET_B(net340),
    .Q(net504));
 sky130_fd_sc_hd__a41o_1 c635 (.A1(net880),
    .A2(net504),
    .A3(net378),
    .A4(net437),
    .B1(net473),
    .X(net505));
 sky130_fd_sc_hd__dfbbp_1 c636 (.CLK(clknet_4_15_0_clk),
    .D(net505),
    .RESET_B(net502),
    .SET_B(net868),
    .Q(net506));
 sky130_fd_sc_hd__sdfstp_1 c637 (.CLK(clknet_4_14_0_clk),
    .D(net499),
    .SCD(net506),
    .SCE(net501),
    .SET_B(net302),
    .Q(net507));
 sky130_fd_sc_hd__mux4_2 c64 (.A0(net730),
    .A1(net720),
    .A2(net731),
    .A3(net1),
    .S0(net724),
    .S1(net706),
    .X(net2));
 sky130_fd_sc_hd__mux4_2 c65 (.A0(net706),
    .A1(net682),
    .A2(net711),
    .A3(net679),
    .S0(net734),
    .S1(net705),
    .X(net3));
 sky130_fd_sc_hd__xnor2_2 c66 (.A(net705),
    .B(net677),
    .Y(net4));
 sky130_fd_sc_hd__buf_1 c660 (.A(net635),
    .X(net508));
 sky130_fd_sc_hd__xnor2_4 c661 (.A(net305),
    .B(net835),
    .Y(net509));
 sky130_fd_sc_hd__xnor2_1 c662 (.A(net180),
    .B(net421),
    .Y(net510));
 sky130_fd_sc_hd__clkbuf_2 c663 (.A(net635),
    .X(net511));
 sky130_fd_sc_hd__xnor2_1 c664 (.A(net832),
    .B(net814),
    .Y(net512));
 sky130_fd_sc_hd__xnor2_2 c665 (.A(net191),
    .B(net509),
    .Y(net513));
 sky130_fd_sc_hd__xnor2_4 c666 (.A(net511),
    .B(net305),
    .Y(net514));
 sky130_fd_sc_hd__xnor2_1 c667 (.A(net510),
    .B(net835),
    .Y(net515));
 sky130_fd_sc_hd__a21bo_1 c668 (.A1(net508),
    .A2(net513),
    .B1_N(net305),
    .X(net516));
 sky130_fd_sc_hd__xnor2_4 c669 (.A(net835),
    .B(net514),
    .Y(net517));
 sky130_fd_sc_hd__xnor2_4 c67 (.A(net682),
    .B(net810),
    .Y(net5));
 sky130_fd_sc_hd__dfsbp_1 c670 (.CLK(clknet_4_5_0_clk),
    .D(net295),
    .SET_B(net517),
    .Q(net519),
    .Q_N(net518));
 sky130_fd_sc_hd__dfstp_1 c671 (.CLK(clknet_4_5_0_clk),
    .D(net512),
    .SET_B(net514),
    .Q(net520));
 sky130_fd_sc_hd__dfstp_1 c672 (.CLK(clknet_4_5_0_clk),
    .D(net512),
    .SET_B(net513),
    .Q(net521));
 sky130_fd_sc_hd__xnor2_1 c673 (.A(net399),
    .B(net521),
    .Y(net522));
 sky130_fd_sc_hd__sdfxbp_1 c674 (.CLK(clknet_4_5_0_clk),
    .D(net884),
    .SCD(net410),
    .SCE(net899),
    .Q(net523));
 sky130_fd_sc_hd__sdfxbp_1 c675 (.CLK(clknet_4_5_0_clk),
    .D(net874),
    .SCD(net521),
    .SCE(net410),
    .Q(net525),
    .Q_N(net524));
 sky130_fd_sc_hd__xnor2_2 c676 (.A(net415),
    .B(net517),
    .Y(net526));
 sky130_fd_sc_hd__xnor2_1 c677 (.A(net508),
    .B(net517),
    .Y(net527));
 sky130_fd_sc_hd__a21bo_1 c678 (.A1(net513),
    .A2(net518),
    .B1_N(net509),
    .X(net528));
 sky130_fd_sc_hd__xnor2_1 c679 (.A(net528),
    .B(net524),
    .Y(net529));
 sky130_fd_sc_hd__xnor2_4 c68 (.A(net679),
    .B(net702),
    .Y(net6));
 sky130_fd_sc_hd__sdfxtp_1 c680 (.CLK(clknet_4_5_0_clk),
    .D(net527),
    .SCD(net521),
    .SCE(net529),
    .Q(net530));
 sky130_fd_sc_hd__a21bo_1 c681 (.A1(net522),
    .A2(net530),
    .B1_N(net811),
    .X(net531));
 sky130_fd_sc_hd__clkbuf_1 c682 (.A(net628),
    .X(net532));
 sky130_fd_sc_hd__xnor2_1 c683 (.A(net531),
    .B(net402),
    .Y(net533));
 sky130_fd_sc_hd__xnor2_1 c684 (.A(net523),
    .B(net402),
    .Y(net534));
 sky130_fd_sc_hd__clkbuf_1 c685 (.A(net883),
    .X(net535));
 sky130_fd_sc_hd__xnor2_2 c686 (.A(net509),
    .B(net440),
    .Y(net536));
 sky130_fd_sc_hd__a21bo_1 c687 (.A1(net315),
    .A2(net307),
    .B1_N(net402),
    .X(net537));
 sky130_fd_sc_hd__a21bo_1 c688 (.A1(net533),
    .A2(net516),
    .B1_N(net440),
    .X(net538));
 sky130_fd_sc_hd__xnor2_2 c689 (.A(net98),
    .B(net811),
    .Y(net539));
 sky130_fd_sc_hd__xnor2_4 c69 (.A(net696),
    .B(net700),
    .Y(net7));
 sky130_fd_sc_hd__sedfxbp_1 c690 (.CLK(clknet_4_7_0_clk),
    .D(net519),
    .DE(net402),
    .SCD(net538),
    .SCE(net539),
    .Q(net541),
    .Q_N(net540));
 sky130_fd_sc_hd__dfstp_1 c691 (.CLK(clknet_4_4_0_clk),
    .D(net515),
    .SET_B(net538),
    .Q(net542));
 sky130_fd_sc_hd__dlrbn_1 c692 (.D(net538),
    .GATE_N(clknet_4_7_0_clk),
    .RESET_B(net895),
    .Q(net543));
 sky130_fd_sc_hd__xnor2_1 c693 (.A(net525),
    .B(net542),
    .Y(net544));
 sky130_fd_sc_hd__dlrbn_1 c694 (.D(net543),
    .GATE_N(clknet_4_7_0_clk),
    .RESET_B(net538),
    .Q(net546),
    .Q_N(net545));
 sky130_fd_sc_hd__xnor2_1 c695 (.A(net542),
    .B(net708),
    .Y(net547));
 sky130_fd_sc_hd__xnor2_1 c696 (.A(net328),
    .B(net539),
    .Y(net548));
 sky130_fd_sc_hd__dlrbp_1 c697 (.D(net214),
    .GATE(clknet_4_5_0_clk),
    .RESET_B(net870),
    .Q(net549));
 sky130_fd_sc_hd__sdfxtp_1 c698 (.CLK(clknet_4_6_0_clk),
    .D(net443),
    .SCD(net547),
    .SCE(net542),
    .Q(net550));
 sky130_fd_sc_hd__dlrbp_1 c699 (.D(net441),
    .GATE(clknet_4_5_0_clk),
    .RESET_B(net516),
    .Q(net551));
 sky130_fd_sc_hd__xnor2_4 c70 (.A(net6),
    .B(net718),
    .Y(net8));
 sky130_fd_sc_hd__xnor2_4 c700 (.A(net549),
    .B(net536),
    .Y(net552));
 sky130_fd_sc_hd__a31o_1 c701 (.A1(net440),
    .A2(net551),
    .A3(net552),
    .B1(net77),
    .X(net553));
 sky130_fd_sc_hd__sedfxbp_1 c702 (.CLK(clknet_4_7_0_clk),
    .D(net553),
    .DE(net519),
    .SCD(net538),
    .SCE(net552),
    .Q(net555),
    .Q_N(net554));
 sky130_fd_sc_hd__a31o_2 c703 (.A1(net550),
    .A2(net532),
    .A3(net552),
    .B1(net540),
    .X(net556));
 sky130_fd_sc_hd__xnor2_1 c704 (.A(net537),
    .B(net544),
    .Y(net557));
 sky130_fd_sc_hd__a31o_1 c705 (.A1(net717),
    .A2(net121),
    .A3(net517),
    .B1(net539),
    .X(net558));
 sky130_fd_sc_hd__a21bo_1 c706 (.A1(net552),
    .A2(net800),
    .B1_N(net644),
    .X(net559));
 sky130_fd_sc_hd__clkbuf_1 c707 (.A(net626),
    .X(net560));
 sky130_fd_sc_hd__a21bo_1 c708 (.A1(net112),
    .A2(net539),
    .B1_N(net552),
    .X(net561));
 sky130_fd_sc_hd__xnor2_1 c709 (.A(net121),
    .B(net454),
    .Y(net562));
 sky130_fd_sc_hd__xnor2_4 c71 (.A(net805),
    .B(net808),
    .Y(net9));
 sky130_fd_sc_hd__xnor2_1 c710 (.A(net516),
    .B(net556),
    .Y(net563));
 sky130_fd_sc_hd__xnor2_1 c711 (.A(net561),
    .B(net800),
    .Y(net564));
 sky130_fd_sc_hd__xnor2_1 c712 (.A(net564),
    .B(net517),
    .Y(net565));
 sky130_fd_sc_hd__a31o_2 c713 (.A1(net560),
    .A2(net544),
    .A3(net556),
    .B1(net554),
    .X(net566));
 sky130_fd_sc_hd__a31o_1 c714 (.A1(net550),
    .A2(net566),
    .A3(net552),
    .B1(net645),
    .X(net567));
 sky130_fd_sc_hd__a31o_1 c715 (.A1(net454),
    .A2(net513),
    .A3(net456),
    .B1(net559),
    .X(net568));
 sky130_fd_sc_hd__xnor2_1 c716 (.A(net456),
    .B(net566),
    .Y(net569));
 sky130_fd_sc_hd__a21bo_1 c717 (.A1(net568),
    .A2(net566),
    .B1_N(net800),
    .X(net570));
 sky130_fd_sc_hd__a31o_1 c718 (.A1(net514),
    .A2(net725),
    .A3(net566),
    .B1(net435),
    .X(net571));
 sky130_fd_sc_hd__a21bo_1 c719 (.A1(net562),
    .A2(net514),
    .B1_N(net561),
    .X(net572));
 sky130_fd_sc_hd__xnor2_2 c72 (.A(net719),
    .B(net4),
    .Y(net10));
 sky130_fd_sc_hd__xnor2_1 c720 (.A(net565),
    .B(net567),
    .Y(net573));
 sky130_fd_sc_hd__buf_1 c721 (.A(net625),
    .X(net574));
 sky130_fd_sc_hd__sdfbbp_1 c722 (.CLK(clknet_4_7_0_clk),
    .D(net570),
    .RESET_B(net535),
    .SCD(net556),
    .SCE(net526),
    .SET_B(net574),
    .Q(net575));
 sky130_fd_sc_hd__a31o_1 c723 (.A1(net812),
    .A2(net301),
    .A3(net556),
    .B1(net574),
    .X(net576));
 sky130_fd_sc_hd__a21bo_1 c724 (.A1(net558),
    .A2(net575),
    .B1_N(net574),
    .X(net577));
 sky130_fd_sc_hd__a21bo_1 c725 (.A1(net569),
    .A2(net576),
    .B1_N(net574),
    .X(net578));
 sky130_fd_sc_hd__sedfxtp_1 c726 (.CLK(clknet_4_6_0_clk),
    .D(net578),
    .DE(net541),
    .SCD(net141),
    .SCE(net674),
    .Q(net579));
 sky130_fd_sc_hd__a21bo_1 c727 (.A1(net534),
    .A2(net545),
    .B1_N(net540),
    .X(net580));
 sky130_fd_sc_hd__clkbuf_1 c728 (.A(net673),
    .X(net581));
 sky130_fd_sc_hd__clkbuf_1 c729 (.A(net882),
    .X(net582));
 sky130_fd_sc_hd__xnor2_2 c73 (.A(net10),
    .B(net728),
    .Y(net11));
 sky130_fd_sc_hd__sdfbbn_1 c730 (.CLK_N(clknet_4_13_0_clk),
    .D(net141),
    .RESET_B(net446),
    .SCD(net555),
    .SCE(net435),
    .SET_B(net871),
    .Q(net584),
    .Q_N(net583));
 sky130_fd_sc_hd__sdfxtp_1 c731 (.CLK(clknet_4_7_0_clk),
    .D(net563),
    .SCD(net582),
    .SCE(net556),
    .Q(net585));
 sky130_fd_sc_hd__a21bo_1 c732 (.A1(net556),
    .A2(net585),
    .B1_N(net435),
    .X(net586));
 sky130_fd_sc_hd__a21bo_1 c733 (.A1(net725),
    .A2(net486),
    .B1_N(net517),
    .X(net587));
 sky130_fd_sc_hd__dfbbn_1 c734 (.CLK_N(clknet_4_6_0_clk),
    .D(net483),
    .RESET_B(net480),
    .SET_B(net566),
    .Q(net588));
 sky130_fd_sc_hd__a21bo_1 c735 (.A1(net517),
    .A2(net587),
    .B1_N(net581),
    .X(net589));
 sky130_fd_sc_hd__a21bo_1 c736 (.A1(net581),
    .A2(net585),
    .B1_N(net725),
    .X(net590));
 sky130_fd_sc_hd__dfbbn_1 c737 (.CLK_N(clknet_4_13_0_clk),
    .D(net361),
    .RESET_B(net566),
    .SET_B(net345),
    .Q(net591));
 sky130_fd_sc_hd__a31o_1 c738 (.A1(net579),
    .A2(net580),
    .A3(net584),
    .B1(net656),
    .X(net592));
 sky130_fd_sc_hd__a31o_1 c739 (.A1(net586),
    .A2(net435),
    .A3(net526),
    .B1(net587),
    .X(net593));
 sky130_fd_sc_hd__xnor2_4 c74 (.A(net809),
    .B(net1),
    .Y(net12));
 sky130_fd_sc_hd__a21bo_1 c740 (.A1(net588),
    .A2(net446),
    .B1_N(net541),
    .X(net594));
 sky130_fd_sc_hd__a31o_1 c741 (.A1(net559),
    .A2(net590),
    .A3(net593),
    .B1(net583),
    .X(net595));
 sky130_fd_sc_hd__dfbbp_1 c742 (.CLK(clknet_4_13_0_clk),
    .D(net594),
    .RESET_B(net591),
    .SET_B(net141),
    .Q(net596));
 sky130_fd_sc_hd__mux4_1 c743 (.A0(net574),
    .A1(net595),
    .A2(net77),
    .A3(net554),
    .S0(net702),
    .S1(net583),
    .X(net597));
 sky130_fd_sc_hd__a21bo_1 c744 (.A1(net469),
    .A2(net592),
    .B1_N(net662),
    .X(net598));
 sky130_fd_sc_hd__a41o_1 c745 (.A1(net596),
    .A2(net592),
    .A3(net556),
    .A4(net559),
    .B1(net704),
    .X(net599));
 sky130_fd_sc_hd__a21bo_1 c746 (.A1(net598),
    .A2(net548),
    .B1_N(net579),
    .X(net600));
 sky130_fd_sc_hd__sdfxbp_1 c747 (.CLK(clknet_4_13_0_clk),
    .D(net600),
    .SCD(net589),
    .SCE(net812),
    .Q(net601));
 sky130_fd_sc_hd__mux4_2 c748 (.A0(net599),
    .A1(net601),
    .A2(net362),
    .A3(net792),
    .S0(net477),
    .S1(net657),
    .X(net602));
 sky130_fd_sc_hd__mux4_1 c749 (.A0(net77),
    .A1(net477),
    .A2(net904),
    .A3(net812),
    .S0(net345),
    .S1(net657),
    .X(net603));
 sky130_fd_sc_hd__xnor2_2 c75 (.A(net11),
    .B(net809),
    .Y(net13));
 sky130_fd_sc_hd__mux4_1 c750 (.A0(net45),
    .A1(net345),
    .A2(net507),
    .A3(net387),
    .S0(net904),
    .S1(clknet_1_1__leaf_net663),
    .X(net604));
 sky130_fd_sc_hd__mux4_1 c751 (.A0(net577),
    .A1(net584),
    .A2(net387),
    .A3(net507),
    .S0(net904),
    .S1(net435),
    .X(net605));
 sky130_fd_sc_hd__mux4_1 c752 (.A0(net478),
    .A1(net362),
    .A2(net487),
    .A3(net77),
    .S0(net904),
    .S1(net584),
    .X(net606));
 sky130_fd_sc_hd__mux4_1 c753 (.A0(net378),
    .A1(net435),
    .A2(net555),
    .A3(net477),
    .S0(net602),
    .S1(clknet_1_0__leaf_net664),
    .X(net607));
 sky130_fd_sc_hd__mux4_1 c754 (.A0(net792),
    .A1(net555),
    .A2(net362),
    .A3(net602),
    .S0(clknet_1_0__leaf_net663),
    .S1(net667),
    .X(net608));
 sky130_fd_sc_hd__mux4_1 c755 (.A0(net109),
    .A1(net472),
    .A2(net904),
    .A3(net665),
    .S0(net666),
    .S1(net668),
    .X(net609));
 sky130_fd_sc_hd__mux4_1 c756 (.A0(net602),
    .A1(net477),
    .A2(net77),
    .A3(clknet_1_1__leaf_net664),
    .S0(net669),
    .S1(net670),
    .X(net610));
 sky130_fd_sc_hd__xnor2_2 c76 (.A(net13),
    .B(net700),
    .Y(net14));
 sky130_fd_sc_hd__xnor2_2 c77 (.A(net14),
    .B(net6),
    .Y(net15));
 sky130_fd_sc_hd__xnor2_2 c78 (.A(net10),
    .B(net734),
    .Y(net16));
 sky130_fd_sc_hd__xnor2_4 c79 (.A(net810),
    .B(net12),
    .Y(net17));
 sky130_fd_sc_hd__xnor2_4 c80 (.A(net17),
    .B(net16),
    .Y(net759));
 sky130_fd_sc_hd__xnor2_2 c81 (.A(net14),
    .B(net759),
    .Y(net18));
 sky130_fd_sc_hd__xnor2_1 c82 (.A(net7),
    .B(net15),
    .Y(net19));
 sky130_fd_sc_hd__a21bo_1 c83 (.A1(net19),
    .A2(net759),
    .B1_N(net18),
    .X(net20));
 sky130_fd_sc_hd__xnor2_1 c84 (.A(net18),
    .B(net7),
    .Y(net21));
 sky130_fd_sc_hd__a21bo_2 c85 (.A1(net21),
    .A2(net19),
    .B1_N(net20),
    .X(net22));
 sky130_fd_sc_hd__a21bo_4 c86 (.A1(net723),
    .A2(net22),
    .B1_N(net21),
    .X(net23));
 sky130_fd_sc_hd__a41o_4 c87 (.A1(net23),
    .A2(net723),
    .A3(net837),
    .A4(net13),
    .B1(net702),
    .X(net24));
 sky130_fd_sc_hd__xnor2_4 c88 (.A(net836),
    .B(net805),
    .Y(net25));
 sky130_fd_sc_hd__xnor2_4 c89 (.A(net803),
    .B(net808),
    .Y(net26));
 sky130_fd_sc_hd__xnor2_1 c90 (.A(net11),
    .B(net26),
    .Y(net27));
 sky130_fd_sc_hd__xnor2_4 c91 (.A(net759),
    .B(net677),
    .Y(net28));
 sky130_fd_sc_hd__xnor2_4 c92 (.A(net9),
    .B(net28),
    .Y(net29));
 sky130_fd_sc_hd__xnor2_4 c93 (.A(net26),
    .B(net803),
    .Y(net30));
 sky130_fd_sc_hd__xnor2_4 c94 (.A(net797),
    .B(net9),
    .Y(net31));
 sky130_fd_sc_hd__xnor2_4 c95 (.A(net29),
    .B(net28),
    .Y(net32));
 sky130_fd_sc_hd__a41o_1 c96 (.A1(net27),
    .A2(net30),
    .A3(net28),
    .A4(net31),
    .B1(net25),
    .X(net33));
 sky130_fd_sc_hd__a21bo_2 c97 (.A1(net20),
    .A2(net728),
    .B1_N(net702),
    .X(net34));
 sky130_fd_sc_hd__xnor2_4 c98 (.A(net25),
    .B(net704),
    .Y(net35));
 sky130_fd_sc_hd__xnor2_4 c99 (.A(net677),
    .B(net726),
    .Y(net36));
 sky130_fd_sc_hd__sedfxtp_1 merge757 (.CLK(clknet_4_1_0_clk),
    .D(net295),
    .DE(net823),
    .SCD(net302),
    .SCE(net301),
    .Q(net611));
 sky130_fd_sc_hd__sdfxbp_1 merge758 (.CLK(clknet_4_2_0_clk),
    .D(net231),
    .SCD(net112),
    .SCE(net97),
    .Q(net613),
    .Q_N(net612));
 sky130_fd_sc_hd__sdfbbn_1 merge759 (.CLK_N(clknet_4_9_0_clk),
    .D(net881),
    .RESET_B(net362),
    .SCD(net159),
    .SCE(net812),
    .SET_B(net374),
    .Q(net615),
    .Q_N(net614));
 sky130_fd_sc_hd__sdfbbp_1 merge760 (.CLK(clknet_4_6_0_clk),
    .D(net327),
    .RESET_B(net141),
    .SCE(net748),
    .SET_B(net715),
    .Q(net466),
    .Q_N(net616));
 sky130_fd_sc_hd__sedfxtp_1 merge761 (.CLK(clknet_4_2_0_clk),
    .D(net334),
    .DE(net335),
    .SCD(net333),
    .SCE(net337),
    .Q(net618));
 sky130_fd_sc_hd__sdfxtp_1 merge762 (.CLK(clknet_4_3_0_clk),
    .D(net858),
    .SCD(net325),
    .SCE(net893),
    .Q(net619));
 sky130_fd_sc_hd__sdfrbp_1 merge763 (.CLK(clknet_4_9_0_clk),
    .D(net15),
    .RESET_B(net741),
    .SCD(net824),
    .SCE(net756),
    .Q(net621),
    .Q_N(net620));
 sky130_fd_sc_hd__sdfrbp_1 merge764 (.CLK(clknet_4_8_0_clk),
    .D(net146),
    .RESET_B(net22),
    .SCD(net713),
    .SCE(net132),
    .Q(net623),
    .Q_N(net622));
 sky130_fd_sc_hd__sdfrtn_1 merge765 (.CLK_N(clknet_4_9_0_clk),
    .D(net739),
    .RESET_B(net704),
    .SCD(net247),
    .SCE(net124),
    .Q(net624));
 sky130_fd_sc_hd__sdfbbn_1 merge766 (.CLK_N(clknet_4_7_0_clk),
    .D(net346),
    .RESET_B(net571),
    .SCD(net573),
    .SCE(net566),
    .SET_B(net644),
    .Q(net626),
    .Q_N(net625));
 sky130_fd_sc_hd__sdfrtp_1 merge767 (.CLK(clknet_4_10_0_clk),
    .D(net169),
    .RESET_B(net754),
    .SCD(net171),
    .SCE(net708),
    .Q(net627));
 sky130_fd_sc_hd__sdfrtp_1 merge768 (.CLK(clknet_4_5_0_clk),
    .D(net402),
    .RESET_B(net214),
    .SCD(net521),
    .SCE(net529),
    .Q(net628));
 sky130_fd_sc_hd__sdfxtp_1 merge769 (.CLK(clknet_4_11_0_clk),
    .D(net160),
    .SCD(net743),
    .SCE(net271),
    .Q(net629));
 sky130_fd_sc_hd__mux4_1 merge770 (.A0(net207),
    .A1(net205),
    .A2(net818),
    .A3(net217),
    .S0(net214),
    .S1(net201),
    .X(net630));
 sky130_fd_sc_hd__sdfrtp_1 merge771 (.CLK(clknet_4_6_0_clk),
    .D(net877),
    .RESET_B(net345),
    .SCD(net451),
    .SCE(net354),
    .Q(net631));
 sky130_fd_sc_hd__sdfsbp_1 merge772 (.CLK(clknet_4_1_0_clk),
    .D(net304),
    .SCD(net77),
    .SCE(net838),
    .SET_B(net403),
    .Q(net633),
    .Q_N(net632));
 sky130_fd_sc_hd__mux4_1 merge773 (.A0(net447),
    .A1(net485),
    .A2(net718),
    .A3(net354),
    .S0(net479),
    .S1(net776),
    .X(net634));
 sky130_fd_sc_hd__dlrtn_1 merge774 (.D(net420),
    .GATE_N(clknet_4_4_0_clk),
    .RESET_B(net410),
    .Q(net635));
 sky130_fd_sc_hd__sdfsbp_1 merge775 (.CLK(clknet_4_1_0_clk),
    .D(net323),
    .SCD(net321),
    .SCE(net423),
    .SET_B(net794),
    .Q(net637),
    .Q_N(net636));
 sky130_fd_sc_hd__mux4_1 merge776 (.A0(net557),
    .A1(net526),
    .A2(net469),
    .A3(net572),
    .S0(net346),
    .S1(net556),
    .X(net638));
 sky130_fd_sc_hd__sdfbbn_1 merge777 (.CLK_N(clknet_4_1_0_clk),
    .D(net343),
    .RESET_B(net885),
    .SCD(net304),
    .SCE(net300),
    .SET_B(net831),
    .Q(net640),
    .Q_N(net639));
 sky130_fd_sc_hd__sdfstp_1 merge778 (.CLK(clknet_4_10_0_clk),
    .D(net889),
    .SCD(net221),
    .SCE(net176),
    .SET_B(net140),
    .Q(net641));
 sky130_fd_sc_hd__sdfbbp_1 merge779 (.CLK(clknet_4_9_0_clk),
    .D(net455),
    .RESET_B(net293),
    .SCD(net335),
    .SCE(net237),
    .SET_B(net648),
    .Q(net643),
    .Q_N(net642));
 sky130_fd_sc_hd__dfxbp_1 s780 (.CLK(clknet_4_10_0_clk),
    .D(net179),
    .Q(net779));
 sky130_fd_sc_hd__dfxbp_1 s781 (.CLK(clknet_4_6_0_clk),
    .D(net244),
    .Q(net645),
    .Q_N(net644));
 sky130_fd_sc_hd__dfxtp_1 s782 (.CLK(clknet_4_8_0_clk),
    .D(net263),
    .Q(net646));
 sky130_fd_sc_hd__dfxtp_1 s783 (.CLK(clknet_4_11_0_clk),
    .D(net280),
    .Q(net647));
 sky130_fd_sc_hd__dfxtp_1 s784 (.CLK(clknet_4_11_0_clk),
    .D(net285),
    .Q(net745));
 sky130_fd_sc_hd__dlclkp_1 s785 (.CLK(clknet_4_10_0_clk),
    .GATE(net286),
    .GCLK(net750));
 sky130_fd_sc_hd__dlclkp_2 s786 (.CLK(clknet_4_10_0_clk),
    .GATE(net287),
    .GCLK(net764));
 sky130_fd_sc_hd__dlclkp_4 s787 (.CLK(clknet_4_2_0_clk),
    .GATE(net326),
    .GCLK(net648));
 sky130_fd_sc_hd__dlxbn_1 s788 (.D(net330),
    .GATE_N(clknet_4_3_0_clk),
    .Q(net649));
 sky130_fd_sc_hd__dlxbn_1 s789 (.D(net355),
    .GATE_N(clknet_4_9_0_clk),
    .Q(net651),
    .Q_N(net650));
 sky130_fd_sc_hd__dlxbp_1 s790 (.D(net356),
    .GATE(clknet_4_12_0_clk),
    .Q(net653),
    .Q_N(net652));
 sky130_fd_sc_hd__dlxtn_1 s791 (.D(net357),
    .GATE_N(clknet_4_12_0_clk),
    .Q(net654));
 sky130_fd_sc_hd__dlxtn_1 s792 (.D(net372),
    .GATE_N(clknet_4_9_0_clk),
    .Q(net655));
 sky130_fd_sc_hd__dlxtn_1 s793 (.D(net377),
    .GATE_N(clknet_4_13_0_clk),
    .Q(net656));
 sky130_fd_sc_hd__dlxtp_1 s794 (.D(net393),
    .GATE(clknet_4_14_0_clk),
    .Q(net657));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s795 (.D(net396),
    .SLEEP_B(clknet_4_14_0_clk),
    .Q(net749));
 sky130_fd_sc_hd__dfxbp_1 s796 (.CLK(clknet_4_4_0_clk),
    .D(net439),
    .Q(net658));
 sky130_fd_sc_hd__dfxbp_1 s797 (.CLK(clknet_4_4_0_clk),
    .D(net442),
    .Q(net659));
 sky130_fd_sc_hd__dfxtp_1 s798 (.CLK(clknet_4_6_0_clk),
    .D(net458),
    .Q(net660));
 sky130_fd_sc_hd__dfxtp_1 s799 (.CLK(clknet_4_14_0_clk),
    .D(net500),
    .Q(net661));
 sky130_fd_sc_hd__dfxtp_1 s800 (.CLK(clknet_4_13_0_clk),
    .D(net597),
    .Q(net662));
 sky130_fd_sc_hd__dlclkp_1 s801 (.CLK(clknet_4_15_0_clk),
    .GATE(net603),
    .GCLK(net663));
 sky130_fd_sc_hd__dlclkp_2 s802 (.CLK(clknet_4_15_0_clk),
    .GATE(net604),
    .GCLK(net664));
 sky130_fd_sc_hd__dlclkp_4 s803 (.CLK(clknet_4_15_0_clk),
    .GATE(net605),
    .GCLK(net665));
 sky130_fd_sc_hd__dlxbn_1 s804 (.D(net606),
    .GATE_N(clknet_4_15_0_clk),
    .Q(net666));
 sky130_fd_sc_hd__dlxbn_1 s805 (.D(net607),
    .GATE_N(clknet_4_15_0_clk),
    .Q(net667));
 sky130_fd_sc_hd__dlxbp_1 s806 (.D(net608),
    .GATE(clknet_4_15_0_clk),
    .Q(net669),
    .Q_N(net668));
 sky130_fd_sc_hd__dlxtn_1 s807 (.D(net609),
    .GATE_N(clknet_4_15_0_clk),
    .Q(net670));
 sky130_fd_sc_hd__dlxtn_2 s808 (.D(net610),
    .GATE_N(clknet_4_15_0_clk));
 sky130_fd_sc_hd__dlxtn_1 s809 (.D(net630),
    .GATE_N(clknet_4_2_0_clk),
    .Q(net671));
 sky130_fd_sc_hd__dlxtp_1 s810 (.D(net634),
    .GATE(clknet_4_12_0_clk),
    .Q(net672));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s811 (.D(net638),
    .SLEEP_B(clknet_4_7_0_clk),
    .Q(net673));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Right_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Right_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Right_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Right_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Right_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Right_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Right_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Right_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Right_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Right_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Right_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Right_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Right_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Right_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Right_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Right_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Right_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Right_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Right_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Right_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Right_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_161 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_162 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_163 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_164 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_165 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_166 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_167 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_168 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_169 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_170 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_171 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_172 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_173 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_174 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_175 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_176 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_177 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_178 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_179 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_180 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_181 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_182 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Left_183 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Left_184 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Left_185 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Left_186 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Left_187 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Left_188 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Left_189 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Left_190 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Left_191 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Left_192 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Left_193 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Left_194 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Left_195 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Left_196 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Left_197 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Left_198 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Left_199 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Left_200 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Left_201 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Left_202 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Left_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1347 ();
 sky130_fd_sc_hd__clkbuf_4 input1 (.A(in0),
    .X(net617));
 sky130_fd_sc_hd__buf_4 input2 (.A(in1),
    .X(net674));
 sky130_fd_sc_hd__buf_2 input3 (.A(in10),
    .X(net675));
 sky130_fd_sc_hd__buf_4 input4 (.A(in11),
    .X(net676));
 sky130_fd_sc_hd__buf_4 input5 (.A(in12),
    .X(net677));
 sky130_fd_sc_hd__clkbuf_4 input6 (.A(in13),
    .X(net678));
 sky130_fd_sc_hd__clkbuf_4 input7 (.A(in14),
    .X(net679));
 sky130_fd_sc_hd__clkbuf_4 input8 (.A(in15),
    .X(net680));
 sky130_fd_sc_hd__buf_2 input9 (.A(in16),
    .X(net681));
 sky130_fd_sc_hd__buf_4 input10 (.A(in17),
    .X(net682));
 sky130_fd_sc_hd__buf_6 input11 (.A(in18),
    .X(net683));
 sky130_fd_sc_hd__clkbuf_2 input12 (.A(in19),
    .X(net684));
 sky130_fd_sc_hd__clkbuf_2 input13 (.A(in2),
    .X(net685));
 sky130_fd_sc_hd__buf_2 input14 (.A(in20),
    .X(net686));
 sky130_fd_sc_hd__clkbuf_2 input15 (.A(in21),
    .X(net687));
 sky130_fd_sc_hd__buf_4 input16 (.A(in22),
    .X(net688));
 sky130_fd_sc_hd__buf_1 input17 (.A(in23),
    .X(net689));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(in24),
    .X(net690));
 sky130_fd_sc_hd__buf_1 input19 (.A(in25),
    .X(net691));
 sky130_fd_sc_hd__buf_1 input20 (.A(in26),
    .X(net692));
 sky130_fd_sc_hd__buf_1 input21 (.A(in27),
    .X(net693));
 sky130_fd_sc_hd__buf_1 input22 (.A(in28),
    .X(net694));
 sky130_fd_sc_hd__clkbuf_2 input23 (.A(in29),
    .X(net695));
 sky130_fd_sc_hd__clkbuf_4 input24 (.A(in3),
    .X(net696));
 sky130_fd_sc_hd__clkbuf_2 input25 (.A(in30),
    .X(net697));
 sky130_fd_sc_hd__clkbuf_2 input26 (.A(in31),
    .X(net698));
 sky130_fd_sc_hd__clkbuf_2 input27 (.A(in32),
    .X(net699));
 sky130_fd_sc_hd__clkbuf_4 input28 (.A(in33),
    .X(net700));
 sky130_fd_sc_hd__clkbuf_2 input29 (.A(in34),
    .X(net701));
 sky130_fd_sc_hd__clkbuf_8 input30 (.A(in35),
    .X(net702));
 sky130_fd_sc_hd__clkbuf_2 input31 (.A(in36),
    .X(net703));
 sky130_fd_sc_hd__buf_4 input32 (.A(in37),
    .X(net704));
 sky130_fd_sc_hd__buf_4 input33 (.A(in38),
    .X(net705));
 sky130_fd_sc_hd__buf_1 input34 (.A(in39),
    .X(net706));
 sky130_fd_sc_hd__buf_2 input35 (.A(in4),
    .X(net707));
 sky130_fd_sc_hd__buf_4 input36 (.A(in40),
    .X(net708));
 sky130_fd_sc_hd__buf_1 input37 (.A(in41),
    .X(net709));
 sky130_fd_sc_hd__buf_1 input38 (.A(in42),
    .X(net710));
 sky130_fd_sc_hd__buf_2 input39 (.A(in43),
    .X(net711));
 sky130_fd_sc_hd__clkbuf_2 input40 (.A(in44),
    .X(net712));
 sky130_fd_sc_hd__buf_1 input41 (.A(in45),
    .X(net713));
 sky130_fd_sc_hd__clkbuf_2 input42 (.A(in46),
    .X(net714));
 sky130_fd_sc_hd__buf_2 input43 (.A(in47),
    .X(net715));
 sky130_fd_sc_hd__buf_2 input44 (.A(in48),
    .X(net716));
 sky130_fd_sc_hd__buf_4 input45 (.A(in49),
    .X(net717));
 sky130_fd_sc_hd__buf_8 input46 (.A(in5),
    .X(net718));
 sky130_fd_sc_hd__buf_1 input47 (.A(in50),
    .X(net719));
 sky130_fd_sc_hd__clkbuf_2 input48 (.A(in51),
    .X(net720));
 sky130_fd_sc_hd__clkbuf_8 input49 (.A(in52),
    .X(net721));
 sky130_fd_sc_hd__clkbuf_2 input50 (.A(in53),
    .X(net722));
 sky130_fd_sc_hd__clkbuf_2 input51 (.A(in54),
    .X(net723));
 sky130_fd_sc_hd__clkbuf_4 input52 (.A(in55),
    .X(net724));
 sky130_fd_sc_hd__clkbuf_4 input53 (.A(in56),
    .X(net725));
 sky130_fd_sc_hd__clkbuf_4 input54 (.A(in57),
    .X(net726));
 sky130_fd_sc_hd__buf_2 input55 (.A(in58),
    .X(net727));
 sky130_fd_sc_hd__buf_2 input56 (.A(in59),
    .X(net728));
 sky130_fd_sc_hd__buf_12 input57 (.A(in6),
    .X(net729));
 sky130_fd_sc_hd__dlymetal6s2s_1 input58 (.A(in60),
    .X(net730));
 sky130_fd_sc_hd__clkbuf_2 input59 (.A(in61),
    .X(net731));
 sky130_fd_sc_hd__clkbuf_4 input60 (.A(in7),
    .X(net732));
 sky130_fd_sc_hd__buf_2 input61 (.A(in8),
    .X(net733));
 sky130_fd_sc_hd__buf_4 input62 (.A(in9),
    .X(net734));
 sky130_fd_sc_hd__buf_2 output63 (.A(net735),
    .X(out0));
 sky130_fd_sc_hd__clkbuf_4 output64 (.A(net736),
    .X(out1));
 sky130_fd_sc_hd__buf_2 output65 (.A(net737),
    .X(out10));
 sky130_fd_sc_hd__buf_2 output66 (.A(net738),
    .X(out11));
 sky130_fd_sc_hd__buf_2 output67 (.A(net739),
    .X(out12));
 sky130_fd_sc_hd__clkbuf_4 output68 (.A(net740),
    .X(out13));
 sky130_fd_sc_hd__buf_2 output69 (.A(net741),
    .X(out14));
 sky130_fd_sc_hd__buf_2 output70 (.A(net742),
    .X(out15));
 sky130_fd_sc_hd__buf_2 output71 (.A(net743),
    .X(out16));
 sky130_fd_sc_hd__buf_2 output72 (.A(net744),
    .X(out17));
 sky130_fd_sc_hd__buf_2 output73 (.A(net745),
    .X(out18));
 sky130_fd_sc_hd__buf_2 output74 (.A(net746),
    .X(out19));
 sky130_fd_sc_hd__buf_2 output75 (.A(net747),
    .X(out2));
 sky130_fd_sc_hd__buf_2 output76 (.A(net748),
    .X(out20));
 sky130_fd_sc_hd__buf_2 output77 (.A(net749),
    .X(out22));
 sky130_fd_sc_hd__clkbuf_1 output78 (.A(clknet_1_1__leaf_net750),
    .X(out23));
 sky130_fd_sc_hd__buf_2 output79 (.A(net751),
    .X(out24));
 sky130_fd_sc_hd__buf_2 output80 (.A(net752),
    .X(out25));
 sky130_fd_sc_hd__buf_2 output81 (.A(net753),
    .X(out26));
 sky130_fd_sc_hd__buf_2 output82 (.A(net754),
    .X(out28));
 sky130_fd_sc_hd__buf_2 output83 (.A(net755),
    .X(out29));
 sky130_fd_sc_hd__buf_2 output84 (.A(net756),
    .X(out30));
 sky130_fd_sc_hd__buf_2 output85 (.A(net757),
    .X(out31));
 sky130_fd_sc_hd__buf_2 output86 (.A(net758),
    .X(out33));
 sky130_fd_sc_hd__buf_2 output87 (.A(net759),
    .X(out34));
 sky130_fd_sc_hd__buf_2 output88 (.A(net760),
    .X(out35));
 sky130_fd_sc_hd__buf_2 output89 (.A(net761),
    .X(out36));
 sky130_fd_sc_hd__buf_2 output90 (.A(net762),
    .X(out37));
 sky130_fd_sc_hd__buf_2 output91 (.A(net763),
    .X(out38));
 sky130_fd_sc_hd__clkbuf_1 output92 (.A(clknet_1_1__leaf_net764),
    .X(out39));
 sky130_fd_sc_hd__buf_2 output93 (.A(net765),
    .X(out4));
 sky130_fd_sc_hd__buf_2 output94 (.A(net766),
    .X(out40));
 sky130_fd_sc_hd__buf_2 output95 (.A(net767),
    .X(out41));
 sky130_fd_sc_hd__buf_2 output96 (.A(net768),
    .X(out42));
 sky130_fd_sc_hd__buf_2 output97 (.A(net769),
    .X(out43));
 sky130_fd_sc_hd__buf_2 output98 (.A(net770),
    .X(out44));
 sky130_fd_sc_hd__buf_2 output99 (.A(net771),
    .X(out45));
 sky130_fd_sc_hd__buf_2 output100 (.A(net811),
    .X(out46));
 sky130_fd_sc_hd__buf_2 output101 (.A(net773),
    .X(out47));
 sky130_fd_sc_hd__buf_2 output102 (.A(net774),
    .X(out48));
 sky130_fd_sc_hd__buf_2 output103 (.A(net775),
    .X(out49));
 sky130_fd_sc_hd__buf_2 output104 (.A(net776),
    .X(out5));
 sky130_fd_sc_hd__buf_2 output105 (.A(net777),
    .X(out50));
 sky130_fd_sc_hd__buf_2 output106 (.A(net778),
    .X(out51));
 sky130_fd_sc_hd__buf_2 output107 (.A(net779),
    .X(out52));
 sky130_fd_sc_hd__buf_2 output108 (.A(net780),
    .X(out53));
 sky130_fd_sc_hd__buf_2 output109 (.A(net781),
    .X(out54));
 sky130_fd_sc_hd__buf_2 output110 (.A(net782),
    .X(out55));
 sky130_fd_sc_hd__buf_2 output111 (.A(net783),
    .X(out56));
 sky130_fd_sc_hd__buf_2 output112 (.A(net784),
    .X(out57));
 sky130_fd_sc_hd__buf_2 output113 (.A(net785),
    .X(out59));
 sky130_fd_sc_hd__buf_2 output114 (.A(net786),
    .X(out6));
 sky130_fd_sc_hd__clkbuf_1 output115 (.A(net787),
    .X(out60));
 sky130_fd_sc_hd__buf_2 output116 (.A(net788),
    .X(out61));
 sky130_fd_sc_hd__buf_2 output117 (.A(net789),
    .X(out7));
 sky130_fd_sc_hd__buf_2 output118 (.A(net790),
    .X(out8));
 sky130_fd_sc_hd__buf_2 output119 (.A(net791),
    .X(out9));
 sky130_fd_sc_hd__buf_4 max_cap120 (.A(net300),
    .X(net792));
 sky130_fd_sc_hd__buf_4 max_cap121 (.A(net292),
    .X(net793));
 sky130_fd_sc_hd__clkbuf_4 fanout122 (.A(net327),
    .X(net794));
 sky130_fd_sc_hd__buf_4 max_cap123 (.A(net911),
    .X(net795));
 sky130_fd_sc_hd__buf_4 max_cap124 (.A(net184),
    .X(net796));
 sky130_fd_sc_hd__buf_8 max_cap125 (.A(net29),
    .X(net797));
 sky130_fd_sc_hd__buf_4 max_cap126 (.A(net93),
    .X(net798));
 sky130_fd_sc_hd__buf_4 max_cap127 (.A(net88),
    .X(net799));
 sky130_fd_sc_hd__clkbuf_4 fanout128 (.A(net446),
    .X(net800));
 sky130_fd_sc_hd__buf_4 max_cap129 (.A(net74),
    .X(net801));
 sky130_fd_sc_hd__buf_4 max_cap130 (.A(net16),
    .X(net802));
 sky130_fd_sc_hd__buf_4 max_cap131 (.A(net12),
    .X(net803));
 sky130_fd_sc_hd__buf_4 max_cap132 (.A(net76),
    .X(net804));
 sky130_fd_sc_hd__buf_4 max_cap133 (.A(net5),
    .X(net805));
 sky130_fd_sc_hd__buf_4 max_cap134 (.A(net187),
    .X(net806));
 sky130_fd_sc_hd__buf_8 max_cap135 (.A(net69),
    .X(net807));
 sky130_fd_sc_hd__buf_4 max_cap136 (.A(net809),
    .X(net808));
 sky130_fd_sc_hd__buf_4 max_cap137 (.A(net6),
    .X(net809));
 sky130_fd_sc_hd__buf_4 max_cap138 (.A(net4),
    .X(net810));
 sky130_fd_sc_hd__clkbuf_8 fanout139 (.A(net772),
    .X(net811));
 sky130_fd_sc_hd__clkbuf_4 fanout140 (.A(net772),
    .X(net812));
 sky130_fd_sc_hd__buf_8 wire141 (.A(net64),
    .X(net813));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net664 (.A(net664),
    .X(clknet_0_net664));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net664 (.A(clknet_0_net664),
    .X(clknet_1_0__leaf_net664));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net664 (.A(clknet_0_net664),
    .X(clknet_1_1__leaf_net664));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net663 (.A(net663),
    .X(clknet_0_net663));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net663 (.A(clknet_0_net663),
    .X(clknet_1_0__leaf_net663));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net663 (.A(clknet_0_net663),
    .X(clknet_1_1__leaf_net663));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net764 (.A(net764),
    .X(clknet_0_net764));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net764 (.A(clknet_0_net764),
    .X(clknet_1_0__leaf_net764));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net764 (.A(clknet_0_net764),
    .X(clknet_1_1__leaf_net764));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net750 (.A(net750),
    .X(clknet_0_net750));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net750 (.A(clknet_0_net750),
    .X(clknet_1_0__leaf_net750));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net750 (.A(clknet_0_net750),
    .X(clknet_1_1__leaf_net750));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer1 (.A(net200),
    .X(net814));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer2 (.A(net200),
    .X(net815));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer3 (.A(net200),
    .X(net816));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer4 (.A(net816),
    .X(net817));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer5 (.A(net817),
    .X(net818));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer6 (.A(net66),
    .X(net819));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer7 (.A(net73),
    .X(net820));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer8 (.A(net820),
    .X(net821));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer9 (.A(net186),
    .X(net822));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer10 (.A(net293),
    .X(net823));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer11 (.A(net293),
    .X(net824));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer12 (.A(net824),
    .X(net825));
 sky130_fd_sc_hd__buf_2 rebuffer13 (.A(net825),
    .X(net826));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer14 (.A(net74),
    .X(net827));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer15 (.A(net827),
    .X(net828));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer16 (.A(net67),
    .X(net829));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer17 (.A(net829),
    .X(net830));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer18 (.A(net830),
    .X(net831));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer19 (.A(net831),
    .X(net832));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer20 (.A(net69),
    .X(net833));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer21 (.A(net64),
    .X(net834));
 sky130_fd_sc_hd__clkbuf_8 rebuffer22 (.A(net83),
    .X(net835));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer23 (.A(net17),
    .X(net836));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer24 (.A(net836),
    .X(net837));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer25 (.A(net195),
    .X(net838));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer26 (.A(net0),
    .X(net839));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer27 (.A(net839),
    .X(net840));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer28 (.A(net181),
    .X(net841));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer29 (.A(net75),
    .X(net842));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer30 (.A(net183),
    .X(net843));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer31 (.A(net183),
    .X(net844));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer32 (.A(net197),
    .X(net845));
 sky130_fd_sc_hd__buf_2 rebuffer33 (.A(net298),
    .X(net846));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer34 (.A(net846),
    .X(net847));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer35 (.A(net847),
    .X(net848));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer36 (.A(net84),
    .X(net849));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer37 (.A(net849),
    .X(net850));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer38 (.A(net850),
    .X(net851));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer39 (.A(net850),
    .X(net852));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer40 (.A(net80),
    .X(net853));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer41 (.A(net135),
    .X(net854));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer42 (.A(net79),
    .X(net855));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer43 (.A(net81),
    .X(net856));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer44 (.A(net856),
    .X(net857));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer45 (.A(net857),
    .X(net858));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer46 (.A(net856),
    .X(net859));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer47 (.A(net81),
    .X(net860));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer48 (.A(net759),
    .X(net861));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer49 (.A(net807),
    .X(net862));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer50 (.A(net729),
    .X(net863));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer51 (.A(net863),
    .X(net864));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(net646),
    .X(net865));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(net275),
    .X(net866));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(net383),
    .X(net867));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(net657),
    .X(net868));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(net632),
    .X(net869));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(net546),
    .X(net870));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(net656),
    .X(net871));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(net348),
    .X(net872));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(net368),
    .X(net873));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(net422),
    .X(net874));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(net238),
    .X(net875));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(net497),
    .X(net876));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(net430),
    .X(net877));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(net359),
    .X(net878));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(net382),
    .X(net879));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(net494),
    .X(net880));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(net149),
    .X(net881));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(net673),
    .X(net882));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(net628),
    .X(net883));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(net520),
    .X(net884));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(net349),
    .X(net885));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(net161),
    .X(net886));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(net164),
    .X(net887));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(net659),
    .X(net888));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(net274),
    .X(net889));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(net647),
    .X(net890));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(net776),
    .X(net891));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(net251),
    .X(net892));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(net311),
    .X(net893));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(net620),
    .X(net894));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(net542),
    .X(net895));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(net232),
    .X(net896));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(net283),
    .X(net897));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(net328),
    .X(net898));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(net518),
    .X(net899));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(net148),
    .X(net900));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(net444),
    .X(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_A (.DIODE(clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(in0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(in1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(in10));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(in11));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(in12));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(in13));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(in14));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(in15));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(in16));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(in17));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(in18));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(in19));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(in2));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(in20));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(in21));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(in22));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(in23));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(in24));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(in25));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(in26));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(in27));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_A (.DIODE(in28));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_A (.DIODE(in29));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_A (.DIODE(in3));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_A (.DIODE(in30));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_A (.DIODE(in31));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_A (.DIODE(in32));
 sky130_fd_sc_hd__diode_2 ANTENNA_input28_A (.DIODE(in33));
 sky130_fd_sc_hd__diode_2 ANTENNA_input29_A (.DIODE(in34));
 sky130_fd_sc_hd__diode_2 ANTENNA_input30_A (.DIODE(in35));
 sky130_fd_sc_hd__diode_2 ANTENNA_input31_A (.DIODE(in36));
 sky130_fd_sc_hd__diode_2 ANTENNA_input32_A (.DIODE(in37));
 sky130_fd_sc_hd__diode_2 ANTENNA_input33_A (.DIODE(in38));
 sky130_fd_sc_hd__diode_2 ANTENNA_input34_A (.DIODE(in39));
 sky130_fd_sc_hd__diode_2 ANTENNA_input35_A (.DIODE(in4));
 sky130_fd_sc_hd__diode_2 ANTENNA_input36_A (.DIODE(in40));
 sky130_fd_sc_hd__diode_2 ANTENNA_input37_A (.DIODE(in41));
 sky130_fd_sc_hd__diode_2 ANTENNA_input38_A (.DIODE(in42));
 sky130_fd_sc_hd__diode_2 ANTENNA_input39_A (.DIODE(in43));
 sky130_fd_sc_hd__diode_2 ANTENNA_input40_A (.DIODE(in44));
 sky130_fd_sc_hd__diode_2 ANTENNA_input41_A (.DIODE(in45));
 sky130_fd_sc_hd__diode_2 ANTENNA_input42_A (.DIODE(in46));
 sky130_fd_sc_hd__diode_2 ANTENNA_input43_A (.DIODE(in47));
 sky130_fd_sc_hd__diode_2 ANTENNA_input44_A (.DIODE(in48));
 sky130_fd_sc_hd__diode_2 ANTENNA_input45_A (.DIODE(in49));
 sky130_fd_sc_hd__diode_2 ANTENNA_input46_A (.DIODE(in5));
 sky130_fd_sc_hd__diode_2 ANTENNA_input47_A (.DIODE(in50));
 sky130_fd_sc_hd__diode_2 ANTENNA_input48_A (.DIODE(in51));
 sky130_fd_sc_hd__diode_2 ANTENNA_input49_A (.DIODE(in52));
 sky130_fd_sc_hd__diode_2 ANTENNA_input50_A (.DIODE(in53));
 sky130_fd_sc_hd__diode_2 ANTENNA_input51_A (.DIODE(in54));
 sky130_fd_sc_hd__diode_2 ANTENNA_input52_A (.DIODE(in55));
 sky130_fd_sc_hd__diode_2 ANTENNA_input53_A (.DIODE(in56));
 sky130_fd_sc_hd__diode_2 ANTENNA_input54_A (.DIODE(in57));
 sky130_fd_sc_hd__diode_2 ANTENNA_input55_A (.DIODE(in58));
 sky130_fd_sc_hd__diode_2 ANTENNA_input56_A (.DIODE(in59));
 sky130_fd_sc_hd__diode_2 ANTENNA_input57_A (.DIODE(in6));
 sky130_fd_sc_hd__diode_2 ANTENNA_input58_A (.DIODE(in60));
 sky130_fd_sc_hd__diode_2 ANTENNA_input59_A (.DIODE(in61));
 sky130_fd_sc_hd__diode_2 ANTENNA_input60_A (.DIODE(in7));
 sky130_fd_sc_hd__diode_2 ANTENNA_input61_A (.DIODE(in8));
 sky130_fd_sc_hd__diode_2 ANTENNA_input62_A (.DIODE(in9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_A0 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_RESET_B (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_A2 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_A2 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c182_B1_N (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_Y (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A0 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_S1 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_A2 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_B1 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_A3 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_B1 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_c190_A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_Y (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge758_SCD (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_A1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c184_A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c183_Y (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_A2 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_X (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c245_A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_A3 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_B (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_A2 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_X (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge765_SCE (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_A1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_S1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_B (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_B (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_X (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c502_B1_N (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_A0 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_B (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_B1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c198_Y (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c208_A (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_B (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_Y (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_A1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_c350_A1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_B (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_c203_Y (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_B (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_A4 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA_c218_A2 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA_c216_B1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_D (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA_c206_Y (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge760_RESET_B (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_c742_SET_B (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_D (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_SCD (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_SET_B (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_c216_X (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge763_D (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_c82_B (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_c77_Y (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_B1_N (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_c218_A4 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_A3 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_A (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_c229_A2 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_Y (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge759_SCD (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_A1 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_A1 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA_c239_SCE (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA_c235_X (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap123_A (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_A2 (.DIODE(net910));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_A1 (.DIODE(net910));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_A3 (.DIODE(net910));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_A2 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA_c269_Y (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA_c311_A (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_B (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA_c277_A1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA_c276_B (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA_c273_Y (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA_c665_A (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA_c278_A1 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA_c276_Y (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_A2 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_A1 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_B1_N (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_B (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_c283_B1_N (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_c277_X (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_A1 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_B (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_Y (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA_c64_X (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_A1 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_A2 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_SCE (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_A1 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_B1_N (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_c311_B (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_c109_A4 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_A1 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_A3 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_SET_B (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_B (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA_c297_B1_N (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_Y (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_A (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_SCE (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_Y (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge770_S0 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge768_RESET_B (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_D (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_SCD (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_Y (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_A1 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_B (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_SCE (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA_c313_B (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_X (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge778_SCD (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_A2 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_D (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_SCD (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_SCE (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_X (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA_c371_A3 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_A (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_c321_Q (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_c610_A1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_A3 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_A2 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_SCD (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_A2 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_A2 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c323_X (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_A1 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_A2 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_B (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_Q (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA_s781_D (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_X (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_A1 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_B1 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_c346_B (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_A (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_Y (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_B1 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_c615_SCE (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_B (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_c350_S0 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_Q_N (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_A2 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_c494_D (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_B (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_B (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_SCE (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_Q (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_D (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_B (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_B1_N (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_A2 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_Y (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge769_SCE (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_SET_B (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_A2 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_B1_N (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA_c372_B (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA_c371_S0 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_S0 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_B1_N (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_SCD (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_Y (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer11_A (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer10_A (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge779_RESET_B (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA_c400_Y (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap120_A (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge777_SCE (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA_c560_B (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA_c532_B (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_A2 (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_S1 (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA_c407_Y (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge757_SCE (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA_c723_A2 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA_c566_A3 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA_c530_B (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_B1_N (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA_c411_A (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA_c408_Y (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge757_SCD (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_SET_B (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_RESET_B (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_SCE (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA_c614_SET_B (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_SCD (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_A3 (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA_c434_SCD (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA_c409_Y (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_A0 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_B1_N (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_A1 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_RESET_B (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA_c411_B (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA_c410_Y (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_B1_N (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_A1 (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_Y (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA_c614_SCD (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_A1 (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_B1 (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_RESET_B (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_A2 (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_A2 (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA_c428_X (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout122_A (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge760_D (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_Y (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_SET_B (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_D (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_A4 (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_A2 (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_SCD (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_A0 (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_X (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge777_D (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_X (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge771_RESET_B (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_A1 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_S0 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_SET_B (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_SCE (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_S1 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_A3 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_A2 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_SET_B (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_Y (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge776_S0 (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge766_D (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_SCD (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_SCE (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_SET_B (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_SCD (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_X (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge773_A3 (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge771_SCE (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA_c458_X (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge759_RESET_B (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A2 (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_A1 (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_A2 (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_A3 (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA_c615_SET_B (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_S0 (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_Y (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_A0 (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_A3 (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_A2 (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_S1 (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_A3 (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_B1_N (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_B1_N (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_X (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_A2 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_A3 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_A4 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_B1_N (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_S0 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_Q (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_A3 (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_A (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA_c547_Y (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_A1 (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_S1 (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA_c739_A2 (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_B1_N (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_SCE (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_B1 (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA_c611_B1_N (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_S0 (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA_c564_A2 (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA_c562_Y (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_A4 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA_c633_A1 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_SCE (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_S0 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_A2 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_A2 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_A2 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA_c565_B (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA_c564_X (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_A0 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_A3 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_A2 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_c109_X (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_A1 (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_A3 (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_A1 (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_S0 (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA_c613_B1 (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_B1 (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_X (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_A2 (.DIODE(net513));
 sky130_fd_sc_hd__diode_2 ANTENNA_c678_A1 (.DIODE(net513));
 sky130_fd_sc_hd__diode_2 ANTENNA_c672_SET_B (.DIODE(net513));
 sky130_fd_sc_hd__diode_2 ANTENNA_c668_A2 (.DIODE(net513));
 sky130_fd_sc_hd__diode_2 ANTENNA_c665_Y (.DIODE(net513));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_A2 (.DIODE(net514));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_A1 (.DIODE(net514));
 sky130_fd_sc_hd__diode_2 ANTENNA_c671_SET_B (.DIODE(net514));
 sky130_fd_sc_hd__diode_2 ANTENNA_c669_B (.DIODE(net514));
 sky130_fd_sc_hd__diode_2 ANTENNA_c666_Y (.DIODE(net514));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_A1 (.DIODE(net517));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_B1_N (.DIODE(net517));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_B (.DIODE(net517));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_A3 (.DIODE(net517));
 sky130_fd_sc_hd__diode_2 ANTENNA_c677_B (.DIODE(net517));
 sky130_fd_sc_hd__diode_2 ANTENNA_c676_B (.DIODE(net517));
 sky130_fd_sc_hd__diode_2 ANTENNA_c670_SET_B (.DIODE(net517));
 sky130_fd_sc_hd__diode_2 ANTENNA_c669_Y (.DIODE(net517));
 sky130_fd_sc_hd__diode_2 ANTENNA_c263_S1 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_c261_B (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_c130_B (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_c127_A (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_c119_B (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_c118_B (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_c117_Y (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge776_A1 (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 ANTENNA_c739_A3 (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_SCE (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 ANTENNA_c676_Y (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 ANTENNA_c746_A2 (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA_c696_Y (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A1 (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_A2 (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_SCD (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA_c702_Q (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge776_S1 (.DIODE(net556));
 sky130_fd_sc_hd__diode_2 ANTENNA_c745_A3 (.DIODE(net556));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_A1 (.DIODE(net556));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_SCE (.DIODE(net556));
 sky130_fd_sc_hd__diode_2 ANTENNA_c723_A3 (.DIODE(net556));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_SCD (.DIODE(net556));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_A3 (.DIODE(net556));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_B (.DIODE(net556));
 sky130_fd_sc_hd__diode_2 ANTENNA_c703_X (.DIODE(net556));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge759_Q_N (.DIODE(net614));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_A (.DIODE(net614));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge777_Q (.DIODE(net640));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_A (.DIODE(net640));
 sky130_fd_sc_hd__diode_2 ANTENNA_s781_Q (.DIODE(net645));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_B1 (.DIODE(net645));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_B (.DIODE(net645));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_A (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_B (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_A (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c136_Y (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c545_B (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_c529_A (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_B1_N (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_B (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_c143_A1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_c140_Y (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge772_SCD (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_A2 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_A3 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_A0 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c743_A2 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c701_B1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_B (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c393_A1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_B (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_X (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_A2 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_A1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_c340_A (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_B (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_A2 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_B1_N (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_X (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_c70_Y (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_S0 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_A (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c215_A2 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c228_A2 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_A (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_Y (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_A0 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_B1_N (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_Y (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_c94_B (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c92_B (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c71_Y (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_A1 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_RESET_B (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_A2 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_SCE (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_B1_N (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_B (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_S0 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_A (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_B1_N (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_Y (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_A1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_c554_B (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_A2 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_Y (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_c267_A (.DIODE(net674));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_X (.DIODE(net674));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_SCE (.DIODE(net674));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_B1_N (.DIODE(net674));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_A1 (.DIODE(net674));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_A (.DIODE(net678));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_X (.DIODE(net678));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_A2 (.DIODE(net678));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_A (.DIODE(net678));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_SCD (.DIODE(net678));
 sky130_fd_sc_hd__diode_2 ANTENNA_c158_B (.DIODE(net678));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_X (.DIODE(net679));
 sky130_fd_sc_hd__diode_2 ANTENNA_c68_A (.DIODE(net679));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_A3 (.DIODE(net679));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_A1 (.DIODE(net679));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_X (.DIODE(net681));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_A (.DIODE(net681));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_B1_N (.DIODE(net681));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_X (.DIODE(net682));
 sky130_fd_sc_hd__diode_2 ANTENNA_c67_A (.DIODE(net682));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_A1 (.DIODE(net682));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_A (.DIODE(net682));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_X (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_A1 (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_B (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_A2 (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_B (.DIODE(net686));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_X (.DIODE(net686));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_A (.DIODE(net686));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_X (.DIODE(net688));
 sky130_fd_sc_hd__diode_2 ANTENNA_c206_B (.DIODE(net688));
 sky130_fd_sc_hd__diode_2 ANTENNA_c198_A (.DIODE(net688));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_A2 (.DIODE(net688));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_X (.DIODE(net691));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_A (.DIODE(net691));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_X (.DIODE(net696));
 sky130_fd_sc_hd__diode_2 ANTENNA_c69_A (.DIODE(net696));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_A (.DIODE(net696));
 sky130_fd_sc_hd__diode_2 ANTENNA_input30_X (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA_c97_B1_N (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA_c87_B1 (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA_c743_S0 (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA_c68_B (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_A1 (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_B1_N (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_A2 (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_B (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA_c253_A0 (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA_input32_X (.DIODE(net704));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge765_RESET_B (.DIODE(net704));
 sky130_fd_sc_hd__diode_2 ANTENNA_c98_B (.DIODE(net704));
 sky130_fd_sc_hd__diode_2 ANTENNA_c745_B1 (.DIODE(net704));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_A2 (.DIODE(net704));
 sky130_fd_sc_hd__diode_2 ANTENNA_c251_A3 (.DIODE(net704));
 sky130_fd_sc_hd__diode_2 ANTENNA_input33_X (.DIODE(net705));
 sky130_fd_sc_hd__diode_2 ANTENNA_c66_A (.DIODE(net705));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_S1 (.DIODE(net705));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_D (.DIODE(net705));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_B1_N (.DIODE(net705));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_B (.DIODE(net705));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_B (.DIODE(net705));
 sky130_fd_sc_hd__diode_2 ANTENNA_input36_X (.DIODE(net708));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge767_SCE (.DIODE(net708));
 sky130_fd_sc_hd__diode_2 ANTENNA_c695_B (.DIODE(net708));
 sky130_fd_sc_hd__diode_2 ANTENNA_c613_A1 (.DIODE(net708));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_S0 (.DIODE(net708));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_B1_N (.DIODE(net708));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_B1_N (.DIODE(net708));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_A3 (.DIODE(net708));
 sky130_fd_sc_hd__diode_2 ANTENNA_c251_A1 (.DIODE(net708));
 sky130_fd_sc_hd__diode_2 ANTENNA_c244_B (.DIODE(net708));
 sky130_fd_sc_hd__diode_2 ANTENNA_input43_X (.DIODE(net715));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge760_SET_B (.DIODE(net715));
 sky130_fd_sc_hd__diode_2 ANTENNA_c611_A1 (.DIODE(net715));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_A2 (.DIODE(net715));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_SCE (.DIODE(net715));
 sky130_fd_sc_hd__diode_2 ANTENNA_input45_X (.DIODE(net717));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_A1 (.DIODE(net717));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_B (.DIODE(net717));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_A3 (.DIODE(net717));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_B (.DIODE(net717));
 sky130_fd_sc_hd__diode_2 ANTENNA_input46_X (.DIODE(net718));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge773_A2 (.DIODE(net718));
 sky130_fd_sc_hd__diode_2 ANTENNA_c70_B (.DIODE(net718));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_SCD (.DIODE(net718));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_A2 (.DIODE(net718));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_A (.DIODE(net718));
 sky130_fd_sc_hd__diode_2 ANTENNA_c531_B (.DIODE(net718));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_B (.DIODE(net718));
 sky130_fd_sc_hd__diode_2 ANTENNA_c129_B1_N (.DIODE(net718));
 sky130_fd_sc_hd__diode_2 ANTENNA_input49_X (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA_c63_S1 (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA_c394_RESET_B (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_B (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_SCE (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_B (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA_c114_B (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA_c113_A (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA_input52_X (.DIODE(net724));
 sky130_fd_sc_hd__diode_2 ANTENNA_c64_S0 (.DIODE(net724));
 sky130_fd_sc_hd__diode_2 ANTENNA_c62_A1 (.DIODE(net724));
 sky130_fd_sc_hd__diode_2 ANTENNA_c251_S0 (.DIODE(net724));
 sky130_fd_sc_hd__diode_2 ANTENNA_c218_B1 (.DIODE(net724));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_A3 (.DIODE(net724));
 sky130_fd_sc_hd__diode_2 ANTENNA_c125_B (.DIODE(net724));
 sky130_fd_sc_hd__diode_2 ANTENNA_c111_B (.DIODE(net724));
 sky130_fd_sc_hd__diode_2 ANTENNA_input53_X (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_B1_N (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_A1 (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_A2 (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_A1 (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_B1_N (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_A4 (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_A2 (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer50_A (.DIODE(net729));
 sky130_fd_sc_hd__diode_2 ANTENNA_c134_A (.DIODE(net912));
 sky130_fd_sc_hd__diode_2 ANTENNA_input57_X (.DIODE(net912));
 sky130_fd_sc_hd__diode_2 ANTENNA_c398_B (.DIODE(net912));
 sky130_fd_sc_hd__diode_2 ANTENNA_c270_B (.DIODE(net912));
 sky130_fd_sc_hd__diode_2 ANTENNA_input62_X (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA_c78_B (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_S0 (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_RESET_B (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_B1_N (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_A2 (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA_c222_A (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA_output63_A (.DIODE(net735));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_SCE (.DIODE(net735));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_X (.DIODE(net735));
 sky130_fd_sc_hd__diode_2 ANTENNA_output64_A (.DIODE(net736));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_X (.DIODE(net736));
 sky130_fd_sc_hd__diode_2 ANTENNA_output67_A (.DIODE(net739));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge765_D (.DIODE(net739));
 sky130_fd_sc_hd__diode_2 ANTENNA_c340_Y (.DIODE(net739));
 sky130_fd_sc_hd__diode_2 ANTENNA_output68_A (.DIODE(net740));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_B1_N (.DIODE(net740));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_B1_N (.DIODE(net740));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_B1_N (.DIODE(net740));
 sky130_fd_sc_hd__diode_2 ANTENNA_c587_X (.DIODE(net740));
 sky130_fd_sc_hd__diode_2 ANTENNA_output69_A (.DIODE(net741));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge763_RESET_B (.DIODE(net741));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_SCD (.DIODE(net741));
 sky130_fd_sc_hd__diode_2 ANTENNA_c392_S0 (.DIODE(net741));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_SCD (.DIODE(net741));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_Y (.DIODE(net741));
 sky130_fd_sc_hd__diode_2 ANTENNA_output70_A (.DIODE(net742));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_A1 (.DIODE(net742));
 sky130_fd_sc_hd__diode_2 ANTENNA_c540_Q (.DIODE(net742));
 sky130_fd_sc_hd__diode_2 ANTENNA_output71_A (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge769_SCD (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_SET_B (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA_c373_A2 (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_X (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA_output74_A (.DIODE(net746));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_A3 (.DIODE(net746));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_A4 (.DIODE(net746));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_B (.DIODE(net746));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_B1_N (.DIODE(net746));
 sky130_fd_sc_hd__diode_2 ANTENNA_c295_X (.DIODE(net746));
 sky130_fd_sc_hd__diode_2 ANTENNA_output76_A (.DIODE(net748));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge760_SCE (.DIODE(net748));
 sky130_fd_sc_hd__diode_2 ANTENNA_c494_SCD (.DIODE(net748));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_SCE (.DIODE(net748));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_X (.DIODE(net748));
 sky130_fd_sc_hd__diode_2 ANTENNA_output81_A (.DIODE(net753));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_A2 (.DIODE(net753));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_S0 (.DIODE(net753));
 sky130_fd_sc_hd__diode_2 ANTENNA_c496_X (.DIODE(net753));
 sky130_fd_sc_hd__diode_2 ANTENNA_output84_A (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge763_SCE (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_A1 (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_A3 (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_SCD (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_Y (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA_output86_A (.DIODE(net758));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_S1 (.DIODE(net758));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_X (.DIODE(net758));
 sky130_fd_sc_hd__diode_2 ANTENNA_output88_A (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA_c494_SCE (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_RESET_B (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_Y (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA_output93_A (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_SCE (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_c393_A2 (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_c370_RESET_B (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_X (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_output95_A (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_c393_A3 (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_B (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_c183_B (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_Y (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_output97_A (.DIODE(net769));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_S1 (.DIODE(net769));
 sky130_fd_sc_hd__diode_2 ANTENNA_c238_SCE (.DIODE(net769));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_X (.DIODE(net769));
 sky130_fd_sc_hd__diode_2 ANTENNA_output98_A (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_B (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_A1 (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_Y (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout140_A (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout139_A (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_c270_Y (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_output103_A (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_A2 (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_B (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_Y (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold78_A (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_output104_A (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge773_S1 (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_B1 (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_SCD (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_B (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_A3 (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_SCE (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_B1 (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_X (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_output105_A (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_c263_S0 (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_c262_SCE (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_c258_B (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_c255_B (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_c253_A2 (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_c248_B (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_c246_Y (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_output110_A (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_c297_A2 (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_c257_B (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_X (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_output114_A (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_c392_A2 (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_c263_A3 (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_c262_SET_B (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_c257_Y (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_output117_A (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_A1 (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_c103_B (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_c101_Y (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_output118_A (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_A2 (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_A2 (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA_c241_B1_N (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA_c226_B (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_X (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA_output119_A (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_A3 (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_SCE (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_c395_A1 (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_c241_A2 (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_c198_B (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_X (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap120_X (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A0 (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_A3 (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_c558_B (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_c559_B1_N (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_c409_B (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout122_X (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_c613_A3 (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_SET_B (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_A3 (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_B1_N (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_A1 (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge775_SET_B (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_c561_SCE (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_B1 (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_c434_SCE (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_B1_N (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap126_X (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_B1_N (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_RESET_B (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_A2 (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_A (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout128_X (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_B1_N (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_B (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_A2 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_B1_N (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_SCE (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c613_A4 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_B1 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_SCD (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_B1_N (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_A (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout139_X (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_B1 (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_output100_A (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_B (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_c681_B1_N (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_S0 (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_S1 (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_B1_N (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_B1 (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_c278_B1_N (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_c277_B1 (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout140_X (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge759_SCE (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_A3 (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_c747_SCE (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_c723_A1 (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_SET_B (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_S1 (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_B1 (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_c369_B1_N (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_c364_B (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_A (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire141_X (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c159_B (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_B1 (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_A1 (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_15_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_14_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_13_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_12_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_11_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_10_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_9_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_8_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_7_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_6_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_5_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_4_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_3_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_2_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_1_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_0_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_X (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c557_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c561_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c563_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c571_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_CLK_N (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c698_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_CLK_N (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge760_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge771_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s781_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s798_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_6_0_clk_X (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_CLK_N (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge759_CLK_N (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge763_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge765_CLK_N (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge779_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s789_GATE_N (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s792_GATE_N (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_9_0_clk_X (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c237_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c238_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c239_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c262_CLK_N (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c394_CLK_N (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge767_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge778_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s780_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s785_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s786_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_10_0_clk_X (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer8_A (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_B (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_B (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer7_X (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_c661_B (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c669_A (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c667_B (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c543_B (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer22_X (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer37_A (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_B (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c234_A2 (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_B (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer36_X (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer51_A (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_A1 (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_B (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_c424_B1_N (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer50_X (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_SET_B (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold78_X (.DIODE(net891));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer52 (.A(net24),
    .X(net902));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer53 (.A(net902),
    .X(net903));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer54 (.A(net602),
    .X(net904));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer55 (.A(net797),
    .X(net905));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer56 (.A(net95),
    .X(net906));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer57 (.A(net906),
    .X(net907));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer58 (.A(net907),
    .X(net908));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer59 (.A(net126),
    .X(net909));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer60 (.A(net185),
    .X(net910));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer61 (.A(net185),
    .X(net911));
 sky130_fd_sc_hd__clkbuf_1 clone62 (.A(in6),
    .X(net912));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_266 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_483 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_303 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_403 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_435 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_476 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_283 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_311 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_284 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_338 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_479 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_456 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_357 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_431 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_488 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_443 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_553 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_163 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_339 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_172 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_476 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_484 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_354 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_102 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_495 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_86 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_609 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_123 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_247 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_403 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_5 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_25 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_95 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_163 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_87 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_456 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_247 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_87 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_102 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_146 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_5 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_143 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_230 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_617 ();
endmodule
