module netlist_1 (clk,
    in0,
    in1,
    in10,
    in11,
    in12,
    in13,
    in14,
    in15,
    in16,
    in17,
    in18,
    in19,
    in2,
    in20,
    in21,
    in22,
    in23,
    in24,
    in3,
    in4,
    in5,
    in6,
    in7,
    in8,
    in9,
    out0,
    out1,
    out10,
    out11,
    out12,
    out13,
    out14,
    out15,
    out16,
    out17,
    out18,
    out19,
    out2,
    out20,
    out21,
    out22,
    out23,
    out24,
    out3,
    out4,
    out5,
    out6,
    out7,
    out8,
    out9,
    rst);
 input clk;
 input in0;
 input in1;
 input in10;
 input in11;
 input in12;
 input in13;
 input in14;
 input in15;
 input in16;
 input in17;
 input in18;
 input in19;
 input in2;
 input in20;
 input in21;
 input in22;
 input in23;
 input in24;
 input in3;
 input in4;
 input in5;
 input in6;
 input in7;
 input in8;
 input in9;
 output out0;
 output out1;
 output out10;
 output out11;
 output out12;
 output out13;
 output out14;
 output out15;
 output out16;
 output out17;
 output out18;
 output out19;
 output out2;
 output out20;
 output out21;
 output out22;
 output out23;
 output out24;
 output out3;
 output out4;
 output out5;
 output out6;
 output out7;
 output out8;
 output out9;
 input rst;

 wire net0;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net629;
 wire net63;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net64;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net65;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net66;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net67;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net68;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net69;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net7;
 wire net70;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net71;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net72;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net73;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net74;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net75;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net76;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net77;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net78;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net79;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net8;
 wire net80;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net81;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net82;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net83;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net84;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net85;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net86;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net87;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net88;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net89;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net9;
 wire net90;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net91;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net92;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net93;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net94;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net95;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net96;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net97;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net98;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net99;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net556;
 wire net628;
 wire net759;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_0_net1020;
 wire clknet_1_0__leaf_net1020;
 wire clknet_1_1__leaf_net1020;
 wire clknet_0_net994;
 wire clknet_1_0__leaf_net994;
 wire clknet_1_1__leaf_net994;
 wire clknet_0_net558;
 wire clknet_1_0__leaf_net558;
 wire clknet_1_1__leaf_net558;
 wire clknet_0_net563;
 wire clknet_1_0__leaf_net563;
 wire clknet_1_1__leaf_net563;
 wire clknet_0_net993;
 wire clknet_1_0__leaf_net993;
 wire clknet_1_1__leaf_net993;
 wire clknet_0_net694;
 wire clknet_1_0__leaf_net694;
 wire clknet_1_1__leaf_net694;
 wire clknet_0_net949;
 wire clknet_1_0__leaf_net949;
 wire clknet_1_1__leaf_net949;
 wire clknet_0_net710;
 wire clknet_1_0__leaf_net710;
 wire clknet_1_1__leaf_net710;
 wire clknet_0_net717;
 wire clknet_1_0__leaf_net717;
 wire clknet_1_1__leaf_net717;
 wire clknet_0_net719;
 wire clknet_1_0__leaf_net719;
 wire clknet_1_1__leaf_net719;
 wire clknet_0_net712;
 wire clknet_1_0__leaf_net712;
 wire clknet_1_1__leaf_net712;
 wire clknet_0_net442;
 wire clknet_1_0__leaf_net442;
 wire clknet_1_1__leaf_net442;
 wire clknet_0_net447;
 wire clknet_1_0__leaf_net447;
 wire clknet_1_1__leaf_net447;
 wire clknet_0_net914;
 wire clknet_1_0__leaf_net914;
 wire clknet_1_1__leaf_net914;
 wire clknet_0_net985;
 wire clknet_1_0__leaf_net985;
 wire clknet_1_1__leaf_net985;
 wire clknet_0_net984;
 wire clknet_1_0__leaf_net984;
 wire clknet_1_1__leaf_net984;
 wire clknet_0_net498;
 wire clknet_1_0__leaf_net498;
 wire clknet_1_1__leaf_net498;
 wire clknet_0_net357;
 wire clknet_1_0__leaf_net357;
 wire clknet_1_1__leaf_net357;
 wire clknet_0_net197;
 wire clknet_1_0__leaf_net197;
 wire clknet_1_1__leaf_net197;
 wire clknet_0_net201;
 wire clknet_1_0__leaf_net201;
 wire clknet_1_1__leaf_net201;
 wire clknet_0_net85;
 wire clknet_1_0__leaf_net85;
 wire clknet_1_1__leaf_net85;
 wire clknet_0_net205;
 wire clknet_1_0__leaf_net205;
 wire clknet_1_1__leaf_net205;
 wire clknet_0_net208;
 wire clknet_1_0__leaf_net208;
 wire clknet_1_1__leaf_net208;
 wire clknet_0_net226;
 wire clknet_1_0__leaf_net226;
 wire clknet_1_1__leaf_net226;
 wire clknet_0_net210;
 wire clknet_1_0__leaf_net210;
 wire clknet_1_1__leaf_net210;
 wire clknet_0_net207;
 wire clknet_1_0__leaf_net207;
 wire clknet_1_1__leaf_net207;
 wire clknet_0_net213;
 wire clknet_1_0__leaf_net213;
 wire clknet_1_1__leaf_net213;
 wire clknet_0_net87;
 wire clknet_1_0__leaf_net87;
 wire clknet_1_1__leaf_net87;
 wire clknet_0_net91;
 wire clknet_1_0__leaf_net91;
 wire clknet_1_1__leaf_net91;
 wire clknet_0_net89;
 wire clknet_1_0__leaf_net89;
 wire clknet_1_1__leaf_net89;
 wire clknet_0_net88;
 wire clknet_1_0__leaf_net88;
 wire clknet_1_1__leaf_net88;
 wire clknet_0_net95;
 wire clknet_1_0__leaf_net95;
 wire clknet_1_1__leaf_net95;
 wire clknet_0_net79;
 wire clknet_1_0__leaf_net79;
 wire clknet_1_1__leaf_net79;
 wire clknet_0_net81;
 wire clknet_1_0__leaf_net81;
 wire clknet_1_1__leaf_net81;
 wire clknet_0_net951;
 wire clknet_1_0__leaf_net951;
 wire clknet_1_1__leaf_net951;
 wire clknet_0_net42;
 wire clknet_1_0__leaf_net42;
 wire clknet_1_1__leaf_net42;
 wire clknet_0_net29;
 wire clknet_1_0__leaf_net29;
 wire clknet_1_1__leaf_net29;
 wire clknet_0_net912;
 wire clknet_1_0__leaf_net912;
 wire clknet_1_1__leaf_net912;
 wire clknet_0_net26;
 wire clknet_1_0__leaf_net26;
 wire clknet_1_1__leaf_net26;
 wire clknet_0_net21;
 wire clknet_1_0__leaf_net21;
 wire clknet_1_1__leaf_net21;
 wire clknet_0_net24;
 wire clknet_1_0__leaf_net24;
 wire clknet_1_1__leaf_net24;
 wire clknet_0_net20;
 wire clknet_1_0__leaf_net20;
 wire clknet_1_1__leaf_net20;
 wire clknet_0_net25;
 wire clknet_1_0__leaf_net25;
 wire clknet_1_1__leaf_net25;
 wire clknet_0_net23;
 wire clknet_1_0__leaf_net23;
 wire clknet_1_1__leaf_net23;
 wire clknet_0_net34;
 wire clknet_1_0__leaf_net34;
 wire clknet_1_1__leaf_net34;
 wire clknet_0_net161;
 wire clknet_1_0__leaf_net161;
 wire clknet_1_1__leaf_net161;
 wire clknet_0_net163;
 wire clknet_1_0__leaf_net163;
 wire clknet_1_1__leaf_net163;
 wire clknet_0_net168;
 wire clknet_1_0__leaf_net168;
 wire clknet_1_1__leaf_net168;
 wire clknet_0_net162;
 wire clknet_1_0__leaf_net162;
 wire clknet_1_1__leaf_net162;
 wire clknet_0_net27;
 wire clknet_1_0__leaf_net27;
 wire clknet_1_1__leaf_net27;
 wire clknet_0_net22;
 wire clknet_1_0__leaf_net22;
 wire clknet_1_1__leaf_net22;
 wire clknet_0_net352;
 wire clknet_1_0__leaf_net352;
 wire clknet_1_1__leaf_net352;
 wire clknet_0_net353;
 wire clknet_1_0__leaf_net353;
 wire clknet_1_1__leaf_net353;
 wire clknet_0_net950;
 wire clknet_1_0__leaf_net950;
 wire clknet_1_1__leaf_net950;
 wire clknet_0_net764;
 wire clknet_1_0__leaf_net764;
 wire clknet_1_1__leaf_net764;
 wire clknet_0_net482;
 wire clknet_1_0__leaf_net482;
 wire clknet_1_1__leaf_net482;
 wire clknet_0_net479;
 wire clknet_1_0__leaf_net479;
 wire clknet_1_1__leaf_net479;
 wire clknet_0_net491;
 wire clknet_1_0__leaf_net491;
 wire clknet_1_1__leaf_net491;
 wire clknet_0_net496;
 wire clknet_1_0__leaf_net496;
 wire clknet_1_1__leaf_net496;
 wire clknet_0_net493;
 wire clknet_1_0__leaf_net493;
 wire clknet_1_1__leaf_net493;
 wire clknet_0_net747;
 wire clknet_1_0__leaf_net747;
 wire clknet_1_1__leaf_net747;
 wire clknet_0_net318;
 wire clknet_1_0__leaf_net318;
 wire clknet_1_1__leaf_net318;
 wire clknet_0_net325;
 wire clknet_1_0__leaf_net325;
 wire clknet_1_1__leaf_net325;
 wire clknet_0_net320;
 wire clknet_1_0__leaf_net320;
 wire clknet_1_1__leaf_net320;
 wire clknet_0_net321;
 wire clknet_1_0__leaf_net321;
 wire clknet_1_1__leaf_net321;
 wire clknet_0_net317;
 wire clknet_1_0__leaf_net317;
 wire clknet_1_1__leaf_net317;
 wire clknet_0_net324;
 wire clknet_1_0__leaf_net324;
 wire clknet_1_1__leaf_net324;
 wire clknet_0_net329;
 wire clknet_1_0__leaf_net329;
 wire clknet_1_1__leaf_net329;
 wire clknet_0_net326;
 wire clknet_1_0__leaf_net326;
 wire clknet_1_1__leaf_net326;
 wire clknet_0_net330;
 wire clknet_1_0__leaf_net330;
 wire clknet_1_1__leaf_net330;
 wire clknet_0_net328;
 wire clknet_1_0__leaf_net328;
 wire clknet_1_1__leaf_net328;
 wire clknet_0_net915;
 wire clknet_1_0__leaf_net915;
 wire clknet_1_1__leaf_net915;
 wire clknet_0_net160;
 wire clknet_1_0__leaf_net160;
 wire clknet_1_1__leaf_net160;
 wire clknet_0_net144;
 wire clknet_1_0__leaf_net144;
 wire clknet_1_1__leaf_net144;
 wire clknet_0_net147;
 wire clknet_1_0__leaf_net147;
 wire clknet_1_1__leaf_net147;
 wire clknet_0_net145;
 wire clknet_1_0__leaf_net145;
 wire clknet_1_1__leaf_net145;
 wire clknet_0_net272;
 wire clknet_1_0__leaf_net272;
 wire clknet_1_1__leaf_net272;
 wire clknet_0_net126;
 wire clknet_1_0__leaf_net126;
 wire clknet_1_1__leaf_net126;
 wire clknet_0_net129;
 wire clknet_1_0__leaf_net129;
 wire clknet_1_1__leaf_net129;
 wire clknet_0_net127;
 wire clknet_1_0__leaf_net127;
 wire clknet_1_1__leaf_net127;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;

 sky130_fd_sc_hd__and3_1 c100 (.A(net76),
    .B(net67),
    .C(net71),
    .X(net77));
 sky130_fd_sc_hd__and3_1 c101 (.A(net57),
    .B(net76),
    .C(net963),
    .X(net78));
 sky130_fd_sc_hd__and2_0 c102 (.A(net73),
    .B(clknet_1_1__leaf_net985),
    .X(net79));
 sky130_fd_sc_hd__and2_1 c103 (.A(net75),
    .B(net69),
    .X(net80));
 sky130_fd_sc_hd__and3_1 c104 (.A(net80),
    .B(net76),
    .C(clknet_1_1__leaf_net79),
    .X(net81));
 sky130_fd_sc_hd__mux4_1 c105 (.A0(net74),
    .A1(clknet_1_0__leaf_net79),
    .A2(net80),
    .A3(clknet_1_0__leaf_net81),
    .S0(net66),
    .S1(net43),
    .X(net82));
 sky130_fd_sc_hd__or4bb_1 c106 (.A(clknet_1_0__leaf_net79),
    .B(net80),
    .C_N(net76),
    .D_N(net67),
    .X(net83));
 sky130_fd_sc_hd__mux4_1 c107 (.A0(net72),
    .A1(net80),
    .A2(net43),
    .A3(net68),
    .S0(clknet_1_1__leaf_net985),
    .S1(net987),
    .X(net84));
 sky130_fd_sc_hd__buf_1 c108 (.A(clknet_1_0__leaf_net985),
    .X(net85));
 sky130_fd_sc_hd__clkbuf_1 c109 (.A(net1040),
    .X(net86));
 sky130_fd_sc_hd__buf_1 c110 (.A(clknet_1_0__leaf_net85),
    .X(net87));
 sky130_fd_sc_hd__and2_0 c111 (.A(clknet_1_0__leaf_net87),
    .B(net73),
    .X(net88));
 sky130_fd_sc_hd__and2_0 c112 (.A(clknet_1_0__leaf_net88),
    .B(clknet_1_0__leaf_net87),
    .X(net89));
 sky130_fd_sc_hd__clkbuf_1 c113 (.A(net910),
    .X(net90));
 sky130_fd_sc_hd__buf_1 c114 (.A(clknet_1_1__leaf_net87),
    .X(net91));
 sky130_fd_sc_hd__buf_1 c115 (.A(net73),
    .X(net92));
 sky130_fd_sc_hd__dlymetal6s2s_1 c116 (.A(net90),
    .X(net93));
 sky130_fd_sc_hd__and3_1 c117 (.A(net90),
    .B(clknet_1_0__leaf_net88),
    .C(net92),
    .X(net94));
 sky130_fd_sc_hd__and2_0 c118 (.A(clknet_1_1__leaf_net88),
    .B(net93),
    .X(net95));
 sky130_fd_sc_hd__and2_0 c119 (.A(net92),
    .B(net93),
    .X(net96));
 sky130_fd_sc_hd__buf_1 c120 (.A(net910),
    .X(net97));
 sky130_fd_sc_hd__dfbbn_1 c121 (.CLK_N(clknet_4_10_0_clk),
    .D(clknet_1_1__leaf_net89),
    .RESET_B(clknet_1_0__leaf_net95),
    .SET_B(net93),
    .Q(net99),
    .Q_N(net98));
 sky130_fd_sc_hd__dfbbn_1 c122 (.CLK_N(clknet_4_10_0_clk),
    .D(net1055),
    .RESET_B(net97),
    .SET_B(clknet_1_1__leaf_net95),
    .Q(net101),
    .Q_N(net100));
 sky130_fd_sc_hd__dfbbp_1 c123 (.CLK(clknet_4_10_0_clk),
    .D(clknet_1_0__leaf_net95),
    .RESET_B(net99),
    .SET_B(net92),
    .Q(net103),
    .Q_N(net102));
 sky130_fd_sc_hd__sdfxbp_1 c124 (.CLK(clknet_4_10_0_clk),
    .D(clknet_1_0__leaf_net95),
    .SCD(net98),
    .SCE(net101),
    .Q(net105),
    .Q_N(net104));
 sky130_fd_sc_hd__sdfrbp_1 c125 (.CLK(clknet_4_10_0_clk),
    .D(clknet_1_0__leaf_net91),
    .RESET_B(net1034),
    .SCD(net100),
    .SCE(clknet_1_1__leaf_net95),
    .Q(net107),
    .Q_N(net106));
 sky130_fd_sc_hd__and3_1 c126 (.A(net93),
    .B(net96),
    .C(net106),
    .X(net108));
 sky130_fd_sc_hd__sdfxbp_1 c127 (.CLK(clknet_4_10_0_clk),
    .D(net97),
    .SCD(net1056),
    .SCE(net108),
    .Q(net110),
    .Q_N(net109));
 sky130_fd_sc_hd__and3_1 c128 (.A(net107),
    .B(net108),
    .C(net109),
    .X(net111));
 sky130_fd_sc_hd__sdfbbn_1 c129 (.CLK_N(clknet_4_10_0_clk),
    .D(net105),
    .RESET_B(net110),
    .SCD(net97),
    .SCE(clknet_1_1__leaf_net95),
    .SET_B(net93),
    .Q(net113),
    .Q_N(net112));
 sky130_fd_sc_hd__and3_1 c130 (.A(net86),
    .B(net113),
    .C(net108),
    .X(net114));
 sky130_fd_sc_hd__a2111o_1 c131 (.A1(net96),
    .A2(net110),
    .B1(net112),
    .C1(net104),
    .D1(clknet_1_1__leaf_net95),
    .X(net115));
 sky130_fd_sc_hd__buf_2 c132 (.A(in18),
    .X(net116));
 sky130_fd_sc_hd__buf_1 c133 (.A(net116),
    .X(net117));
 sky130_fd_sc_hd__and3_1 c134 (.A(net117),
    .B(net1002),
    .C(net116),
    .X(net118));
 sky130_fd_sc_hd__and2_0 c135 (.A(net116),
    .B(net117),
    .X(net119));
 sky130_fd_sc_hd__clkbuf_1 c136 (.A(net907),
    .X(net120));
 sky130_fd_sc_hd__and2_0 c137 (.A(net116),
    .B(net120),
    .X(net121));
 sky130_fd_sc_hd__and2_1 c138 (.A(net117),
    .B(net116),
    .X(net122));
 sky130_fd_sc_hd__buf_1 c139 (.A(net907),
    .X(net123));
 sky130_fd_sc_hd__and3_1 c140 (.A(net121),
    .B(net123),
    .C(net116),
    .X(net124));
 sky130_fd_sc_hd__buf_1 c141 (.A(clknet_1_0__leaf_net915),
    .X(net125));
 sky130_fd_sc_hd__buf_1 c142 (.A(clknet_1_0__leaf_net915),
    .X(net126));
 sky130_fd_sc_hd__and3_1 c143 (.A(clknet_1_1__leaf_net126),
    .B(net116),
    .C(net121),
    .X(net127));
 sky130_fd_sc_hd__mux4_1 c144 (.A0(clknet_1_1__leaf_net127),
    .A1(net117),
    .A2(net122),
    .A3(clknet_1_0__leaf_net126),
    .S0(net116),
    .S1(net119),
    .X(net128));
 sky130_fd_sc_hd__and3_1 c145 (.A(net1011),
    .B(clknet_1_0__leaf_net126),
    .C(net870),
    .X(net129));
 sky130_fd_sc_hd__and3_2 c146 (.A(net120),
    .B(net1005),
    .C(net556),
    .X(net130));
 sky130_fd_sc_hd__buf_1 c147 (.A(net980),
    .X(net131));
 sky130_fd_sc_hd__clkbuf_1 c148 (.A(net976),
    .X(net132));
 sky130_fd_sc_hd__mux4_1 c149 (.A0(clknet_1_0__leaf_net129),
    .A1(net131),
    .A2(net130),
    .A3(net123),
    .S0(net116),
    .S1(clknet_1_1__leaf_net126),
    .X(net133));
 sky130_fd_sc_hd__clkbuf_1 c150 (.A(net932),
    .X(net134));
 sky130_fd_sc_hd__and3_1 c151 (.A(net996),
    .B(net132),
    .C(clknet_1_0__leaf_net126),
    .X(net135));
 sky130_fd_sc_hd__mux4_1 c152 (.A0(net133),
    .A1(net123),
    .A2(clknet_1_1__leaf_net129),
    .A3(clknet_1_1__leaf_net126),
    .S0(net130),
    .S1(net116),
    .X(net136));
 sky130_fd_sc_hd__and3_1 c153 (.A(net135),
    .B(net134),
    .C(net136),
    .X(net137));
 sky130_fd_sc_hd__buf_1 c154 (.A(net1006),
    .X(net138));
 sky130_fd_sc_hd__buf_1 c155 (.A(net138),
    .X(net139));
 sky130_fd_sc_hd__and2_2 c156 (.A(net139),
    .B(net138),
    .X(net140));
 sky130_fd_sc_hd__clkbuf_1 c157 (.A(net975),
    .X(net141));
 sky130_fd_sc_hd__and2_2 c158 (.A(net139),
    .B(net999),
    .X(net142));
 sky130_fd_sc_hd__clkbuf_1 c159 (.A(net975),
    .X(net143));
 sky130_fd_sc_hd__buf_1 c160 (.A(clknet_1_1__leaf_net915),
    .X(net144));
 sky130_fd_sc_hd__and2_0 c161 (.A(clknet_1_0__leaf_net144),
    .B(net138),
    .X(net145));
 sky130_fd_sc_hd__buf_1 c162 (.A(net916),
    .X(net146));
 sky130_fd_sc_hd__and3_1 c163 (.A(net143),
    .B(clknet_1_0__leaf_net144),
    .C(net146),
    .X(net147));
 sky130_fd_sc_hd__sdfbbp_1 c164 (.CLK(clknet_4_13_0_clk),
    .D(net146),
    .RESET_B(clknet_1_0__leaf_net147),
    .SCD(net139),
    .SCE(net142),
    .SET_B(net140),
    .Q(net149),
    .Q_N(net148));
 sky130_fd_sc_hd__buf_1 c165 (.A(clknet_1_1__leaf_net915),
    .X(net150));
 sky130_fd_sc_hd__and3_1 c166 (.A(net149),
    .B(net143),
    .C(clknet_1_1__leaf_net145),
    .X(net151));
 sky130_fd_sc_hd__clkbuf_1 c167 (.A(net957),
    .X(net152));
 sky130_fd_sc_hd__clkbuf_1 c168 (.A(net976),
    .X(net153));
 sky130_fd_sc_hd__mux4_1 c169 (.A0(clknet_1_1__leaf_net144),
    .A1(clknet_1_1__leaf_net147),
    .A2(net149),
    .A3(net138),
    .S0(net13),
    .S1(net139),
    .X(net154));
 sky130_fd_sc_hd__or4bb_1 c170 (.A(net153),
    .B(net146),
    .C_N(net148),
    .D_N(net142),
    .X(net155));
 sky130_fd_sc_hd__and3_1 c171 (.A(net141),
    .B(net146),
    .C(net938),
    .X(net156));
 sky130_fd_sc_hd__mux4_1 c172 (.A0(clknet_1_0__leaf_net147),
    .A1(net153),
    .A2(net138),
    .A3(net140),
    .S0(net142),
    .S1(net938),
    .X(net157));
 sky130_fd_sc_hd__and3_1 c173 (.A(net150),
    .B(net156),
    .C(net153),
    .X(net158));
 sky130_fd_sc_hd__and2_0 c174 (.A(net156),
    .B(net907),
    .X(net159));
 sky130_fd_sc_hd__and3_1 c175 (.A(net158),
    .B(net159),
    .C(net146),
    .X(net160));
 sky130_fd_sc_hd__and2_0 c176 (.A(clknet_1_1__leaf_net42),
    .B(net948),
    .X(net161));
 sky130_fd_sc_hd__and2_0 c177 (.A(clknet_1_1__leaf_net145),
    .B(clknet_1_0__leaf_net161),
    .X(net162));
 sky130_fd_sc_hd__and2_0 c178 (.A(net1015),
    .B(clknet_1_1__leaf_net161),
    .X(net163));
 sky130_fd_sc_hd__clkbuf_1 c179 (.A(net904),
    .X(net164));
 sky130_fd_sc_hd__buf_1 c180 (.A(net904),
    .X(net165));
 sky130_fd_sc_hd__buf_1 c181 (.A(net976),
    .X(net166));
 sky130_fd_sc_hd__and2_0 c182 (.A(net166),
    .B(net165),
    .X(net167));
 sky130_fd_sc_hd__and2_0 c183 (.A(clknet_1_0__leaf_net163),
    .B(net166),
    .X(net168));
 sky130_fd_sc_hd__and2_0 c184 (.A(net167),
    .B(clknet_1_0__leaf_net163),
    .X(net169));
 sky130_fd_sc_hd__clkbuf_1 c185 (.A(net942),
    .X(net170));
 sky130_fd_sc_hd__buf_1 c186 (.A(net947),
    .X(net171));
 sky130_fd_sc_hd__and3_1 c187 (.A(clknet_1_1__leaf_net168),
    .B(net166),
    .C(net165),
    .X(net172));
 sky130_fd_sc_hd__mux4_1 c188 (.A0(clknet_1_1__leaf_net163),
    .A1(clknet_1_1__leaf_net168),
    .A2(net171),
    .A3(net165),
    .S0(net166),
    .S1(net904),
    .X(net173));
 sky130_fd_sc_hd__a2111o_1 c189 (.A1(net171),
    .A2(net166),
    .B1(clknet_1_1__leaf_net163),
    .C1(clknet_1_1__leaf_net162),
    .D1(net904),
    .X(net174));
 sky130_fd_sc_hd__clkbuf_1 c190 (.A(net954),
    .X(net175));
 sky130_fd_sc_hd__and3_1 c191 (.A(net166),
    .B(net170),
    .C(net171),
    .X(net176));
 sky130_fd_sc_hd__and2_0 c192 (.A(net170),
    .B(net171),
    .X(net177));
 sky130_fd_sc_hd__and2_0 c193 (.A(net164),
    .B(net177),
    .X(net178));
 sky130_fd_sc_hd__clkbuf_1 c194 (.A(net947),
    .X(net179));
 sky130_fd_sc_hd__and2_0 c195 (.A(net175),
    .B(net179),
    .X(net180));
 sky130_fd_sc_hd__and2_0 c196 (.A(net177),
    .B(net180),
    .X(net181));
 sky130_fd_sc_hd__and2_0 c197 (.A(clknet_1_1__leaf_net161),
    .B(net178),
    .X(net182));
 sky130_fd_sc_hd__clkbuf_2 c198 (.A(net930),
    .X(net183));
 sky130_fd_sc_hd__buf_1 c199 (.A(net183),
    .X(net184));
 sky130_fd_sc_hd__clkbuf_1 c200 (.A(net930),
    .X(net185));
 sky130_fd_sc_hd__clkbuf_1 c201 (.A(net183),
    .X(net186));
 sky130_fd_sc_hd__and2_2 c202 (.A(net186),
    .B(net183),
    .X(net187));
 sky130_fd_sc_hd__and2_0 c203 (.A(net185),
    .B(net187),
    .X(net188));
 sky130_fd_sc_hd__and2_0 c204 (.A(net43),
    .B(net187),
    .X(net189));
 sky130_fd_sc_hd__and2_0 c205 (.A(net186),
    .B(net183),
    .X(net190));
 sky130_fd_sc_hd__and2_0 c206 (.A(net184),
    .B(net183),
    .X(net191));
 sky130_fd_sc_hd__buf_1 c207 (.A(net944),
    .X(net192));
 sky130_fd_sc_hd__and2_1 c208 (.A(net187),
    .B(net882),
    .X(net193));
 sky130_fd_sc_hd__clkbuf_1 c209 (.A(net974),
    .X(net194));
 sky130_fd_sc_hd__and2_0 c210 (.A(net192),
    .B(net882),
    .X(net195));
 sky130_fd_sc_hd__or4bb_1 c211 (.A(net187),
    .B(net193),
    .C_N(clknet_1_1__leaf_net42),
    .D_N(net183),
    .X(net196));
 sky130_fd_sc_hd__buf_1 c212 (.A(clknet_1_1__leaf_net984),
    .X(net197));
 sky130_fd_sc_hd__and3_1 c213 (.A(net193),
    .B(clknet_1_0__leaf_net197),
    .C(net979),
    .X(net198));
 sky130_fd_sc_hd__clkbuf_1 c214 (.A(net942),
    .X(net199));
 sky130_fd_sc_hd__or4bb_1 c215 (.A(net194),
    .B(net186),
    .C_N(clknet_1_0__leaf_net197),
    .D_N(net183),
    .X(net200));
 sky130_fd_sc_hd__and3_1 c216 (.A(net200),
    .B(net199),
    .C(clknet_1_1__leaf_net197),
    .X(net201));
 sky130_fd_sc_hd__a2111o_1 c217 (.A1(net195),
    .A2(net192),
    .B1(clknet_1_1__leaf_net201),
    .C1(net199),
    .D1(net979),
    .X(net202));
 sky130_fd_sc_hd__clkbuf_1 c218 (.A(net974),
    .X(net203));
 sky130_fd_sc_hd__a2111o_1 c219 (.A1(net203),
    .A2(net192),
    .B1(clknet_1_0__leaf_net201),
    .C1(net187),
    .D1(net956),
    .X(net204));
 sky130_fd_sc_hd__buf_1 c220 (.A(clknet_1_1__leaf_net85),
    .X(net205));
 sky130_fd_sc_hd__buf_1 c221 (.A(net771),
    .X(net206));
 sky130_fd_sc_hd__and2_0 c222 (.A(net206),
    .B(clknet_1_0__leaf_net205),
    .X(net207));
 sky130_fd_sc_hd__and2_0 c223 (.A(clknet_1_0__leaf_net205),
    .B(net206),
    .X(net208));
 sky130_fd_sc_hd__buf_1 c224 (.A(clknet_1_1__leaf_net207),
    .X(net209));
 sky130_fd_sc_hd__and2_0 c225 (.A(clknet_1_0__leaf_net208),
    .B(net987),
    .X(net210));
 sky130_fd_sc_hd__and2_0 c226 (.A(clknet_1_1__leaf_net205),
    .B(clknet_1_0__leaf_net207),
    .X(net211));
 sky130_fd_sc_hd__and3_1 c227 (.A(net206),
    .B(clknet_1_0__leaf_net208),
    .C(clknet_1_0__leaf_net210),
    .X(net212));
 sky130_fd_sc_hd__and2_0 c228 (.A(clknet_1_0__leaf_net207),
    .B(net206),
    .X(net213));
 sky130_fd_sc_hd__clkbuf_1 c229 (.A(net771),
    .X(net214));
 sky130_fd_sc_hd__clkbuf_1 c230 (.A(net778),
    .X(net215));
 sky130_fd_sc_hd__buf_1 c231 (.A(net809),
    .X(net216));
 sky130_fd_sc_hd__and2_0 c232 (.A(net215),
    .B(net216),
    .X(net217));
 sky130_fd_sc_hd__and2_0 c233 (.A(net206),
    .B(net214),
    .X(net218));
 sky130_fd_sc_hd__and2_0 c234 (.A(net216),
    .B(net218),
    .X(net219));
 sky130_fd_sc_hd__and2_0 c235 (.A(net217),
    .B(net216),
    .X(net220));
 sky130_fd_sc_hd__and3_1 c236 (.A(net214),
    .B(net220),
    .C(net879),
    .X(net221));
 sky130_fd_sc_hd__sdfxtp_1 c237 (.CLK(clknet_4_14_0_clk),
    .D(net218),
    .SCD(net221),
    .SCE(clknet_1_1__leaf_net208),
    .Q(net222));
 sky130_fd_sc_hd__and3_1 c238 (.A(net220),
    .B(net1045),
    .C(net221),
    .X(net223));
 sky130_fd_sc_hd__or4bb_1 c239 (.A(net209),
    .B(net1045),
    .C_N(net221),
    .D_N(net220),
    .X(net224));
 sky130_fd_sc_hd__and3_1 c240 (.A(net216),
    .B(net221),
    .C(net942),
    .X(net225));
 sky130_fd_sc_hd__or4bb_1 c241 (.A(clknet_1_1__leaf_net208),
    .B(net222),
    .C_N(net878),
    .D_N(net901),
    .X(net226));
 sky130_fd_sc_hd__buf_1 c242 (.A(net959),
    .X(net227));
 sky130_fd_sc_hd__and2_2 c243 (.A(net227),
    .B(net100),
    .X(net228));
 sky130_fd_sc_hd__and2_1 c244 (.A(net227),
    .B(net959),
    .X(net229));
 sky130_fd_sc_hd__and2_0 c245 (.A(net228),
    .B(net229),
    .X(net230));
 sky130_fd_sc_hd__and2_1 c246 (.A(net1065),
    .B(net228),
    .X(net231));
 sky130_fd_sc_hd__clkbuf_2 c247 (.A(net909),
    .X(net232));
 sky130_fd_sc_hd__clkbuf_1 c248 (.A(net909),
    .X(net233));
 sky130_fd_sc_hd__buf_1 c249 (.A(net928),
    .X(net234));
 sky130_fd_sc_hd__and2_1 c25 (.A(net1008),
    .B(net1006),
    .X(net0));
 sky130_fd_sc_hd__sdfxtp_1 c250 (.CLK(clknet_4_11_0_clk),
    .D(net230),
    .SCD(net232),
    .SCE(net234),
    .Q(net235));
 sky130_fd_sc_hd__and2_0 c251 (.A(net235),
    .B(net233),
    .X(net236));
 sky130_fd_sc_hd__and2_0 c252 (.A(net236),
    .B(net233),
    .X(net237));
 sky130_fd_sc_hd__a2111o_1 c253 (.A1(net103),
    .A2(net1051),
    .B1(net234),
    .C1(net231),
    .D1(net227),
    .X(net238));
 sky130_fd_sc_hd__sdfrtn_1 c254 (.CLK_N(clknet_4_10_0_clk),
    .D(net237),
    .RESET_B(net1044),
    .SCD(net231),
    .SCE(net959),
    .Q(net239));
 sky130_fd_sc_hd__sdfrtp_1 c255 (.CLK(clknet_4_10_0_clk),
    .D(net237),
    .RESET_B(net231),
    .SCD(net232),
    .SCE(net234),
    .Q(net240));
 sky130_fd_sc_hd__and3_1 c256 (.A(net234),
    .B(net240),
    .C(net236),
    .X(net241));
 sky130_fd_sc_hd__and2_0 c257 (.A(net239),
    .B(net227),
    .X(net242));
 sky130_fd_sc_hd__and2_0 c258 (.A(net241),
    .B(net242),
    .X(net243));
 sky130_fd_sc_hd__and2_1 c259 (.A(net101),
    .B(net227),
    .X(net244));
 sky130_fd_sc_hd__and2_0 c26 (.A(net8),
    .B(net1009),
    .X(net1));
 sky130_fd_sc_hd__a2111o_1 c260 (.A1(net244),
    .A2(net232),
    .B1(net228),
    .C1(net229),
    .D1(net243),
    .X(net245));
 sky130_fd_sc_hd__mux4_1 c261 (.A0(net243),
    .A1(net244),
    .A2(net239),
    .A3(net228),
    .S0(net232),
    .S1(net888),
    .X(net246));
 sky130_fd_sc_hd__a2111o_1 c262 (.A1(net240),
    .A2(net235),
    .B1(net244),
    .C1(net228),
    .D1(net1063),
    .X(net247));
 sky130_fd_sc_hd__sdfbbn_1 c263 (.CLK_N(clknet_4_8_0_clk),
    .D(net247),
    .RESET_B(net241),
    .SCD(net244),
    .SCE(net889),
    .SET_B(net988),
    .Q(net249),
    .Q_N(net248));
 sky130_fd_sc_hd__buf_1 c264 (.A(net870),
    .X(net250));
 sky130_fd_sc_hd__clkbuf_2 c265 (.A(net250),
    .X(net251));
 sky130_fd_sc_hd__buf_1 c266 (.A(net251),
    .X(net252));
 sky130_fd_sc_hd__dlymetal6s2s_1 c267 (.A(net906),
    .X(net253));
 sky130_fd_sc_hd__buf_1 c268 (.A(net253),
    .X(net254));
 sky130_fd_sc_hd__and2_0 c269 (.A(net250),
    .B(net253),
    .X(net255));
 sky130_fd_sc_hd__and2_1 c27 (.A(net759),
    .B(net1006),
    .X(net2));
 sky130_fd_sc_hd__and2_0 c270 (.A(net255),
    .B(net253),
    .X(net256));
 sky130_fd_sc_hd__clkbuf_1 c271 (.A(net906),
    .X(net257));
 sky130_fd_sc_hd__buf_1 c272 (.A(net257),
    .X(net258));
 sky130_fd_sc_hd__and2_0 c273 (.A(net258),
    .B(net251),
    .X(net259));
 sky130_fd_sc_hd__and3_1 c274 (.A(net253),
    .B(net251),
    .C(net1001),
    .X(net260));
 sky130_fd_sc_hd__clkbuf_1 c275 (.A(net926),
    .X(net261));
 sky130_fd_sc_hd__and2_0 c276 (.A(net251),
    .B(net253),
    .X(net262));
 sky130_fd_sc_hd__clkbuf_1 c277 (.A(net1046),
    .X(net263));
 sky130_fd_sc_hd__clkbuf_2 c278 (.A(net925),
    .X(net264));
 sky130_fd_sc_hd__buf_1 c279 (.A(clknet_1_1__leaf_net994),
    .X(net265));
 sky130_fd_sc_hd__and3_1 c28 (.A(net1007),
    .B(net8),
    .C(net1000),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 c280 (.A(net925),
    .X(net266));
 sky130_fd_sc_hd__and3_1 c281 (.A(net266),
    .B(net255),
    .C(net264),
    .X(net267));
 sky130_fd_sc_hd__mux4_1 c282 (.A0(net265),
    .A1(net267),
    .A2(net260),
    .A3(net266),
    .S0(net251),
    .S1(net253),
    .X(net268));
 sky130_fd_sc_hd__and3_1 c283 (.A(net264),
    .B(net251),
    .C(net946),
    .X(net269));
 sky130_fd_sc_hd__and3_1 c284 (.A(net269),
    .B(net266),
    .C(net258),
    .X(net270));
 sky130_fd_sc_hd__and3_1 c285 (.A(net250),
    .B(net262),
    .C(net946),
    .X(net271));
 sky130_fd_sc_hd__and2_0 c286 (.A(net264),
    .B(clknet_1_0__leaf_net145),
    .X(net272));
 sky130_fd_sc_hd__buf_1 c287 (.A(net933),
    .X(net273));
 sky130_fd_sc_hd__and2_0 c288 (.A(net273),
    .B(net264),
    .X(net274));
 sky130_fd_sc_hd__clkbuf_1 c289 (.A(net933),
    .X(net275));
 sky130_fd_sc_hd__and2_0 c29 (.A(net2),
    .B(net0),
    .X(net4));
 sky130_fd_sc_hd__and2_1 c290 (.A(net275),
    .B(net273),
    .X(net276));
 sky130_fd_sc_hd__and2_1 c291 (.A(net254),
    .B(net276),
    .X(net277));
 sky130_fd_sc_hd__buf_1 c292 (.A(net277),
    .X(net278));
 sky130_fd_sc_hd__clkbuf_2 c293 (.A(net943),
    .X(net279));
 sky130_fd_sc_hd__sdfxtp_1 c294 (.CLK(clknet_4_5_0_clk),
    .D(net273),
    .SCD(net278),
    .SCE(net279),
    .Q(net280));
 sky130_fd_sc_hd__and2_0 c295 (.A(net277),
    .B(net273),
    .X(net281));
 sky130_fd_sc_hd__and3_1 c296 (.A(net276),
    .B(net277),
    .C(net280),
    .X(net282));
 sky130_fd_sc_hd__and2_0 c297 (.A(net280),
    .B(net279),
    .X(net283));
 sky130_fd_sc_hd__dlymetal6s2s_1 c298 (.A(net966),
    .X(net284));
 sky130_fd_sc_hd__clkbuf_1 c299 (.A(net926),
    .X(net285));
 sky130_fd_sc_hd__and3_1 c30 (.A(net1014),
    .B(net1004),
    .C(net998),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 c300 (.A(net941),
    .X(net286));
 sky130_fd_sc_hd__and3_1 c301 (.A(net286),
    .B(net279),
    .C(net284),
    .X(net287));
 sky130_fd_sc_hd__a2111o_1 c302 (.A1(net279),
    .A2(net278),
    .B1(net264),
    .C1(net287),
    .D1(net277),
    .X(net288));
 sky130_fd_sc_hd__and3_1 c303 (.A(net278),
    .B(net287),
    .C(net284),
    .X(net289));
 sky130_fd_sc_hd__and3_1 c304 (.A(net287),
    .B(net279),
    .C(net286),
    .X(net290));
 sky130_fd_sc_hd__mux4_1 c305 (.A0(net290),
    .A1(net286),
    .A2(net278),
    .A3(net279),
    .S0(net284),
    .S1(net977),
    .X(net291));
 sky130_fd_sc_hd__a2111o_1 c306 (.A1(net285),
    .A2(net280),
    .B1(net290),
    .C1(clknet_1_0__leaf_net272),
    .D1(net977),
    .X(net292));
 sky130_fd_sc_hd__sdfbbn_1 c307 (.CLK_N(clknet_4_6_0_clk),
    .D(net282),
    .RESET_B(net290),
    .SCD(net287),
    .SCE(net279),
    .SET_B(net906),
    .Q(net294),
    .Q_N(net293));
 sky130_fd_sc_hd__buf_1 c308 (.A(net876),
    .X(net295));
 sky130_fd_sc_hd__and2_1 c309 (.A(net295),
    .B(net294),
    .X(net296));
 sky130_fd_sc_hd__and2_0 c31 (.A(net5),
    .B(net2),
    .X(net6));
 sky130_fd_sc_hd__and2_1 c310 (.A(net295),
    .B(net293),
    .X(net297));
 sky130_fd_sc_hd__and2_1 c311 (.A(net297),
    .B(net295),
    .X(net298));
 sky130_fd_sc_hd__buf_1 c312 (.A(net875),
    .X(net299));
 sky130_fd_sc_hd__and2_1 c313 (.A(net297),
    .B(net298),
    .X(net300));
 sky130_fd_sc_hd__and2_0 c314 (.A(net296),
    .B(net299),
    .X(net301));
 sky130_fd_sc_hd__and2_2 c315 (.A(net298),
    .B(net956),
    .X(net302));
 sky130_fd_sc_hd__buf_1 c316 (.A(net916),
    .X(net303));
 sky130_fd_sc_hd__clkbuf_1 c317 (.A(net955),
    .X(net304));
 sky130_fd_sc_hd__buf_1 c318 (.A(net945),
    .X(net305));
 sky130_fd_sc_hd__and2_0 c319 (.A(net298),
    .B(net299),
    .X(net306));
 sky130_fd_sc_hd__or4bb_1 c32 (.A(net4),
    .B(net6),
    .C_N(net3),
    .D_N(net1006),
    .X(net7));
 sky130_fd_sc_hd__buf_1 c320 (.A(net966),
    .X(net307));
 sky130_fd_sc_hd__and3_1 c321 (.A(net299),
    .B(net303),
    .C(net293),
    .X(net308));
 sky130_fd_sc_hd__and3_1 c322 (.A(net308),
    .B(net296),
    .C(net295),
    .X(net309));
 sky130_fd_sc_hd__mux4_1 c323 (.A0(net303),
    .A1(net296),
    .A2(net308),
    .A3(net307),
    .S0(net302),
    .S1(net305),
    .X(net310));
 sky130_fd_sc_hd__and3_1 c324 (.A(net298),
    .B(net307),
    .C(net876),
    .X(net311));
 sky130_fd_sc_hd__clkbuf_1 c325 (.A(net973),
    .X(net312));
 sky130_fd_sc_hd__clkbuf_1 c326 (.A(net929),
    .X(net313));
 sky130_fd_sc_hd__mux4_1 c327 (.A0(net304),
    .A1(net309),
    .A2(net308),
    .A3(net313),
    .S0(net297),
    .S1(net302),
    .X(net314));
 sky130_fd_sc_hd__or4bb_1 c328 (.A(net312),
    .B(net297),
    .C_N(net313),
    .D_N(net990),
    .X(net315));
 sky130_fd_sc_hd__or4bb_1 c329 (.A(net315),
    .B(net313),
    .C_N(net301),
    .D_N(net990),
    .X(net316));
 sky130_fd_sc_hd__and2_1 c33 (.A(net1010),
    .B(net1003),
    .X(net8));
 sky130_fd_sc_hd__buf_1 c330 (.A(clknet_1_0__leaf_net747),
    .X(net317));
 sky130_fd_sc_hd__buf_1 c331 (.A(clknet_1_1__leaf_net747),
    .X(net318));
 sky130_fd_sc_hd__buf_1 c332 (.A(clknet_1_0__leaf_net318),
    .X(net319));
 sky130_fd_sc_hd__and2_0 c333 (.A(net319),
    .B(clknet_1_1__leaf_net317),
    .X(net320));
 sky130_fd_sc_hd__and2_0 c334 (.A(clknet_1_0__leaf_net320),
    .B(clknet_1_0__leaf_net317),
    .X(net321));
 sky130_fd_sc_hd__dlymetal6s2s_1 c335 (.A(net908),
    .X(net322));
 sky130_fd_sc_hd__clkbuf_1 c336 (.A(net923),
    .X(net323));
 sky130_fd_sc_hd__and2_0 c337 (.A(clknet_1_1__leaf_net317),
    .B(net956),
    .X(net324));
 sky130_fd_sc_hd__and2_0 c338 (.A(clknet_1_1__leaf_net320),
    .B(clknet_1_1__leaf_net318),
    .X(net325));
 sky130_fd_sc_hd__buf_1 c339 (.A(clknet_1_0__leaf_net950),
    .X(net326));
 sky130_fd_sc_hd__sdfrbp_1 c34 (.CLK(clknet_4_14_0_clk),
    .D(net0),
    .RESET_B(net7),
    .SCD(net2),
    .SCE(net1006),
    .Q(net10),
    .Q_N(net9));
 sky130_fd_sc_hd__and2_0 c340 (.A(clknet_1_0__leaf_net324),
    .B(clknet_1_0__leaf_net326),
    .X(net327));
 sky130_fd_sc_hd__and2_0 c341 (.A(net323),
    .B(clknet_1_0__leaf_net326),
    .X(net328));
 sky130_fd_sc_hd__and2_0 c342 (.A(net191),
    .B(clknet_1_1__leaf_net324),
    .X(net329));
 sky130_fd_sc_hd__and3_1 c343 (.A(clknet_1_1__leaf_net328),
    .B(clknet_1_1__leaf_net326),
    .C(net322),
    .X(net330));
 sky130_fd_sc_hd__clkbuf_1 c344 (.A(net935),
    .X(net331));
 sky130_fd_sc_hd__and2_0 c345 (.A(net322),
    .B(clknet_1_0__leaf_net328),
    .X(net332));
 sky130_fd_sc_hd__clkbuf_2 c346 (.A(net923),
    .X(net333));
 sky130_fd_sc_hd__clkbuf_1 c347 (.A(net856),
    .X(net334));
 sky130_fd_sc_hd__or4bb_1 c348 (.A(clknet_1_0__leaf_net318),
    .B(net334),
    .C_N(clknet_1_1__leaf_net330),
    .D_N(net322),
    .X(net335));
 sky130_fd_sc_hd__and3_1 c349 (.A(net331),
    .B(net332),
    .C(net333),
    .X(net336));
 sky130_fd_sc_hd__clkbuf_1 c35 (.A(net930),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 c350 (.A(net945),
    .X(net337));
 sky130_fd_sc_hd__or4bb_1 c351 (.A(net335),
    .B(net337),
    .C_N(net333),
    .D_N(clknet_1_1__leaf_net324),
    .X(net338));
 sky130_fd_sc_hd__dlymetal6s2s_1 c352 (.A(net948),
    .X(net339));
 sky130_fd_sc_hd__buf_1 c353 (.A(net339),
    .X(net340));
 sky130_fd_sc_hd__and2_0 c354 (.A(net340),
    .B(net339),
    .X(net341));
 sky130_fd_sc_hd__buf_1 c355 (.A(net948),
    .X(net342));
 sky130_fd_sc_hd__and2_0 c356 (.A(net342),
    .B(net340),
    .X(net343));
 sky130_fd_sc_hd__and2_1 c357 (.A(net340),
    .B(net342),
    .X(net344));
 sky130_fd_sc_hd__and2_1 c358 (.A(net342),
    .B(net343),
    .X(net345));
 sky130_fd_sc_hd__clkbuf_1 c359 (.A(net827),
    .X(net346));
 sky130_fd_sc_hd__and3_1 c36 (.A(net10),
    .B(net11),
    .C(net0),
    .X(net12));
 sky130_fd_sc_hd__buf_1 c360 (.A(net967),
    .X(net347));
 sky130_fd_sc_hd__mux4_1 c361 (.A0(net333),
    .A1(net345),
    .A2(net343),
    .A3(net347),
    .S0(net340),
    .S1(net339),
    .X(net348));
 sky130_fd_sc_hd__and3_1 c362 (.A(net347),
    .B(net344),
    .C(net333),
    .X(net349));
 sky130_fd_sc_hd__and2_0 c363 (.A(net341),
    .B(net342),
    .X(net350));
 sky130_fd_sc_hd__a2111o_1 c364 (.A1(net350),
    .A2(net344),
    .B1(net342),
    .C1(net346),
    .D1(net339),
    .X(net351));
 sky130_fd_sc_hd__buf_1 c365 (.A(clknet_1_1__leaf_net951),
    .X(net352));
 sky130_fd_sc_hd__and2_0 c366 (.A(net344),
    .B(clknet_1_0__leaf_net352),
    .X(net353));
 sky130_fd_sc_hd__and2_0 c367 (.A(clknet_1_1__leaf_net352),
    .B(net983),
    .X(net354));
 sky130_fd_sc_hd__or4bb_1 c368 (.A(net316),
    .B(clknet_1_0__leaf_net352),
    .C_N(clknet_1_0__leaf_net353),
    .D_N(net345),
    .X(net355));
 sky130_fd_sc_hd__and2_0 c369 (.A(net983),
    .B(clknet_1_0__leaf_net984),
    .X(net356));
 sky130_fd_sc_hd__and3_4 c37 (.A(net1),
    .B(net10),
    .C(net1006),
    .X(net13));
 sky130_fd_sc_hd__and2_0 c370 (.A(net356),
    .B(net340),
    .X(net357));
 sky130_fd_sc_hd__and2_0 c371 (.A(net354),
    .B(clknet_1_1__leaf_net357),
    .X(net358));
 sky130_fd_sc_hd__buf_1 c372 (.A(clknet_1_1__leaf_net984),
    .X(net359));
 sky130_fd_sc_hd__buf_1 c373 (.A(net778),
    .X(net360));
 sky130_fd_sc_hd__and2_0 c374 (.A(net228),
    .B(net989),
    .X(net361));
 sky130_fd_sc_hd__buf_2 c375 (.A(net229),
    .X(net362));
 sky130_fd_sc_hd__and2_0 c376 (.A(net339),
    .B(net232),
    .X(net363));
 sky130_fd_sc_hd__clkbuf_1 c377 (.A(net761),
    .X(net364));
 sky130_fd_sc_hd__and2_2 c378 (.A(net232),
    .B(net229),
    .X(net365));
 sky130_fd_sc_hd__buf_1 c379 (.A(net761),
    .X(net366));
 sky130_fd_sc_hd__or4bb_1 c38 (.A(net12),
    .B(net6),
    .C_N(net11),
    .D_N(net13),
    .X(net14));
 sky130_fd_sc_hd__buf_1 c380 (.A(clknet_1_1__leaf_net950),
    .X(net367));
 sky130_fd_sc_hd__and2_0 c381 (.A(net363),
    .B(net229),
    .X(net368));
 sky130_fd_sc_hd__clkbuf_1 c382 (.A(net980),
    .X(net369));
 sky130_fd_sc_hd__and3_1 c383 (.A(net362),
    .B(net361),
    .C(net364),
    .X(net370));
 sky130_fd_sc_hd__clkbuf_1 c384 (.A(net983),
    .X(net371));
 sky130_fd_sc_hd__or4bb_1 c385 (.A(net361),
    .B(net365),
    .C_N(net362),
    .D_N(net366),
    .X(net372));
 sky130_fd_sc_hd__and2_1 c386 (.A(net366),
    .B(net945),
    .X(net373));
 sky130_fd_sc_hd__and2_0 c387 (.A(net371),
    .B(net373),
    .X(net374));
 sky130_fd_sc_hd__buf_1 c388 (.A(clknet_1_0__leaf_net985),
    .X(net375));
 sky130_fd_sc_hd__clkbuf_1 c389 (.A(net827),
    .X(net376));
 sky130_fd_sc_hd__clkbuf_1 c39 (.A(net930),
    .X(net15));
 sky130_fd_sc_hd__and2_0 c390 (.A(net373),
    .B(net931),
    .X(net377));
 sky130_fd_sc_hd__and2_1 c391 (.A(net373),
    .B(net374),
    .X(net378));
 sky130_fd_sc_hd__a2111o_1 c392 (.A1(net374),
    .A2(net377),
    .B1(net378),
    .C1(net362),
    .D1(net373),
    .X(net379));
 sky130_fd_sc_hd__buf_1 c393 (.A(net940),
    .X(net380));
 sky130_fd_sc_hd__dfbbn_1 c394 (.CLK_N(clknet_4_9_0_clk),
    .D(net364),
    .RESET_B(net1068),
    .SET_B(net378),
    .Q(net382),
    .Q_N(net381));
 sky130_fd_sc_hd__mux4_1 c395 (.A0(net375),
    .A1(net380),
    .A2(net377),
    .A3(net382),
    .S0(net378),
    .S1(net362),
    .X(net383));
 sky130_fd_sc_hd__dlymetal6s2s_1 c396 (.A(net264),
    .X(net384));
 sky130_fd_sc_hd__clkbuf_1 c397 (.A(net384),
    .X(net385));
 sky130_fd_sc_hd__clkbuf_1 c398 (.A(net385),
    .X(net386));
 sky130_fd_sc_hd__clkbuf_1 c399 (.A(net756),
    .X(net387));
 sky130_fd_sc_hd__a2111o_1 c40 (.A1(net7),
    .A2(net628),
    .B1(net15),
    .C1(net12),
    .D1(net1042),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 c400 (.A(net756),
    .X(net388));
 sky130_fd_sc_hd__and2_1 c401 (.A(net385),
    .B(net388),
    .X(net389));
 sky130_fd_sc_hd__clkbuf_1 c402 (.A(net781),
    .X(net390));
 sky130_fd_sc_hd__and2_0 c403 (.A(net384),
    .B(net387),
    .X(net391));
 sky130_fd_sc_hd__and2_1 c404 (.A(net387),
    .B(net384),
    .X(net392));
 sky130_fd_sc_hd__clkbuf_1 c405 (.A(net392),
    .X(net393));
 sky130_fd_sc_hd__clkbuf_1 c406 (.A(net1032),
    .X(net394));
 sky130_fd_sc_hd__clkbuf_1 c407 (.A(net937),
    .X(net395));
 sky130_fd_sc_hd__clkbuf_1 c408 (.A(net1031),
    .X(net396));
 sky130_fd_sc_hd__and2_1 c409 (.A(net391),
    .B(net396),
    .X(net397));
 sky130_fd_sc_hd__mux4_1 c41 (.A0(net15),
    .A1(net12),
    .A2(net9),
    .A3(net13),
    .S0(net1007),
    .S1(net929),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 c410 (.A(net937),
    .X(net398));
 sky130_fd_sc_hd__and2_1 c411 (.A(net390),
    .B(net398),
    .X(net399));
 sky130_fd_sc_hd__clkbuf_1 c412 (.A(net936),
    .X(net400));
 sky130_fd_sc_hd__and3_1 c413 (.A(net396),
    .B(net399),
    .C(net388),
    .X(net401));
 sky130_fd_sc_hd__clkbuf_1 c414 (.A(net936),
    .X(net402));
 sky130_fd_sc_hd__and3_1 c415 (.A(net397),
    .B(net400),
    .C(net392),
    .X(net403));
 sky130_fd_sc_hd__and3_2 c416 (.A(net388),
    .B(net400),
    .C(net1059),
    .X(net404));
 sky130_fd_sc_hd__and3_1 c417 (.A(net391),
    .B(net401),
    .C(net399),
    .X(net405));
 sky130_fd_sc_hd__buf_1 c418 (.A(net294),
    .X(net406));
 sky130_fd_sc_hd__clkbuf_2 c419 (.A(net406),
    .X(net407));
 sky130_fd_sc_hd__a2111o_1 c42 (.A1(net8),
    .A2(net13),
    .B1(net1006),
    .C1(net929),
    .D1(net1042),
    .X(net18));
 sky130_fd_sc_hd__and2_0 c420 (.A(net407),
    .B(net406),
    .X(net408));
 sky130_fd_sc_hd__and2_0 c421 (.A(net404),
    .B(net407),
    .X(net409));
 sky130_fd_sc_hd__and2_0 c422 (.A(net284),
    .B(net407),
    .X(net410));
 sky130_fd_sc_hd__and2_2 c423 (.A(net402),
    .B(net406),
    .X(net411));
 sky130_fd_sc_hd__clkbuf_1 c424 (.A(net773),
    .X(net412));
 sky130_fd_sc_hd__and2_0 c425 (.A(net411),
    .B(net407),
    .X(net413));
 sky130_fd_sc_hd__and2_1 c426 (.A(net412),
    .B(net411),
    .X(net414));
 sky130_fd_sc_hd__clkbuf_1 c427 (.A(net773),
    .X(net415));
 sky130_fd_sc_hd__clkbuf_1 c428 (.A(net935),
    .X(net416));
 sky130_fd_sc_hd__or4bb_1 c429 (.A(net413),
    .B(net407),
    .C_N(net411),
    .D_N(net416),
    .X(net417));
 sky130_fd_sc_hd__and3_1 c43 (.A(net3),
    .B(net15),
    .C(net954),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_1 c430 (.A(net981),
    .X(net418));
 sky130_fd_sc_hd__and2_0 c431 (.A(net407),
    .B(net960),
    .X(net419));
 sky130_fd_sc_hd__and2_1 c432 (.A(net418),
    .B(net411),
    .X(net420));
 sky130_fd_sc_hd__and2_1 c433 (.A(net416),
    .B(net411),
    .X(net421));
 sky130_fd_sc_hd__clkbuf_1 c434 (.A(net1039),
    .X(net422));
 sky130_fd_sc_hd__and3_1 c435 (.A(net422),
    .B(net411),
    .C(net407),
    .X(net423));
 sky130_fd_sc_hd__buf_2 c436 (.A(net908),
    .X(net424));
 sky130_fd_sc_hd__clkbuf_1 c437 (.A(net807),
    .X(net425));
 sky130_fd_sc_hd__mux4_1 c438 (.A0(net425),
    .A1(net411),
    .A2(net423),
    .A3(net407),
    .S0(net424),
    .S1(net421),
    .X(net426));
 sky130_fd_sc_hd__mux4_1 c439 (.A0(net423),
    .A1(net414),
    .A2(net425),
    .A3(net420),
    .S0(net424),
    .S1(net960),
    .X(net427));
 sky130_fd_sc_hd__buf_1 c44 (.A(clknet_1_0__leaf_net42),
    .X(net20));
 sky130_fd_sc_hd__buf_1 c440 (.A(net991),
    .X(net428));
 sky130_fd_sc_hd__and2_0 c441 (.A(net428),
    .B(net990),
    .X(net429));
 sky130_fd_sc_hd__clkbuf_1 c442 (.A(net428),
    .X(net430));
 sky130_fd_sc_hd__and2_1 c443 (.A(net428),
    .B(net429),
    .X(net431));
 sky130_fd_sc_hd__buf_1 c444 (.A(net934),
    .X(net432));
 sky130_fd_sc_hd__clkbuf_1 c445 (.A(net934),
    .X(net433));
 sky130_fd_sc_hd__and2_1 c446 (.A(net432),
    .B(net430),
    .X(net434));
 sky130_fd_sc_hd__clkbuf_1 c447 (.A(net1054),
    .X(net435));
 sky130_fd_sc_hd__clkbuf_2 c448 (.A(net922),
    .X(net436));
 sky130_fd_sc_hd__clkbuf_1 c449 (.A(net871),
    .X(net437));
 sky130_fd_sc_hd__and2_0 c45 (.A(clknet_1_1__leaf_net20),
    .B(clknet_1_0__leaf_net42),
    .X(net21));
 sky130_fd_sc_hd__and3_1 c450 (.A(net437),
    .B(net431),
    .C(net428),
    .X(net438));
 sky130_fd_sc_hd__and2_1 c451 (.A(net429),
    .B(net437),
    .X(net439));
 sky130_fd_sc_hd__buf_1 c452 (.A(net958),
    .X(net440));
 sky130_fd_sc_hd__buf_1 c453 (.A(clknet_1_1__leaf_net949),
    .X(net441));
 sky130_fd_sc_hd__and3_1 c454 (.A(net441),
    .B(net440),
    .C(net436),
    .X(net442));
 sky130_fd_sc_hd__and2_0 c455 (.A(clknet_1_0__leaf_net442),
    .B(net440),
    .X(net443));
 sky130_fd_sc_hd__and3_1 c456 (.A(net436),
    .B(net440),
    .C(clknet_1_1__leaf_net442),
    .X(net444));
 sky130_fd_sc_hd__dfbbn_1 c457 (.CLK_N(clknet_4_3_0_clk),
    .D(net430),
    .RESET_B(net431),
    .SET_B(clknet_1_0__leaf_net442),
    .Q(net446),
    .Q_N(net445));
 sky130_fd_sc_hd__and3_1 c458 (.A(net444),
    .B(clknet_1_1__leaf_net442),
    .C(net446),
    .X(net447));
 sky130_fd_sc_hd__and3_1 c459 (.A(net446),
    .B(net436),
    .C(net440),
    .X(net448));
 sky130_fd_sc_hd__buf_1 c46 (.A(clknet_1_0__leaf_net951),
    .X(net22));
 sky130_fd_sc_hd__a2111o_1 c460 (.A1(clknet_1_0__leaf_net447),
    .A2(net448),
    .B1(clknet_1_1__leaf_net442),
    .C1(net436),
    .D1(net445),
    .X(net449));
 sky130_fd_sc_hd__mux4_1 c461 (.A0(net443),
    .A1(net431),
    .A2(clknet_1_1__leaf_net447),
    .A3(net434),
    .S0(net436),
    .S1(net957),
    .X(net450));
 sky130_fd_sc_hd__clkbuf_2 c462 (.A(net856),
    .X(net451));
 sky130_fd_sc_hd__clkbuf_1 c463 (.A(net451),
    .X(net452));
 sky130_fd_sc_hd__and2_1 c464 (.A(net452),
    .B(net1070),
    .X(net453));
 sky130_fd_sc_hd__buf_1 c465 (.A(net760),
    .X(net454));
 sky130_fd_sc_hd__clkbuf_2 c466 (.A(net760),
    .X(net455));
 sky130_fd_sc_hd__and3_1 c467 (.A(net440),
    .B(net455),
    .C(net451),
    .X(net456));
 sky130_fd_sc_hd__clkbuf_1 c468 (.A(net922),
    .X(net457));
 sky130_fd_sc_hd__and2_0 c469 (.A(net455),
    .B(net451),
    .X(net458));
 sky130_fd_sc_hd__and2_0 c47 (.A(net1013),
    .B(clknet_1_0__leaf_net20),
    .X(net23));
 sky130_fd_sc_hd__and2_0 c470 (.A(net452),
    .B(net957),
    .X(net459));
 sky130_fd_sc_hd__and2_2 c471 (.A(net455),
    .B(net454),
    .X(net460));
 sky130_fd_sc_hd__and2_1 c472 (.A(net458),
    .B(net460),
    .X(net461));
 sky130_fd_sc_hd__a2111o_1 c473 (.A1(net456),
    .A2(net457),
    .B1(net461),
    .C1(net454),
    .D1(net451),
    .X(net462));
 sky130_fd_sc_hd__clkbuf_1 c474 (.A(net917),
    .X(net463));
 sky130_fd_sc_hd__mux4_1 c475 (.A0(net452),
    .A1(net455),
    .A2(net461),
    .A3(net460),
    .S0(net333),
    .S1(net451),
    .X(net464));
 sky130_fd_sc_hd__clkbuf_1 c476 (.A(net944),
    .X(net465));
 sky130_fd_sc_hd__and2_0 c477 (.A(net465),
    .B(net965),
    .X(net466));
 sky130_fd_sc_hd__a2111o_1 c478 (.A1(net457),
    .A2(net455),
    .B1(net463),
    .C1(net456),
    .D1(net460),
    .X(net467));
 sky130_fd_sc_hd__and2_0 c479 (.A(net463),
    .B(net455),
    .X(net468));
 sky130_fd_sc_hd__and2_0 c48 (.A(clknet_1_0__leaf_net22),
    .B(clknet_1_1__leaf_net21),
    .X(net24));
 sky130_fd_sc_hd__mux4_1 c480 (.A0(net468),
    .A1(net463),
    .A2(net461),
    .A3(net456),
    .S0(net460),
    .S1(net455),
    .X(net469));
 sky130_fd_sc_hd__and2_0 c481 (.A(net466),
    .B(net939),
    .X(net470));
 sky130_fd_sc_hd__and3_1 c482 (.A(net454),
    .B(net470),
    .C(net460),
    .X(net471));
 sky130_fd_sc_hd__a2111o_1 c483 (.A1(net465),
    .A2(net470),
    .B1(net471),
    .C1(net467),
    .D1(net455),
    .X(net472));
 sky130_fd_sc_hd__buf_1 c484 (.A(net360),
    .X(net473));
 sky130_fd_sc_hd__clkbuf_1 c485 (.A(net473),
    .X(net474));
 sky130_fd_sc_hd__and2_0 c486 (.A(net474),
    .B(net360),
    .X(net475));
 sky130_fd_sc_hd__buf_1 c487 (.A(net473),
    .X(net476));
 sky130_fd_sc_hd__and2_0 c488 (.A(net476),
    .B(net473),
    .X(net477));
 sky130_fd_sc_hd__and2_1 c489 (.A(net473),
    .B(net476),
    .X(net478));
 sky130_fd_sc_hd__and2_0 c49 (.A(clknet_1_0__leaf_net20),
    .B(clknet_1_0__leaf_net23),
    .X(net25));
 sky130_fd_sc_hd__buf_1 c490 (.A(clknet_1_0__leaf_net764),
    .X(net479));
 sky130_fd_sc_hd__buf_1 c491 (.A(clknet_1_1__leaf_net764),
    .X(net480));
 sky130_fd_sc_hd__buf_2 c492 (.A(net966),
    .X(net481));
 sky130_fd_sc_hd__and3_1 c493 (.A(net480),
    .B(net481),
    .C(net476),
    .X(net482));
 sky130_fd_sc_hd__dfbbp_1 c494 (.CLK(clknet_4_6_0_clk),
    .D(net475),
    .RESET_B(clknet_1_1__leaf_net479),
    .SET_B(net473),
    .Q(net484),
    .Q_N(net483));
 sky130_fd_sc_hd__and3_1 c495 (.A(clknet_1_0__leaf_net482),
    .B(net481),
    .C(net474),
    .X(net485));
 sky130_fd_sc_hd__buf_1 c496 (.A(net967),
    .X(net486));
 sky130_fd_sc_hd__clkbuf_1 c497 (.A(net966),
    .X(net487));
 sky130_fd_sc_hd__buf_1 c498 (.A(net917),
    .X(net488));
 sky130_fd_sc_hd__clkbuf_1 c499 (.A(net923),
    .X(net489));
 sky130_fd_sc_hd__and2_0 c50 (.A(clknet_1_0__leaf_net42),
    .B(clknet_1_0__leaf_net20),
    .X(net26));
 sky130_fd_sc_hd__or4bb_1 c500 (.A(net489),
    .B(net484),
    .C_N(net360),
    .D_N(net488),
    .X(net490));
 sky130_fd_sc_hd__and3_1 c501 (.A(clknet_1_0__leaf_net479),
    .B(net487),
    .C(net490),
    .X(net491));
 sky130_fd_sc_hd__and3_1 c502 (.A(net467),
    .B(net487),
    .C(clknet_1_0__leaf_net482),
    .X(net492));
 sky130_fd_sc_hd__or4bb_1 c503 (.A(clknet_1_1__leaf_net491),
    .B(net486),
    .C_N(net481),
    .D_N(net943),
    .X(net493));
 sky130_fd_sc_hd__or4bb_1 c504 (.A(net490),
    .B(clknet_1_1__leaf_net493),
    .C_N(net488),
    .D_N(net473),
    .X(net494));
 sky130_fd_sc_hd__and3_1 c505 (.A(net487),
    .B(clknet_1_0__leaf_net493),
    .C(net490),
    .X(net495));
 sky130_fd_sc_hd__and2_0 c506 (.A(clknet_1_0__leaf_net491),
    .B(net481),
    .X(net496));
 sky130_fd_sc_hd__and2_0 c507 (.A(net481),
    .B(net381),
    .X(net497));
 sky130_fd_sc_hd__and2_0 c508 (.A(net481),
    .B(clknet_1_0__leaf_net984),
    .X(net498));
 sky130_fd_sc_hd__clkbuf_1 c509 (.A(net751),
    .X(net499));
 sky130_fd_sc_hd__buf_1 c51 (.A(clknet_1_0__leaf_net951),
    .X(net27));
 sky130_fd_sc_hd__buf_1 c510 (.A(net751),
    .X(net500));
 sky130_fd_sc_hd__and2_1 c511 (.A(net382),
    .B(net500),
    .X(net501));
 sky130_fd_sc_hd__and3_1 c512 (.A(net376),
    .B(clknet_1_0__leaf_net498),
    .C(net501),
    .X(net502));
 sky130_fd_sc_hd__and3_1 c513 (.A(clknet_1_1__leaf_net498),
    .B(net382),
    .C(net942),
    .X(net503));
 sky130_fd_sc_hd__and2_1 c514 (.A(net501),
    .B(net481),
    .X(net1026));
 sky130_fd_sc_hd__and2_0 c515 (.A(net500),
    .B(net501),
    .X(net504));
 sky130_fd_sc_hd__and3_1 c516 (.A(net504),
    .B(clknet_1_0__leaf_net496),
    .C(net501),
    .X(net505));
 sky130_fd_sc_hd__and2_0 c517 (.A(net502),
    .B(net499),
    .X(net506));
 sky130_fd_sc_hd__sdfxbp_1 c518 (.CLK(clknet_4_6_0_clk),
    .D(clknet_1_1__leaf_net498),
    .SCD(net500),
    .SCE(clknet_1_1__leaf_net496),
    .Q(net508),
    .Q_N(net507));
 sky130_fd_sc_hd__and2_1 c519 (.A(net497),
    .B(net504),
    .X(net509));
 sky130_fd_sc_hd__or4bb_1 c52 (.A(clknet_1_1__leaf_net24),
    .B(clknet_1_1__leaf_net22),
    .C_N(clknet_1_0__leaf_net27),
    .D_N(clknet_1_1__leaf_net20),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_2 c520 (.A(net973),
    .X(net510));
 sky130_fd_sc_hd__and3_1 c521 (.A(net509),
    .B(net508),
    .C(net510),
    .X(net511));
 sky130_fd_sc_hd__and3_1 c522 (.A(net503),
    .B(net507),
    .C(net509),
    .X(net512));
 sky130_fd_sc_hd__and3_1 c523 (.A(net500),
    .B(net509),
    .C(net965),
    .X(net513));
 sky130_fd_sc_hd__and3_1 c524 (.A(net506),
    .B(net510),
    .C(net504),
    .X(net514));
 sky130_fd_sc_hd__or4bb_1 c525 (.A(net501),
    .B(net509),
    .C_N(net481),
    .D_N(net958),
    .X(net515));
 sky130_fd_sc_hd__clkbuf_1 c526 (.A(net944),
    .X(net516));
 sky130_fd_sc_hd__and3_1 c527 (.A(net508),
    .B(net516),
    .C(net510),
    .X(net517));
 sky130_fd_sc_hd__buf_1 c528 (.A(net753),
    .X(net518));
 sky130_fd_sc_hd__buf_1 c529 (.A(net518),
    .X(net519));
 sky130_fd_sc_hd__and3_1 c53 (.A(clknet_1_0__leaf_net23),
    .B(clknet_1_0__leaf_net22),
    .C(clknet_1_0__leaf_net42),
    .X(net29));
 sky130_fd_sc_hd__and2_0 c530 (.A(net519),
    .B(net518),
    .X(net520));
 sky130_fd_sc_hd__and2_1 c531 (.A(net519),
    .B(net518),
    .X(net521));
 sky130_fd_sc_hd__and3_1 c532 (.A(net521),
    .B(net519),
    .C(net518),
    .X(net522));
 sky130_fd_sc_hd__buf_1 c533 (.A(net752),
    .X(net523));
 sky130_fd_sc_hd__and2_1 c534 (.A(net520),
    .B(net521),
    .X(net524));
 sky130_fd_sc_hd__buf_2 c535 (.A(net793),
    .X(net525));
 sky130_fd_sc_hd__and2_2 c536 (.A(net518),
    .B(net521),
    .X(net526));
 sky130_fd_sc_hd__buf_1 c537 (.A(net787),
    .X(net527));
 sky130_fd_sc_hd__sdfxbp_1 c538 (.CLK(clknet_4_0_0_clk),
    .D(net524),
    .SCD(net527),
    .SCE(net526),
    .Q(net529),
    .Q_N(net528));
 sky130_fd_sc_hd__sdfxtp_1 c539 (.CLK(clknet_4_0_0_clk),
    .D(net521),
    .SCD(net525),
    .SCE(net526),
    .Q(net530));
 sky130_fd_sc_hd__buf_1 c54 (.A(net923),
    .X(net30));
 sky130_fd_sc_hd__and3_1 c540 (.A(net518),
    .B(net527),
    .C(net525),
    .X(net531));
 sky130_fd_sc_hd__and3_1 c541 (.A(net523),
    .B(net1035),
    .C(net531),
    .X(net532));
 sky130_fd_sc_hd__and3_1 c542 (.A(net529),
    .B(net1035),
    .C(net520),
    .X(net533));
 sky130_fd_sc_hd__mux4_1 c543 (.A0(net526),
    .A1(net532),
    .A2(net524),
    .A3(net533),
    .S0(net530),
    .S1(net518),
    .X(net534));
 sky130_fd_sc_hd__and3_1 c544 (.A(net533),
    .B(net525),
    .C(net529),
    .X(net535));
 sky130_fd_sc_hd__and3_1 c545 (.A(net1035),
    .B(net533),
    .C(net532),
    .X(net536));
 sky130_fd_sc_hd__a2111o_1 c546 (.A1(net533),
    .A2(net532),
    .B1(net885),
    .C1(clknet_1_0__leaf_net914),
    .D1(net1061),
    .X(net537));
 sky130_fd_sc_hd__and3_1 c547 (.A(net531),
    .B(net532),
    .C(net952),
    .X(net538));
 sky130_fd_sc_hd__mux4_1 c548 (.A0(net532),
    .A1(net538),
    .A2(net528),
    .A3(net526),
    .S0(net527),
    .S1(net1061),
    .X(net539));
 sky130_fd_sc_hd__sdfbbp_1 c549 (.CLK(clknet_4_0_0_clk),
    .D(net538),
    .RESET_B(net526),
    .SCD(net884),
    .SCE(clknet_1_0__leaf_net914),
    .SET_B(net1048),
    .Q(net541),
    .Q_N(net540));
 sky130_fd_sc_hd__buf_1 c55 (.A(net981),
    .X(net31));
 sky130_fd_sc_hd__and2_0 c550 (.A(net424),
    .B(net991),
    .X(net542));
 sky130_fd_sc_hd__buf_1 c551 (.A(net542),
    .X(net543));
 sky130_fd_sc_hd__clkbuf_1 c552 (.A(net543),
    .X(net544));
 sky130_fd_sc_hd__clkbuf_1 c553 (.A(net543),
    .X(net545));
 sky130_fd_sc_hd__clkbuf_1 c554 (.A(net972),
    .X(net546));
 sky130_fd_sc_hd__and2_0 c555 (.A(net542),
    .B(net525),
    .X(net547));
 sky130_fd_sc_hd__clkbuf_1 c556 (.A(net525),
    .X(net548));
 sky130_fd_sc_hd__buf_1 c557 (.A(net972),
    .X(net549));
 sky130_fd_sc_hd__and2_0 c558 (.A(net547),
    .B(net549),
    .X(net550));
 sky130_fd_sc_hd__and2_0 c559 (.A(net549),
    .B(net546),
    .X(net551));
 sky130_fd_sc_hd__a2111o_1 c56 (.A1(net31),
    .A2(clknet_1_1__leaf_net29),
    .B1(net30),
    .C1(net1006),
    .D1(clknet_1_1__leaf_net20),
    .X(net32));
 sky130_fd_sc_hd__and2_0 c560 (.A(net551),
    .B(net549),
    .X(net552));
 sky130_fd_sc_hd__and3_1 c561 (.A(net548),
    .B(net552),
    .C(net549),
    .X(net553));
 sky130_fd_sc_hd__and2_0 c562 (.A(net546),
    .B(net548),
    .X(net554));
 sky130_fd_sc_hd__and3_1 c563 (.A(net550),
    .B(net552),
    .C(net404),
    .X(net555));
 sky130_fd_sc_hd__and3_1 c564 (.A(net553),
    .B(net525),
    .X(net873));
 sky130_fd_sc_hd__and3_1 c565 (.A(net545),
    .B(net549),
    .C(net553),
    .X(net557));
 sky130_fd_sc_hd__buf_1 c566 (.A(clknet_1_0__leaf_net994),
    .X(net558));
 sky130_fd_sc_hd__and2_0 c567 (.A(clknet_1_1__leaf_net558),
    .B(net549),
    .X(net559));
 sky130_fd_sc_hd__and3_1 c568 (.A(net553),
    .B(clknet_1_0__leaf_net558),
    .C(net424),
    .X(net560));
 sky130_fd_sc_hd__and2_0 c569 (.A(net559),
    .B(net921),
    .X(net561));
 sky130_fd_sc_hd__buf_6 c57 (.A(net902),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_1 c570 (.A(net921),
    .X(net562));
 sky130_fd_sc_hd__and3_1 c571 (.A(net561),
    .B(net562),
    .C(net873),
    .X(net563));
 sky130_fd_sc_hd__clkbuf_2 c572 (.A(net775),
    .X(net564));
 sky130_fd_sc_hd__and2_0 c573 (.A(net564),
    .B(net970),
    .X(net565));
 sky130_fd_sc_hd__buf_1 c574 (.A(net775),
    .X(net566));
 sky130_fd_sc_hd__clkbuf_1 c575 (.A(net566),
    .X(net567));
 sky130_fd_sc_hd__clkbuf_1 c576 (.A(net919),
    .X(net568));
 sky130_fd_sc_hd__and2_0 c577 (.A(net567),
    .B(net566),
    .X(net569));
 sky130_fd_sc_hd__and2_0 c578 (.A(net568),
    .B(net564),
    .X(net570));
 sky130_fd_sc_hd__buf_1 c579 (.A(net448),
    .X(net571));
 sky130_fd_sc_hd__and3_1 c58 (.A(net33),
    .B(clknet_1_0__leaf_net27),
    .C(clknet_1_1__leaf_net23),
    .X(net34));
 sky130_fd_sc_hd__and3_1 c580 (.A(net564),
    .B(net571),
    .C(net567),
    .X(net572));
 sky130_fd_sc_hd__clkbuf_1 c581 (.A(net978),
    .X(net573));
 sky130_fd_sc_hd__clkbuf_1 c582 (.A(net964),
    .X(net574));
 sky130_fd_sc_hd__and3_1 c583 (.A(net571),
    .B(net570),
    .C(net564),
    .X(net575));
 sky130_fd_sc_hd__and3_1 c584 (.A(net574),
    .B(net566),
    .C(net573),
    .X(net576));
 sky130_fd_sc_hd__and2_0 c585 (.A(net576),
    .B(net571),
    .X(net577));
 sky130_fd_sc_hd__clkbuf_1 c586 (.A(net943),
    .X(net578));
 sky130_fd_sc_hd__and3_1 c587 (.A(net573),
    .B(net578),
    .C(net574),
    .X(net579));
 sky130_fd_sc_hd__and3_1 c588 (.A(net569),
    .B(net570),
    .C(net565),
    .X(net580));
 sky130_fd_sc_hd__and3_1 c589 (.A(net580),
    .B(net576),
    .C(net577),
    .X(net581));
 sky130_fd_sc_hd__sdfbbn_1 c59 (.CLK_N(clknet_4_11_0_clk),
    .D(clknet_1_0__leaf_net26),
    .RESET_B(clknet_1_1__leaf_net34),
    .SCD(net13),
    .SCE(clknet_1_1__leaf_net27),
    .SET_B(clknet_1_1__leaf_net912),
    .Q(net36),
    .Q_N(net35));
 sky130_fd_sc_hd__and3_1 c590 (.A(net1067),
    .B(net580),
    .C(net576),
    .X(net582));
 sky130_fd_sc_hd__a2111o_1 c591 (.A1(net579),
    .A2(net572),
    .B1(net564),
    .C1(net566),
    .D1(net883),
    .X(net583));
 sky130_fd_sc_hd__a2111o_1 c592 (.A1(net580),
    .A2(net576),
    .B1(net564),
    .C1(net883),
    .D1(net975),
    .X(net584));
 sky130_fd_sc_hd__and2_0 c593 (.A(net975),
    .B(net978),
    .X(net585));
 sky130_fd_sc_hd__dlymetal6s2s_1 c594 (.A(net939),
    .X(net586));
 sky130_fd_sc_hd__buf_1 c595 (.A(net586),
    .X(net587));
 sky130_fd_sc_hd__clkbuf_1 c596 (.A(net586),
    .X(net588));
 sky130_fd_sc_hd__and2_1 c597 (.A(net587),
    .B(net586),
    .X(net589));
 sky130_fd_sc_hd__and2_0 c598 (.A(net587),
    .B(net586),
    .X(net590));
 sky130_fd_sc_hd__clkbuf_1 c599 (.A(net908),
    .X(net591));
 sky130_fd_sc_hd__and3_1 c60 (.A(net30),
    .B(clknet_1_1__leaf_net27),
    .C(net35),
    .X(net37));
 sky130_fd_sc_hd__and2_1 c600 (.A(net460),
    .B(net588),
    .X(net592));
 sky130_fd_sc_hd__sdfxtp_1 c601 (.CLK(clknet_4_7_0_clk),
    .D(net592),
    .SCD(net589),
    .SCE(net586),
    .Q(net593));
 sky130_fd_sc_hd__buf_1 c602 (.A(net908),
    .X(net594));
 sky130_fd_sc_hd__and3_1 c603 (.A(net588),
    .B(net589),
    .C(net594),
    .X(net595));
 sky130_fd_sc_hd__and3_1 c604 (.A(net593),
    .B(net594),
    .C(net892),
    .X(net596));
 sky130_fd_sc_hd__and2_0 c605 (.A(net591),
    .B(net593),
    .X(net597));
 sky130_fd_sc_hd__and3_1 c606 (.A(net592),
    .B(net591),
    .C(net594),
    .X(net598));
 sky130_fd_sc_hd__clkbuf_1 c607 (.A(net892),
    .X(net599));
 sky130_fd_sc_hd__and2_0 c608 (.A(net586),
    .B(net599),
    .X(net600));
 sky130_fd_sc_hd__and2_1 c609 (.A(net600),
    .B(net597),
    .X(net601));
 sky130_fd_sc_hd__or4bb_1 c61 (.A(net36),
    .B(clknet_1_1__leaf_net27),
    .C_N(clknet_1_1__leaf_net34),
    .D_N(clknet_1_1__leaf_net912),
    .X(net38));
 sky130_fd_sc_hd__sdfxtp_1 c610 (.CLK(clknet_4_7_0_clk),
    .D(net590),
    .SCD(net594),
    .SCE(net587),
    .Q(net602));
 sky130_fd_sc_hd__and3_1 c611 (.A(net597),
    .B(net591),
    .C(net602),
    .X(net603));
 sky130_fd_sc_hd__mux4_1 c612 (.A0(net603),
    .A1(net588),
    .A2(net594),
    .A3(net602),
    .S0(net592),
    .S1(net1064),
    .X(net604));
 sky130_fd_sc_hd__and3_1 c613 (.A(net596),
    .B(net602),
    .C(net992),
    .X(net605));
 sky130_fd_sc_hd__or4bb_1 c614 (.A(net602),
    .B(net605),
    .C_N(net594),
    .D_N(net1052),
    .X(net606));
 sky130_fd_sc_hd__or4bb_1 c615 (.A(net599),
    .B(net606),
    .C_N(net602),
    .D_N(net1052),
    .X(net607));
 sky130_fd_sc_hd__buf_1 c616 (.A(net978),
    .X(net608));
 sky130_fd_sc_hd__buf_1 c617 (.A(net608),
    .X(net609));
 sky130_fd_sc_hd__buf_1 c618 (.A(net609),
    .X(net610));
 sky130_fd_sc_hd__clkbuf_1 c619 (.A(net905),
    .X(net611));
 sky130_fd_sc_hd__a2111o_1 c62 (.A1(clknet_1_0__leaf_net34),
    .A2(net31),
    .B1(clknet_1_1__leaf_net22),
    .C1(clknet_1_0__leaf_net20),
    .D1(net979),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_1 c620 (.A(net911),
    .X(net612));
 sky130_fd_sc_hd__buf_1 c621 (.A(net911),
    .X(net613));
 sky130_fd_sc_hd__buf_1 c622 (.A(net905),
    .X(net614));
 sky130_fd_sc_hd__and3_1 c623 (.A(net612),
    .B(net613),
    .C(net614),
    .X(net615));
 sky130_fd_sc_hd__and2_0 c624 (.A(net614),
    .B(net977),
    .X(net616));
 sky130_fd_sc_hd__and2_0 c625 (.A(net615),
    .B(net608),
    .X(net617));
 sky130_fd_sc_hd__and2_0 c626 (.A(net609),
    .B(net612),
    .X(net618));
 sky130_fd_sc_hd__and2_0 c627 (.A(net616),
    .B(net614),
    .X(net619));
 sky130_fd_sc_hd__and2_1 c628 (.A(net613),
    .B(net977),
    .X(net1019));
 sky130_fd_sc_hd__buf_1 c629 (.A(net911),
    .X(net620));
 sky130_fd_sc_hd__a2111o_1 c63 (.A1(net36),
    .A2(clknet_1_0__leaf_net34),
    .B1(clknet_1_1__leaf_net23),
    .C1(clknet_1_0__leaf_net912),
    .D1(net927),
    .X(net40));
 sky130_fd_sc_hd__and2_1 c630 (.A(net617),
    .B(net616),
    .X(net621));
 sky130_fd_sc_hd__and2_0 c631 (.A(net615),
    .B(net620),
    .X(net622));
 sky130_fd_sc_hd__and2_1 c632 (.A(net619),
    .B(net620),
    .X(net623));
 sky130_fd_sc_hd__clkbuf_1 c633 (.A(net919),
    .X(net624));
 sky130_fd_sc_hd__or4bb_1 c634 (.A(net611),
    .B(net623),
    .C_N(net617),
    .D_N(net621),
    .X(net625));
 sky130_fd_sc_hd__clkbuf_1 c635 (.A(net941),
    .X(net626));
 sky130_fd_sc_hd__and3_1 c636 (.A(net622),
    .B(net626),
    .C(net868),
    .X(net627));
 sky130_fd_sc_hd__mux4_1 c637 (.A0(net627),
    .A1(net626),
    .A2(net611),
    .A3(net621),
    .S0(net610),
    .X(net868));
 sky130_fd_sc_hd__or4bb_1 c64 (.A(clknet_1_1__leaf_net26),
    .B(net30),
    .C_N(clknet_1_1__leaf_net34),
    .D_N(net927),
    .X(net41));
 sky130_fd_sc_hd__buf_1 c65 (.A(clknet_1_1__leaf_net951),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_2 c651 (.A(net1021),
    .X(net1025));
 sky130_fd_sc_hd__clkbuf_2 c652 (.A(net1057),
    .X(net1022));
 sky130_fd_sc_hd__and3_1 c653 (.A(net1022),
    .B(net517),
    .C(net867),
    .X(net1024));
 sky130_fd_sc_hd__or4bb_1 c654 (.A(net1024),
    .B(net1025),
    .C_N(net510),
    .D_N(net1022),
    .X(net1027));
 sky130_fd_sc_hd__and3_1 c655 (.A(net510),
    .B(net1025),
    .C(net1024),
    .X(net1030));
 sky130_fd_sc_hd__sdfrtp_1 c656 (.CLK(clknet_4_4_0_clk),
    .D(net1030),
    .RESET_B(net1022),
    .SCD(net1024),
    .SCE(net1025),
    .Q(net1023));
 sky130_fd_sc_hd__mux4_1 c657 (.A0(net1023),
    .A1(net1025),
    .A2(net1030),
    .A3(net1024),
    .S0(net1022),
    .S1(net510),
    .X(net629));
 sky130_fd_sc_hd__mux4_1 c658 (.A0(net621),
    .A1(net1022),
    .A2(net1023),
    .A3(net1024),
    .S0(net1025),
    .S1(clknet_1_1__leaf_net1020),
    .X(net630));
 sky130_fd_sc_hd__mux4_1 c659 (.A0(net1025),
    .A1(net1023),
    .A2(net1022),
    .A3(net1024),
    .S0(net1021),
    .S1(clknet_1_0__leaf_net1020),
    .X(net1018));
 sky130_fd_sc_hd__clkbuf_2 c66 (.A(net948),
    .X(net43));
 sky130_fd_sc_hd__buf_1 c660 (.A(net541),
    .X(net631));
 sky130_fd_sc_hd__clkbuf_1 c661 (.A(net631),
    .X(net632));
 sky130_fd_sc_hd__clkbuf_1 c662 (.A(net631),
    .X(net633));
 sky130_fd_sc_hd__and2_1 c663 (.A(net633),
    .B(net631),
    .X(net634));
 sky130_fd_sc_hd__clkbuf_1 c664 (.X(net635));
 sky130_fd_sc_hd__and2_0 c665 (.A(net633),
    .B(net631),
    .X(net636));
 sky130_fd_sc_hd__clkbuf_1 c666 (.A(net769),
    .X(net637));
 sky130_fd_sc_hd__clkbuf_1 c667 (.A(net1069),
    .X(net638));
 sky130_fd_sc_hd__buf_1 c668 (.A(net803),
    .X(net639));
 sky130_fd_sc_hd__and2_1 c669 (.A(net638),
    .B(net639),
    .X(net640));
 sky130_fd_sc_hd__buf_1 c67 (.A(net43),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_1 c670 (.A(net1049),
    .X(net641));
 sky130_fd_sc_hd__and2_0 c671 (.A(net635),
    .B(net633),
    .X(net642));
 sky130_fd_sc_hd__clkbuf_1 c672 (.A(net819),
    .X(net643));
 sky130_fd_sc_hd__and2_0 c673 (.A(net643),
    .B(net641),
    .X(net644));
 sky130_fd_sc_hd__and2_0 c674 (.A(net401),
    .B(net640),
    .X(net645));
 sky130_fd_sc_hd__and2_0 c675 (.A(net640),
    .B(net643),
    .X(net646));
 sky130_fd_sc_hd__or4bb_1 c676 (.A(net645),
    .B(net646),
    .C_N(net640),
    .D_N(net540),
    .X(net647));
 sky130_fd_sc_hd__and2_0 c677 (.A(net641),
    .B(net644),
    .X(net648));
 sky130_fd_sc_hd__and2_0 c678 (.A(net644),
    .B(net646),
    .X(net649));
 sky130_fd_sc_hd__clkbuf_1 c679 (.A(net824),
    .X(net650));
 sky130_fd_sc_hd__and2_1 c68 (.A(net1033),
    .B(net44),
    .X(net45));
 sky130_fd_sc_hd__or4bb_1 c680 (.A(net1050),
    .B(net640),
    .C_N(net645),
    .D_N(net634),
    .X(net651));
 sky130_fd_sc_hd__and2_0 c681 (.A(net650),
    .B(net872),
    .X(net652));
 sky130_fd_sc_hd__buf_1 c682 (.X(net653));
 sky130_fd_sc_hd__buf_1 c683 (.A(net758),
    .X(net654));
 sky130_fd_sc_hd__and2_0 c684 (.A(net639),
    .B(net654),
    .X(net655));
 sky130_fd_sc_hd__and2_0 c685 (.A(net654),
    .B(net653),
    .X(net656));
 sky130_fd_sc_hd__and2_0 c686 (.A(net654),
    .B(net653),
    .X(net657));
 sky130_fd_sc_hd__and2_0 c687 (.A(net653),
    .B(net639),
    .X(net658));
 sky130_fd_sc_hd__and2_1 c688 (.A(net655),
    .B(net639),
    .X(net659));
 sky130_fd_sc_hd__buf_1 c689 (.A(net788),
    .X(net660));
 sky130_fd_sc_hd__clkbuf_1 c69 (.A(net44),
    .X(net46));
 sky130_fd_sc_hd__and2_2 c690 (.A(net658),
    .B(net659),
    .X(net661));
 sky130_fd_sc_hd__and2_0 c691 (.A(net657),
    .B(net653),
    .X(net662));
 sky130_fd_sc_hd__and2_0 c692 (.A(net653),
    .B(net662),
    .X(net663));
 sky130_fd_sc_hd__clkbuf_1 c693 (.A(net964),
    .X(net664));
 sky130_fd_sc_hd__dfbbn_1 c694 (.CLK_N(clknet_4_2_0_clk),
    .D(net656),
    .RESET_B(net660),
    .SET_B(net661),
    .Q(net666),
    .Q_N(net665));
 sky130_fd_sc_hd__and2_0 c695 (.A(net659),
    .B(net654),
    .X(net667));
 sky130_fd_sc_hd__clkbuf_1 c696 (.A(net802),
    .X(net668));
 sky130_fd_sc_hd__and3_1 c697 (.A(net660),
    .B(net668),
    .C(net665),
    .X(net669));
 sky130_fd_sc_hd__and3_1 c698 (.A(net658),
    .B(net656),
    .C(net669),
    .X(net670));
 sky130_fd_sc_hd__and3_1 c699 (.A(net670),
    .B(net669),
    .C(net652),
    .X(net671));
 sky130_fd_sc_hd__and2_1 c70 (.A(net44),
    .B(net43),
    .X(net47));
 sky130_fd_sc_hd__and3_1 c700 (.A(net666),
    .B(net668),
    .C(net671),
    .X(net672));
 sky130_fd_sc_hd__dfbbn_1 c701 (.CLK_N(clknet_4_2_0_clk),
    .D(net671),
    .RESET_B(net670),
    .SET_B(net659),
    .Q(net674),
    .Q_N(net673));
 sky130_fd_sc_hd__or4bb_1 c702 (.A(net667),
    .B(net674),
    .C_N(net660),
    .D_N(net654),
    .X(net675));
 sky130_fd_sc_hd__or4bb_1 c703 (.A(net655),
    .B(net673),
    .C_N(net659),
    .D_N(net924),
    .X(net676));
 sky130_fd_sc_hd__buf_1 c704 (.A(net762),
    .X(net677));
 sky130_fd_sc_hd__clkbuf_1 c705 (.A(net677),
    .X(net678));
 sky130_fd_sc_hd__clkbuf_1 c706 (.A(net762),
    .X(net679));
 sky130_fd_sc_hd__clkbuf_1 c707 (.A(net971),
    .X(net680));
 sky130_fd_sc_hd__clkbuf_1 c708 (.A(net971),
    .X(net681));
 sky130_fd_sc_hd__clkbuf_1 c709 (.A(net680),
    .X(net682));
 sky130_fd_sc_hd__buf_1 c71 (.A(net777),
    .X(net48));
 sky130_fd_sc_hd__buf_2 c710 (.A(net1031),
    .X(net683));
 sky130_fd_sc_hd__and2_2 c711 (.A(net677),
    .B(net683),
    .X(net684));
 sky130_fd_sc_hd__and3_1 c712 (.A(net681),
    .B(net683),
    .C(net684),
    .X(net685));
 sky130_fd_sc_hd__buf_1 c713 (.A(net803),
    .X(net686));
 sky130_fd_sc_hd__and2_0 c714 (.A(net678),
    .B(net684),
    .X(net687));
 sky130_fd_sc_hd__and2_0 c715 (.A(net662),
    .B(net683),
    .X(net688));
 sky130_fd_sc_hd__and2_1 c716 (.A(net682),
    .B(net684),
    .X(net689));
 sky130_fd_sc_hd__and2_0 c717 (.A(net687),
    .B(net686),
    .X(net690));
 sky130_fd_sc_hd__clkbuf_1 c718 (.A(net978),
    .X(net691));
 sky130_fd_sc_hd__clkbuf_1 c719 (.A(net957),
    .X(net692));
 sky130_fd_sc_hd__buf_1 c72 (.A(net901),
    .X(net49));
 sky130_fd_sc_hd__mux4_1 c720 (.A0(net692),
    .A1(net685),
    .A2(net688),
    .A3(net689),
    .S0(net684),
    .S1(net686),
    .X(net693));
 sky130_fd_sc_hd__or4bb_1 c721 (.A(net691),
    .B(net684),
    .C_N(net689),
    .D_N(clknet_1_0__leaf_net993),
    .X(net694));
 sky130_fd_sc_hd__mux4_1 c722 (.A0(net679),
    .A1(clknet_1_1__leaf_net694),
    .A2(net661),
    .A3(net689),
    .S0(net683),
    .S1(clknet_1_1__leaf_net993),
    .X(net695));
 sky130_fd_sc_hd__or4bb_1 c723 (.A(clknet_1_0__leaf_net694),
    .B(net689),
    .C_N(net684),
    .D_N(net968),
    .X(net696));
 sky130_fd_sc_hd__or4bb_1 c724 (.A(net686),
    .B(clknet_1_1__leaf_net694),
    .C_N(net689),
    .D_N(net968),
    .X(net697));
 sky130_fd_sc_hd__or4bb_1 c725 (.A(net689),
    .B(clknet_1_0__leaf_net694),
    .C_N(net669),
    .D_N(clknet_1_1__leaf_net914),
    .X(net698));
 sky130_fd_sc_hd__clkbuf_1 c726 (.A(net767),
    .X(net699));
 sky130_fd_sc_hd__clkbuf_1 c727 (.A(net767),
    .X(net700));
 sky130_fd_sc_hd__buf_1 c728 (.A(net699),
    .X(net701));
 sky130_fd_sc_hd__and2_1 c729 (.A(net700),
    .B(net701),
    .X(net702));
 sky130_fd_sc_hd__clkbuf_1 c73 (.A(net777),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_1 c730 (.A(net701),
    .X(net703));
 sky130_fd_sc_hd__and2_0 c731 (.A(net702),
    .B(net701),
    .X(net704));
 sky130_fd_sc_hd__and2_0 c732 (.A(net683),
    .B(net702),
    .X(net705));
 sky130_fd_sc_hd__and2_1 c733 (.A(net701),
    .B(net700),
    .X(net706));
 sky130_fd_sc_hd__clkbuf_1 c734 (.A(net961),
    .X(net707));
 sky130_fd_sc_hd__clkbuf_1 c735 (.A(net964),
    .X(net708));
 sky130_fd_sc_hd__and3_1 c736 (.A(net702),
    .B(net708),
    .C(net703),
    .X(net709));
 sky130_fd_sc_hd__buf_1 c737 (.A(clknet_1_0__leaf_net949),
    .X(net710));
 sky130_fd_sc_hd__and2_0 c738 (.A(net703),
    .B(net702),
    .X(net711));
 sky130_fd_sc_hd__and2_0 c739 (.A(net706),
    .B(clknet_1_1__leaf_net710),
    .X(net712));
 sky130_fd_sc_hd__and2_0 c74 (.A(net48),
    .B(net49),
    .X(net51));
 sky130_fd_sc_hd__and3_1 c740 (.A(net708),
    .B(net711),
    .C(net705),
    .X(net713));
 sky130_fd_sc_hd__and3_1 c741 (.A(net585),
    .B(net705),
    .C(net706),
    .X(net714));
 sky130_fd_sc_hd__sdfbbn_1 c742 (.CLK_N(clknet_4_0_0_clk),
    .D(clknet_1_0__leaf_net710),
    .RESET_B(net683),
    .SCD(clknet_1_0__leaf_net712),
    .SCE(net953),
    .SET_B(net1038),
    .Q(net716),
    .Q_N(net715));
 sky130_fd_sc_hd__and3_1 c743 (.A(clknet_1_0__leaf_net710),
    .B(net716),
    .C(net969),
    .X(net717));
 sky130_fd_sc_hd__clkbuf_1 c744 (.A(net964),
    .X(net718));
 sky130_fd_sc_hd__or4bb_1 c745 (.A(net707),
    .B(net716),
    .C_N(clknet_1_0__leaf_net717),
    .D_N(net702),
    .X(net719));
 sky130_fd_sc_hd__buf_1 c746 (.A(net983),
    .X(net720));
 sky130_fd_sc_hd__mux4_1 c747 (.A0(clknet_1_0__leaf_net719),
    .A1(clknet_1_0__leaf_net717),
    .A2(net720),
    .A3(net683),
    .S0(net718),
    .S1(clknet_1_1__leaf_net914),
    .X(net721));
 sky130_fd_sc_hd__and2_2 c748 (.A(net614),
    .B(net867),
    .X(net722));
 sky130_fd_sc_hd__and2_0 c749 (.A(net722),
    .B(net614),
    .X(net723));
 sky130_fd_sc_hd__clkbuf_1 c75 (.A(net855),
    .X(net52));
 sky130_fd_sc_hd__and2_0 c750 (.A(net718),
    .B(net722),
    .X(net724));
 sky130_fd_sc_hd__and2_0 c751 (.A(net720),
    .B(net953),
    .X(net725));
 sky130_fd_sc_hd__and2_0 c752 (.A(net725),
    .B(net722),
    .X(net1028));
 sky130_fd_sc_hd__and2_0 c753 (.A(net724),
    .B(net722),
    .X(net726));
 sky130_fd_sc_hd__and2_2 c754 (.A(net720),
    .B(net722),
    .X(net727));
 sky130_fd_sc_hd__and2_1 c755 (.A(net722),
    .B(net727),
    .X(net728));
 sky130_fd_sc_hd__dfbbp_1 c756 (.CLK(clknet_4_1_0_clk),
    .D(net614),
    .RESET_B(net728),
    .SET_B(net727),
    .Q(net730),
    .Q_N(net729));
 sky130_fd_sc_hd__or4bb_1 c757 (.A(net723),
    .B(net727),
    .C_N(net729),
    .D_N(clknet_1_0__leaf_net949),
    .X(net731));
 sky130_fd_sc_hd__clkbuf_1 c758 (.A(net920),
    .X(net732));
 sky130_fd_sc_hd__and2_1 c759 (.A(net730),
    .B(net732),
    .X(net1017));
 sky130_fd_sc_hd__and2_0 c76 (.A(net50),
    .B(net49),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_1 c760 (.A(net920),
    .X(net733));
 sky130_fd_sc_hd__and2_0 c761 (.A(net725),
    .B(net733),
    .X(net734));
 sky130_fd_sc_hd__a2111o_1 c762 (.A1(net726),
    .A2(net728),
    .B1(net723),
    .C1(net1017),
    .D1(net722),
    .X(net735));
 sky130_fd_sc_hd__and3_1 c763 (.A(net733),
    .B(net730),
    .C(net727),
    .X(net736));
 sky130_fd_sc_hd__and3_2 c764 (.A(net734),
    .B(net722),
    .C(net727),
    .X(net737));
 sky130_fd_sc_hd__clkbuf_1 c765 (.A(net911),
    .X(net738));
 sky130_fd_sc_hd__clkbuf_1 c766 (.A(net961),
    .X(net739));
 sky130_fd_sc_hd__sdfbbn_1 c767 (.CLK_N(clknet_4_1_0_clk),
    .D(net732),
    .RESET_B(net736),
    .SCD(net727),
    .SCE(net737),
    .SET_B(net722),
    .Q(net1016),
    .Q_N(net740));
 sky130_fd_sc_hd__mux4_1 c768 (.A0(net728),
    .A1(net739),
    .A2(net1017),
    .A3(net740),
    .S0(net737),
    .S1(net727),
    .X(net741));
 sky130_fd_sc_hd__and3_1 c769 (.A(net727),
    .B(net725),
    .C(net905),
    .X(net1029));
 sky130_fd_sc_hd__buf_1 c77 (.A(net976),
    .X(net54));
 sky130_fd_sc_hd__buf_1 c78 (.A(net900),
    .X(net55));
 sky130_fd_sc_hd__and3_1 c79 (.A(net51),
    .B(net53),
    .C(net55),
    .X(net56));
 sky130_fd_sc_hd__and3_2 c80 (.A(net56),
    .B(net44),
    .C(net53),
    .X(net57));
 sky130_fd_sc_hd__and3_1 c81 (.A(net37),
    .B(net56),
    .C(net54),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_1 c82 (.A(net941),
    .X(net59));
 sky130_fd_sc_hd__and3_1 c83 (.A(net52),
    .B(net54),
    .C(net55),
    .X(net60));
 sky130_fd_sc_hd__and3_1 c84 (.A(net59),
    .B(net55),
    .C(net60),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_1 c85 (.A(net941),
    .X(net62));
 sky130_fd_sc_hd__or4bb_1 c86 (.A(net53),
    .B(net60),
    .C_N(net55),
    .D_N(net57),
    .X(net63));
 sky130_fd_sc_hd__a2111o_1 c87 (.A1(net62),
    .A2(net60),
    .B1(net57),
    .C1(net55),
    .X(net64));
 sky130_fd_sc_hd__buf_1 c88 (.A(net43),
    .X(net65));
 sky130_fd_sc_hd__buf_1 c89 (.A(net65),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_2 c90 (.A(net65),
    .X(net67));
 sky130_fd_sc_hd__buf_1 c91 (.A(net931),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_1 c92 (.A(net931),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_1 c93 (.A(net982),
    .X(net70));
 sky130_fd_sc_hd__and2_1 c94 (.A(net69),
    .B(net68),
    .X(net71));
 sky130_fd_sc_hd__and2_0 c95 (.A(net71),
    .B(net68),
    .X(net72));
 sky130_fd_sc_hd__buf_1 c96 (.A(net808),
    .X(net73));
 sky130_fd_sc_hd__clkbuf_1 c97 (.A(net982),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_1 c98 (.A(net928),
    .X(net75));
 sky130_fd_sc_hd__and2_1 c99 (.A(net75),
    .B(net71),
    .X(net76));
 sky130_fd_sc_hd__mux4_1 merge782 (.A0(net7),
    .A1(net995),
    .A2(net3),
    .A3(net11),
    .S0(net12),
    .S1(net13),
    .X(net742));
 sky130_fd_sc_hd__and3_1 merge783 (.A(clknet_1_1__leaf_net226),
    .B(clknet_1_1__leaf_net325),
    .C(net339),
    .X(net743));
 sky130_fd_sc_hd__or4bb_1 merge784 (.A(net252),
    .B(net251),
    .C_N(net256),
    .D_N(net253),
    .X(net744));
 sky130_fd_sc_hd__or4bb_1 merge785 (.A(net118),
    .B(net117),
    .C_N(net122),
    .D_N(net997),
    .X(net745));
 sky130_fd_sc_hd__or4bb_1 merge786 (.A(clknet_1_0__leaf_net89),
    .B(net94),
    .C_N(net93),
    .D_N(clknet_1_0__leaf_net95),
    .X(net746));
 sky130_fd_sc_hd__buf_1 merge787 (.A(clknet_1_0__leaf_net950),
    .X(net747));
 sky130_fd_sc_hd__and3_1 merge788 (.A(net430),
    .B(net431),
    .C(net432),
    .X(net748));
 sky130_fd_sc_hd__or4bb_1 merge789 (.A(net731),
    .B(net729),
    .C_N(net1017),
    .D_N(net726),
    .X(net749));
 sky130_fd_sc_hd__and3_1 merge790 (.A(net609),
    .B(net610),
    .C(net608),
    .X(net750));
 sky130_fd_sc_hd__clkbuf_1 merge791 (.A(net940),
    .X(net751));
 sky130_fd_sc_hd__sdfxbp_1 merge792 (.CLK(clknet_4_0_0_clk),
    .D(net405),
    .SCD(net522),
    .SCE(net519),
    .Q(net753),
    .Q_N(net752));
 sky130_fd_sc_hd__and3_1 merge793 (.A(net139),
    .B(net140),
    .C(net142),
    .X(net754));
 sky130_fd_sc_hd__or4bb_1 merge794 (.A(clknet_1_1__leaf_net160),
    .B(clknet_1_0__leaf_net161),
    .C_N(clknet_1_1__leaf_net162),
    .D_N(net13),
    .X(net755));
 sky130_fd_sc_hd__clkbuf_1 merge795 (.A(net781),
    .X(net756));
 sky130_fd_sc_hd__or4bb_1 merge796 (.A(clknet_1_0__leaf_net162),
    .B(net181),
    .C_N(net297),
    .D_N(net956),
    .X(net757));
 sky130_fd_sc_hd__sdfxbp_1 merge797 (.CLK(clknet_4_2_0_clk),
    .D(net652),
    .SCD(clknet_1_1__leaf_net563),
    .Q(net653),
    .Q_N(net758));
 sky130_fd_sc_hd__clkbuf_1 merge798 (.A(net955),
    .X(net760));
 sky130_fd_sc_hd__clkbuf_1 merge799 (.A(net929),
    .X(net761));
 sky130_fd_sc_hd__clkbuf_1 merge800 (.A(net940),
    .X(net762));
 sky130_fd_sc_hd__and3_1 merge801 (.A(net544),
    .B(net543),
    .C(net991),
    .X(net763));
 sky130_fd_sc_hd__buf_1 merge802 (.A(clknet_1_1__leaf_net950),
    .X(net764));
 sky130_fd_sc_hd__and3_1 merge803 (.A(net182),
    .B(net184),
    .C(net57),
    .X(net765));
 sky130_fd_sc_hd__or4bb_1 merge804 (.A(net65),
    .B(net67),
    .C_N(net66),
    .D_N(net68),
    .X(net766));
 sky130_fd_sc_hd__clkbuf_1 merge805 (.A(net958),
    .X(net767));
 sky130_fd_sc_hd__or4bb_1 merge806 (.A(clknet_1_0__leaf_net226),
    .B(net230),
    .C_N(net231),
    .D_N(net959),
    .X(net768));
 sky130_fd_sc_hd__sdfxtp_1 merge807 (.CLK(clknet_4_0_0_clk),
    .D(net634),
    .SCD(net525),
    .Q(net635));
 sky130_fd_sc_hd__and3_1 merge808 (.A(net19),
    .B(net1006),
    .C(net13),
    .X(net770));
 sky130_fd_sc_hd__clkbuf_1 merge809 (.A(net980),
    .X(net771));
 sky130_fd_sc_hd__or4bb_1 merge810 (.A(net590),
    .B(net460),
    .C_N(net593),
    .D_N(net575),
    .X(net772));
 sky130_fd_sc_hd__buf_1 merge811 (.A(net932),
    .X(net773));
 sky130_fd_sc_hd__and3_1 merge812 (.A(clknet_1_1__leaf_net272),
    .B(net264),
    .C(net273),
    .X(net774));
 sky130_fd_sc_hd__clkbuf_1 merge813 (.A(net940),
    .X(net775));
 sky130_fd_sc_hd__mux4_1 merge814 (.A0(net589),
    .A1(net1019),
    .A2(net381),
    .A3(net517),
    .S0(net621),
    .S1(net1025),
    .X(net776));
 sky130_fd_sc_hd__clkbuf_1 merge815 (.A(net944),
    .X(net777));
 sky130_fd_sc_hd__sdfrtp_1 merge816 (.CLK(clknet_4_14_0_clk),
    .D(net359),
    .RESET_B(net358),
    .SCD(clknet_1_0__leaf_net213),
    .SCE(clknet_1_1__leaf_net207),
    .Q(net778));
 sky130_fd_sc_hd__or4bb_1 merge817 (.A(net601),
    .B(net433),
    .C_N(net439),
    .D_N(clknet_1_1__leaf_net949),
    .X(net779));
 sky130_fd_sc_hd__or4bb_1 merge818 (.A(net119),
    .B(net123),
    .C_N(net140),
    .D_N(net142),
    .X(net780));
 sky130_fd_sc_hd__clkbuf_1 merge819 (.A(net871),
    .X(net781));
 sky130_fd_sc_hd__or4bb_1 merge820 (.A(net176),
    .B(clknet_1_0__leaf_net168),
    .C_N(net169),
    .D_N(net165),
    .X(net782));
 sky130_fd_sc_hd__or4bb_1 merge821 (.A(net389),
    .B(net386),
    .C_N(net434),
    .D_N(net432),
    .X(net783));
 sky130_fd_sc_hd__or4bb_1 merge822 (.A(net300),
    .B(net302),
    .C_N(net138),
    .D_N(net142),
    .X(net784));
 sky130_fd_sc_hd__or4bb_1 merge823 (.A(clknet_1_1__leaf_net317),
    .B(clknet_1_0__leaf_net325),
    .C_N(net45),
    .D_N(net47),
    .X(net785));
 sky130_fd_sc_hd__or4bb_1 merge824 (.A(net296),
    .B(net302),
    .C_N(net336),
    .D_N(net327),
    .X(net786));
 sky130_fd_sc_hd__sdfsbp_1 merge825 (.CLK(clknet_4_0_0_clk),
    .D(net659),
    .SCD(clknet_1_0__leaf_net563),
    .SCE(net522),
    .SET_B(net526),
    .Q(net788),
    .Q_N(net787));
 sky130_fd_sc_hd__or4bb_1 merge826 (.A(net190),
    .B(net193),
    .C_N(net165),
    .D_N(clknet_1_0__leaf_net168),
    .X(net789));
 sky130_fd_sc_hd__or4bb_1 merge827 (.A(net349),
    .B(net484),
    .C_N(net346),
    .D_N(net345),
    .X(net790));
 sky130_fd_sc_hd__or4bb_1 merge828 (.A(net453),
    .B(net456),
    .C_N(net435),
    .D_N(net434),
    .X(net791));
 sky130_fd_sc_hd__sdfsbp_1 merge829 (.CLK(clknet_4_5_0_clk),
    .D(net524),
    .SCD(net523),
    .SCE(net261),
    .SET_B(net252),
    .Q(net793),
    .Q_N(net792));
 sky130_fd_sc_hd__or4bb_1 merge830 (.A(net690),
    .B(net683),
    .C_N(net565),
    .D_N(net572),
    .X(net794));
 sky130_fd_sc_hd__or4bb_1 merge831 (.A(net189),
    .B(net184),
    .C_N(net461),
    .D_N(net455),
    .X(net795));
 sky130_fd_sc_hd__or4bb_1 merge832 (.A(net301),
    .B(net300),
    .C_N(net451),
    .D_N(net453),
    .X(net796));
 sky130_fd_sc_hd__or4bb_1 merge833 (.A(net322),
    .B(clknet_1_1__leaf_net321),
    .C_N(clknet_1_0__leaf_net29),
    .D_N(clknet_1_0__leaf_net24),
    .X(net797));
 sky130_fd_sc_hd__or4bb_1 merge834 (.A(net260),
    .B(net259),
    .C_N(net281),
    .D_N(net284),
    .X(net798));
 sky130_fd_sc_hd__or4bb_1 merge835 (.A(clknet_1_0__leaf_net272),
    .B(net276),
    .C_N(net577),
    .D_N(net576),
    .X(net799));
 sky130_fd_sc_hd__or4bb_1 merge836 (.A(net566),
    .B(clknet_1_0__leaf_net563),
    .C_N(net610),
    .D_N(net1019),
    .X(net800));
 sky130_fd_sc_hd__or4bb_1 merge837 (.A(net705),
    .B(net701),
    .C_N(net737),
    .D_N(net738),
    .X(net801));
 sky130_fd_sc_hd__sdfstp_1 merge838 (.CLK(clknet_4_2_0_clk),
    .D(net664),
    .SCD(net661),
    .SCE(net632),
    .SET_B(net634),
    .Q(net802));
 sky130_fd_sc_hd__sdfstp_1 merge839 (.CLK(clknet_4_2_0_clk),
    .D(net636),
    .SCD(net634),
    .SCE(net661),
    .SET_B(net684),
    .Q(net803));
 sky130_fd_sc_hd__or4bb_1 merge840 (.A(net306),
    .B(net302),
    .C_N(net274),
    .D_N(clknet_1_1__leaf_net272),
    .X(net804));
 sky130_fd_sc_hd__or4bb_1 merge841 (.A(net362),
    .B(net365),
    .C_N(clknet_1_0__leaf_net321),
    .D_N(clknet_1_1__leaf_net324),
    .X(net805));
 sky130_fd_sc_hd__or4bb_1 merge842 (.A(net483),
    .B(clknet_1_1__leaf_net482),
    .C_N(net476),
    .D_N(net478),
    .X(net806));
 sky130_fd_sc_hd__sdfstp_1 merge843 (.CLK(clknet_4_2_0_clk),
    .D(net637),
    .SCD(net634),
    .SCE(net421),
    .SET_B(net422),
    .Q(net807));
 sky130_fd_sc_hd__sedfxbp_1 merge844 (.CLK(clknet_4_11_0_clk),
    .D(net211),
    .DE(net66),
    .SCD(net71),
    .SCE(net1066),
    .Q(net809),
    .Q_N(net808));
 sky130_fd_sc_hd__or4bb_1 merge845 (.A(net572),
    .B(net569),
    .C_N(net704),
    .D_N(net706),
    .X(net810));
 sky130_fd_sc_hd__or4bb_1 merge846 (.A(net65),
    .B(net57),
    .C_N(net68),
    .D_N(net67),
    .X(net811));
 sky130_fd_sc_hd__or4bb_1 merge847 (.A(clknet_1_1__leaf_net197),
    .B(clknet_1_0__leaf_net201),
    .C_N(clknet_1_0__leaf_net162),
    .D_N(net187),
    .X(net812));
 sky130_fd_sc_hd__or4bb_1 merge848 (.A(net165),
    .B(clknet_1_0__leaf_net160),
    .C_N(net45),
    .D_N(net48),
    .X(net813));
 sky130_fd_sc_hd__a2111o_1 merge849 (.A1(net608),
    .A2(net610),
    .B1(net609),
    .C1(net613),
    .D1(net943),
    .X(net814));
 sky130_fd_sc_hd__or4bb_1 merge850 (.A(net486),
    .B(net478),
    .C_N(net459),
    .D_N(net965),
    .X(net815));
 sky130_fd_sc_hd__or4bb_1 merge851 (.A(net67),
    .B(net68),
    .C_N(clknet_1_1__leaf_net91),
    .D_N(net231),
    .X(net816));
 sky130_fd_sc_hd__or4bb_1 merge852 (.A(net392),
    .B(net386),
    .C_N(clknet_1_1__leaf_net563),
    .D_N(net924),
    .X(net817));
 sky130_fd_sc_hd__sedfxbp_1 merge853 (.CLK(clknet_4_2_0_clk),
    .D(net642),
    .DE(net639),
    .SCD(net424),
    .SCE(net434),
    .Q(net819),
    .Q_N(net818));
 sky130_fd_sc_hd__or4bb_1 merge854 (.A(net389),
    .B(net392),
    .C_N(clknet_1_0__leaf_net25),
    .D_N(clknet_1_0__leaf_net912),
    .X(net820));
 sky130_fd_sc_hd__or4bb_1 merge855 (.A(net406),
    .B(net414),
    .C_N(clknet_1_0__leaf_net330),
    .D_N(clknet_1_0__leaf_net329),
    .X(net821));
 sky130_fd_sc_hd__mux4_1 merge856 (.A0(net618),
    .A1(net613),
    .A2(net617),
    .A3(net728),
    .S0(net737),
    .S1(net905),
    .X(net822));
 sky130_fd_sc_hd__or4bb_1 merge857 (.A(clknet_1_0__leaf_net321),
    .B(clknet_1_0__leaf_net317),
    .C_N(net415),
    .D_N(net420),
    .X(net823));
 sky130_fd_sc_hd__sedfxtp_1 merge858 (.CLK(clknet_4_2_0_clk),
    .D(net649),
    .DE(net419),
    .SCD(net414),
    .SCE(net872),
    .Q(net824));
 sky130_fd_sc_hd__or4bb_1 merge859 (.A(clknet_1_0__leaf_net21),
    .B(clknet_1_1__leaf_net25),
    .C_N(net408),
    .D_N(net414),
    .X(net825));
 sky130_fd_sc_hd__or4bb_1 merge860 (.A(net219),
    .B(net345),
    .C_N(net13),
    .D_N(clknet_1_1__leaf_net20),
    .X(net826));
 sky130_fd_sc_hd__sedfxtp_1 merge861 (.CLK(clknet_4_9_0_clk),
    .D(net369),
    .DE(net362),
    .SCD(net343),
    .SCE(net345),
    .Q(net827));
 sky130_fd_sc_hd__a2111o_1 merge862 (.A1(net228),
    .A2(net365),
    .B1(net70),
    .C1(clknet_1_0__leaf_net81),
    .D1(net963),
    .X(net828));
 sky130_fd_sc_hd__and3_1 merge863 (.A(net669),
    .B(net575),
    .C(net676),
    .X(net829));
 sky130_fd_sc_hd__a2111o_1 merge864 (.A1(net394),
    .A2(net389),
    .B1(net392),
    .C1(net393),
    .D1(net397),
    .X(net830));
 sky130_fd_sc_hd__mux4_1 merge865 (.A0(net125),
    .A1(net123),
    .A2(net122),
    .A3(net140),
    .S0(net142),
    .S1(net870),
    .X(net831));
 sky130_fd_sc_hd__mux4_1 merge866 (.A0(clknet_1_0__leaf_net357),
    .A1(clknet_1_1__leaf_net353),
    .A2(net347),
    .A3(net188),
    .S0(net187),
    .S1(net183),
    .X(net832));
 sky130_fd_sc_hd__mux4_1 merge867 (.A0(net47),
    .A1(net43),
    .A2(net46),
    .A3(net49),
    .S0(net54),
    .S1(net979),
    .X(net833));
 sky130_fd_sc_hd__mux4_1 merge868 (.A0(clknet_1_1__leaf_net329),
    .A1(clknet_1_0__leaf_net324),
    .A2(net322),
    .A3(net488),
    .S0(net481),
    .S1(net478),
    .X(net834));
 sky130_fd_sc_hd__mux4_1 merge869 (.A0(clknet_1_1__leaf_net42),
    .A1(net47),
    .A2(net45),
    .A3(net509),
    .S0(net922),
    .S1(net958),
    .X(net835));
 sky130_fd_sc_hd__mux4_1 merge870 (.A0(net311),
    .A1(net305),
    .A2(net307),
    .A3(net249),
    .S0(net362),
    .S1(net365),
    .X(net836));
 sky130_fd_sc_hd__mux4_1 merge871 (.A0(net366),
    .A1(net365),
    .A2(clknet_1_1__leaf_net712),
    .A3(clknet_1_1__leaf_net717),
    .S0(clknet_1_1__leaf_net719),
    .S1(net945),
    .X(net837));
 sky130_fd_sc_hd__mux4_1 merge872 (.A0(net67),
    .A1(clknet_1_1__leaf_net210),
    .A2(clknet_1_1__leaf_net213),
    .A3(net130),
    .S0(net118),
    .S1(net124),
    .X(net838));
 sky130_fd_sc_hd__a2111o_1 merge873 (.A1(net395),
    .A2(net399),
    .B1(net397),
    .C1(net398),
    .D1(net390),
    .X(net839));
 sky130_fd_sc_hd__mux4_1 merge874 (.A0(net151),
    .A1(net152),
    .A2(net142),
    .A3(net124),
    .S0(net131),
    .S1(net130),
    .X(net840));
 sky130_fd_sc_hd__mux4_1 merge875 (.A0(net554),
    .A1(net553),
    .A2(net252),
    .A3(net258),
    .S0(net254),
    .S1(net1037),
    .X(net841));
 sky130_fd_sc_hd__mux4_1 merge876 (.A0(net709),
    .A1(net708),
    .A2(net706),
    .A3(net439),
    .S0(net436),
    .S1(net970),
    .X(net842));
 sky130_fd_sc_hd__a2111o_1 merge877 (.A1(net259),
    .A2(net257),
    .B1(net260),
    .C1(net263),
    .D1(net264),
    .X(net843));
 sky130_fd_sc_hd__mux4_1 merge878 (.A0(net663),
    .A1(net660),
    .A2(net661),
    .A3(clknet_1_1__leaf_net717),
    .S0(net715),
    .S1(net709),
    .X(net844));
 sky130_fd_sc_hd__mux4_1 merge879 (.A0(net428),
    .A1(clknet_1_1__leaf_net563),
    .A2(net564),
    .A3(net378),
    .S0(net248),
    .S1(net931),
    .X(net845));
 sky130_fd_sc_hd__mux4_1 merge880 (.A0(net688),
    .A1(net689),
    .A2(net683),
    .A3(net1012),
    .S0(clknet_1_0__leaf_net145),
    .S1(net140),
    .X(net846));
 sky130_fd_sc_hd__mux4_1 merge881 (.A0(net368),
    .A1(net366),
    .A2(net362),
    .A3(clknet_1_1__leaf_net81),
    .S0(net84),
    .S1(clknet_1_0__leaf_net85),
    .X(net847));
 sky130_fd_sc_hd__mux4_1 merge882 (.A0(net367),
    .A1(net509),
    .A2(net300),
    .A3(net303),
    .S0(net308),
    .S1(net965),
    .X(net848));
 sky130_fd_sc_hd__mux4_1 merge883 (.A0(net410),
    .A1(net411),
    .A2(net409),
    .A3(net132),
    .S0(clknet_1_0__leaf_net127),
    .S1(net130),
    .X(net849));
 sky130_fd_sc_hd__mux4_1 merge884 (.A0(net307),
    .A1(net302),
    .A2(net477),
    .A3(net476),
    .S0(net478),
    .S1(net990),
    .X(net850));
 sky130_fd_sc_hd__mux4_1 merge885 (.A0(net624),
    .A1(net623),
    .A2(net620),
    .A3(net283),
    .S0(net278),
    .S1(net1058),
    .X(net851));
 sky130_fd_sc_hd__mux4_1 merge886 (.A0(net676),
    .A1(net575),
    .A2(net677),
    .A3(clknet_1_0__leaf_net498),
    .S0(clknet_1_0__leaf_net496),
    .S1(net481),
    .X(net852));
 sky130_fd_sc_hd__a2111o_1 merge887 (.A1(net49),
    .A2(net57),
    .B1(net52),
    .C1(net61),
    .D1(net58),
    .X(net853));
 sky130_fd_sc_hd__and2_0 merge888 (.A(net696),
    .B(net697),
    .X(net854));
 sky130_fd_sc_hd__dfrbp_1 merge889 (.CLK(clknet_4_12_0_clk),
    .D(net338),
    .RESET_B(net785),
    .Q(net856),
    .Q_N(net855));
 sky130_fd_sc_hd__and2_0 merge890 (.A(net714),
    .B(net721),
    .X(net857));
 sky130_fd_sc_hd__and2_0 merge891 (.A(net38),
    .B(net40),
    .X(net858));
 sky130_fd_sc_hd__and2_0 merge892 (.A(net462),
    .B(net464),
    .X(net859));
 sky130_fd_sc_hd__and2_0 merge893 (.A(net154),
    .B(net157),
    .X(net860));
 sky130_fd_sc_hd__and2_0 merge894 (.A(net78),
    .B(net83),
    .X(net861));
 sky130_fd_sc_hd__and2_0 merge895 (.A(net672),
    .B(net675),
    .X(net862));
 sky130_fd_sc_hd__and2_0 merge896 (.A(net173),
    .B(net174),
    .X(net863));
 sky130_fd_sc_hd__and2_0 merge897 (.A(net288),
    .B(net289),
    .X(net864));
 sky130_fd_sc_hd__and2_1 merge898 (.A(net417),
    .B(net426),
    .X(net865));
 sky130_fd_sc_hd__and2_0 merge899 (.A(net348),
    .B(net351),
    .X(net866));
 sky130_fd_sc_hd__dfrbp_1 merge900 (.CLK(clknet_4_4_0_clk),
    .D(net625),
    .Q(net868),
    .Q_N(net867));
 sky130_fd_sc_hd__and2_0 merge901 (.A(net111),
    .B(net115),
    .X(net869));
 sky130_fd_sc_hd__dfrtn_1 merge902 (.CLK_N(clknet_4_7_0_clk),
    .D(net128),
    .RESET_B(net137),
    .Q(net870));
 sky130_fd_sc_hd__dfrtp_1 merge903 (.CLK(clknet_4_8_0_clk),
    .D(net403),
    .RESET_B(net783),
    .Q(net871));
 sky130_fd_sc_hd__dfrtp_1 merge904 (.CLK(clknet_4_2_0_clk),
    .D(net647),
    .RESET_B(net651),
    .Q(net872));
 sky130_fd_sc_hd__dfrtp_1 merge905 (.CLK(clknet_4_4_0_clk),
    .RESET_B(net1060),
    .Q(net873));
 sky130_fd_sc_hd__and2_0 merge906 (.A(net14),
    .B(net17),
    .X(net874));
 sky130_fd_sc_hd__dfsbp_1 merge907 (.CLK(clknet_4_13_0_clk),
    .D(net310),
    .SET_B(net757),
    .Q(net876),
    .Q_N(net875));
 sky130_fd_sc_hd__and2_0 merge908 (.A(net196),
    .B(net198),
    .X(net877));
 sky130_fd_sc_hd__dfsbp_1 merge909 (.CLK(clknet_4_14_0_clk),
    .D(net212),
    .SET_B(net223),
    .Q(net879),
    .Q_N(net878));
 sky130_fd_sc_hd__and2_0 merge910 (.A(net735),
    .B(net741),
    .X(net880));
 sky130_fd_sc_hd__dfstp_1 merge911 (.CLK(clknet_4_5_0_clk),
    .D(net776),
    .SET_B(net630),
    .Q(net1021));
 sky130_fd_sc_hd__and2_0 merge912 (.A(net505),
    .B(net511),
    .X(net881));
 sky130_fd_sc_hd__dfstp_1 merge913 (.CLK(clknet_4_15_0_clk),
    .D(net63),
    .Q(net64));
 sky130_fd_sc_hd__dfstp_1 merge914 (.CLK(clknet_4_4_0_clk),
    .D(net581),
    .SET_B(net582),
    .Q(net883));
 sky130_fd_sc_hd__dlrbn_1 merge915 (.D(net534),
    .GATE_N(clknet_4_0_0_clk),
    .RESET_B(net1062),
    .Q(net885),
    .Q_N(net884));
 sky130_fd_sc_hd__and2_0 merge916 (.A(net485),
    .B(net492),
    .X(net886));
 sky130_fd_sc_hd__and2_0 merge917 (.A(net372),
    .B(net379),
    .X(net887));
 sky130_fd_sc_hd__dlrbn_1 merge918 (.D(net245),
    .GATE_N(clknet_4_10_0_clk),
    .RESET_B(net238),
    .Q(net889),
    .Q_N(net888));
 sky130_fd_sc_hd__and2_0 merge919 (.A(net268),
    .B(net270),
    .X(net890));
 sky130_fd_sc_hd__dlrbp_1 merge920 (.D(net595),
    .GATE(clknet_4_7_0_clk),
    .RESET_B(net598),
    .Q(net892),
    .Q_N(net891));
 sky130_fd_sc_hd__and2_0 merge921 (.A(net438),
    .B(net450),
    .X(net893));
 sky130_fd_sc_hd__and2_0 merge922 (.A(net863),
    .B(net18),
    .X(net894));
 sky130_fd_sc_hd__and2_0 merge923 (.A(net584),
    .B(net495),
    .X(net895));
 sky130_fd_sc_hd__and2_0 merge924 (.A(net469),
    .B(net472),
    .X(net896));
 sky130_fd_sc_hd__and2_0 merge925 (.A(net202),
    .B(net204),
    .X(net897));
 sky130_fd_sc_hd__and2_0 merge926 (.A(net494),
    .B(net224),
    .X(net898));
 sky130_fd_sc_hd__and2_1 merge927 (.A(net291),
    .B(net271),
    .X(net899));
 sky130_fd_sc_hd__dlrbp_1 merge928 (.D(net225),
    .GATE(clknet_4_14_0_clk),
    .RESET_B(net833),
    .Q(net901),
    .Q_N(net900));
 sky130_fd_sc_hd__dlrtn_2 merge929 (.D(net817),
    .GATE_N(clknet_4_8_0_clk),
    .RESET_B(net820),
    .Q(net902));
 sky130_fd_sc_hd__and2_0 merge930 (.A(net355),
    .B(net383),
    .X(net903));
 sky130_fd_sc_hd__dlrtn_1 merge931 (.D(net172),
    .GATE_N(clknet_4_13_0_clk),
    .RESET_B(net755),
    .Q(net904));
 sky130_fd_sc_hd__dlrtn_1 merge932 (.D(net814),
    .GATE_N(clknet_4_1_0_clk),
    .RESET_B(net880),
    .Q(net905));
 sky130_fd_sc_hd__dlrtp_1 merge933 (.D(net292),
    .GATE(clknet_4_5_0_clk),
    .RESET_B(net744),
    .Q(net906));
 sky130_fd_sc_hd__dlrtp_1 merge934 (.D(net860),
    .GATE(clknet_4_13_0_clk),
    .RESET_B(net745),
    .Q(net907));
 sky130_fd_sc_hd__dlrtp_1 merge935 (.D(net823),
    .GATE(clknet_4_7_0_clk),
    .RESET_B(net772),
    .Q(net908));
 sky130_fd_sc_hd__edfxbp_1 merge936 (.CLK(clknet_4_10_0_clk),
    .D(net746),
    .DE(net768),
    .Q(net910),
    .Q_N(net909));
 sky130_fd_sc_hd__edfxtp_1 merge937 (.CLK(clknet_4_1_0_clk),
    .D(net750),
    .DE(net822),
    .Q(net911));
 sky130_fd_sc_hd__sdlclkp_1 merge938 (.CLK(clknet_4_9_0_clk),
    .GATE(net28),
    .SCE(net32),
    .GCLK(net912));
 sky130_fd_sc_hd__and2_0 merge939 (.A(net512),
    .B(net513),
    .X(net913));
 sky130_fd_sc_hd__sdlclkp_2 merge940 (.CLK(clknet_4_0_0_clk),
    .GATE(net854),
    .SCE(net535),
    .GCLK(net914));
 sky130_fd_sc_hd__sdlclkp_4 merge941 (.CLK(clknet_4_7_0_clk),
    .GATE(net780),
    .SCE(net831),
    .GCLK(net915));
 sky130_fd_sc_hd__dfrbp_1 merge942 (.CLK(clknet_4_12_0_clk),
    .D(net815),
    .RESET_B(net784),
    .Q(net917),
    .Q_N(net916));
 sky130_fd_sc_hd__and2_0 merge943 (.A(net514),
    .B(net913),
    .X(net918));
 sky130_fd_sc_hd__dfrbp_1 merge944 (.CLK(clknet_4_1_0_clk),
    .D(net749),
    .RESET_B(net800),
    .Q(net920),
    .Q_N(net919));
 sky130_fd_sc_hd__dfrtn_1 merge945 (.CLK_N(clknet_4_4_0_clk),
    .D(net557),
    .RESET_B(net560),
    .Q(net921));
 sky130_fd_sc_hd__dfrtp_2 merge946 (.CLK(clknet_4_6_0_clk),
    .D(net515),
    .RESET_B(net791),
    .Q(net922));
 sky130_fd_sc_hd__dfrtp_1 merge947 (.CLK(clknet_4_9_0_clk),
    .D(net797),
    .RESET_B(net834),
    .Q(net923));
 sky130_fd_sc_hd__dfrtp_2 merge948 (.CLK(clknet_4_0_0_clk),
    .D(net862),
    .RESET_B(net1036),
    .Q(net924));
 sky130_fd_sc_hd__dfsbp_1 merge949 (.CLK(clknet_4_5_0_clk),
    .D(net798),
    .SET_B(net1047),
    .Q(net926),
    .Q_N(net925));
 sky130_fd_sc_hd__dfsbp_1 merge950 (.CLK(clknet_4_9_0_clk),
    .D(net816),
    .SET_B(net39),
    .Q(net928),
    .Q_N(net927));
 sky130_fd_sc_hd__dfstp_2 merge951 (.CLK(clknet_4_14_0_clk),
    .D(net836),
    .SET_B(net1043),
    .Q(net929));
 sky130_fd_sc_hd__dfstp_1 merge952 (.CLK(clknet_4_14_0_clk),
    .D(net765),
    .SET_B(net742),
    .Q(net930));
 sky130_fd_sc_hd__dfstp_1 merge953 (.CLK(clknet_4_9_0_clk),
    .D(net887),
    .SET_B(net766),
    .Q(net931));
 sky130_fd_sc_hd__dlrbn_1 merge954 (.D(net774),
    .GATE_N(clknet_4_6_0_clk),
    .RESET_B(net849),
    .Q(net933),
    .Q_N(net932));
 sky130_fd_sc_hd__dlrbn_1 merge955 (.D(net821),
    .GATE_N(clknet_4_9_0_clk),
    .RESET_B(net748),
    .Q(net935),
    .Q_N(net934));
 sky130_fd_sc_hd__dlrbp_1 merge956 (.D(net830),
    .GATE(clknet_4_8_0_clk),
    .RESET_B(net839),
    .Q(net937),
    .Q_N(net936));
 sky130_fd_sc_hd__dlrbp_1 merge957 (.D(net896),
    .GATE(clknet_4_7_0_clk),
    .RESET_B(net155),
    .Q(net939),
    .Q_N(net938));
 sky130_fd_sc_hd__dlrtn_1 merge958 (.D(net845),
    .GATE_N(clknet_4_3_0_clk),
    .RESET_B(net852),
    .Q(net940));
 sky130_fd_sc_hd__dlrtn_2 merge959 (.D(net853),
    .GATE_N(clknet_4_6_0_clk),
    .RESET_B(net851),
    .Q(net941));
 sky130_fd_sc_hd__dlrtn_2 merge960 (.D(net789),
    .GATE_N(clknet_4_15_0_clk),
    .RESET_B(net898),
    .Q(net942));
 sky130_fd_sc_hd__dlrtp_1 merge961 (.D(net886),
    .GATE(clknet_4_4_0_clk),
    .RESET_B(net799),
    .Q(net943));
 sky130_fd_sc_hd__dlrtp_1 merge962 (.D(net835),
    .GATE(clknet_4_12_0_clk),
    .RESET_B(net795),
    .Q(net944));
 sky130_fd_sc_hd__dlrtp_1 merge963 (.D(net370),
    .GATE(clknet_4_8_0_clk),
    .RESET_B(net786),
    .Q(net945));
 sky130_fd_sc_hd__edfxbp_1 merge964 (.CLK(clknet_4_7_0_clk),
    .D(net782),
    .DE(net890),
    .Q(net947),
    .Q_N(net946));
 sky130_fd_sc_hd__edfxtp_1 merge965 (.CLK(clknet_4_14_0_clk),
    .D(net743),
    .DE(net41),
    .Q(net948));
 sky130_fd_sc_hd__sdlclkp_1 merge966 (.CLK(clknet_4_3_0_clk),
    .GATE(net698),
    .SCE(net842),
    .GCLK(net949));
 sky130_fd_sc_hd__sdlclkp_2 merge967 (.CLK(clknet_4_12_0_clk),
    .GATE(net850),
    .SCE(net805),
    .GCLK(net950));
 sky130_fd_sc_hd__sdlclkp_4 merge968 (.CLK(clknet_4_14_0_clk),
    .GATE(net826),
    .SCE(net770),
    .GCLK(net951));
 sky130_fd_sc_hd__dfrbp_1 merge969 (.CLK(clknet_4_1_0_clk),
    .D(net857),
    .RESET_B(net537),
    .Q(net953),
    .Q_N(net952));
 sky130_fd_sc_hd__dfrbp_1 merge970 (.CLK(clknet_4_15_0_clk),
    .D(net796),
    .RESET_B(net894),
    .Q(net955),
    .Q_N(net954));
 sky130_fd_sc_hd__dfrtn_1 merge971 (.CLK_N(clknet_4_13_0_clk),
    .D(net899),
    .RESET_B(net897),
    .Q(net956));
 sky130_fd_sc_hd__dfrtp_4 merge972 (.CLK(clknet_4_3_0_clk),
    .D(net449),
    .RESET_B(net846),
    .Q(net957));
 sky130_fd_sc_hd__dfrtp_4 merge973 (.CLK(clknet_4_6_0_clk),
    .D(net779),
    .RESET_B(net918),
    .Q(net958));
 sky130_fd_sc_hd__dfrtp_1 merge974 (.CLK(clknet_4_11_0_clk),
    .D(net869),
    .RESET_B(net1041),
    .Q(net959));
 sky130_fd_sc_hd__dfsbp_1 merge975 (.CLK(clknet_4_1_0_clk),
    .D(net801),
    .SET_B(net865),
    .Q(net961),
    .Q_N(net960));
 sky130_fd_sc_hd__dfsbp_1 merge976 (.CLK(clknet_4_14_0_clk),
    .D(net77),
    .SET_B(net874),
    .Q(net963),
    .Q_N(net962));
 sky130_fd_sc_hd__dfstp_1 merge977 (.CLK(clknet_4_1_0_clk),
    .D(net810),
    .SET_B(net844),
    .Q(net964));
 sky130_fd_sc_hd__dfstp_1 merge978 (.CLK(clknet_4_6_0_clk),
    .D(net859),
    .SET_B(net881),
    .Q(net965));
 sky130_fd_sc_hd__dfstp_1 merge979 (.CLK(clknet_4_7_0_clk),
    .D(net804),
    .SET_B(net806),
    .Q(net966));
 sky130_fd_sc_hd__dlrbn_1 merge980 (.D(net695),
    .GATE_N(clknet_4_3_0_clk),
    .RESET_B(net790),
    .Q(net968),
    .Q_N(net967));
 sky130_fd_sc_hd__dlrbn_1 merge981 (.D(net893),
    .GATE_N(clknet_4_1_0_clk),
    .RESET_B(net713),
    .Q(net970),
    .Q_N(net969));
 sky130_fd_sc_hd__dlrbp_1 merge982 (.D(net763),
    .GATE(clknet_4_4_0_clk),
    .RESET_B(net829),
    .Q(net972),
    .Q_N(net971));
 sky130_fd_sc_hd__dlrbp_1 merge983 (.D(net812),
    .GATE(clknet_4_12_0_clk),
    .RESET_B(net848),
    .Q(net974),
    .Q_N(net973));
 sky130_fd_sc_hd__dlrtn_1 merge984 (.D(net583),
    .GATE_N(clknet_4_7_0_clk),
    .RESET_B(net754),
    .Q(net975));
 sky130_fd_sc_hd__dlrtn_1 merge985 (.D(net840),
    .GATE_N(clknet_4_13_0_clk),
    .RESET_B(net813),
    .Q(net976));
 sky130_fd_sc_hd__dlrtn_1 merge986 (.D(net864),
    .GATE_N(clknet_4_7_0_clk),
    .RESET_B(net1053),
    .Q(net977));
 sky130_fd_sc_hd__dlrtp_1 merge987 (.D(net895),
    .GATE(clknet_4_3_0_clk),
    .RESET_B(net794),
    .Q(net978));
 sky130_fd_sc_hd__dlrtp_1 merge988 (.D(net877),
    .GATE(clknet_4_15_0_clk),
    .RESET_B(net858),
    .Q(net979));
 sky130_fd_sc_hd__dlrtp_2 merge989 (.D(net838),
    .GATE(clknet_4_15_0_clk),
    .RESET_B(net847),
    .Q(net980));
 sky130_fd_sc_hd__edfxbp_1 merge990 (.CLK(clknet_4_8_0_clk),
    .D(net811),
    .DE(net825),
    .Q(net982),
    .Q_N(net981));
 sky130_fd_sc_hd__edfxtp_1 merge991 (.CLK(clknet_4_9_0_clk),
    .D(net866),
    .DE(net837),
    .Q(net983));
 sky130_fd_sc_hd__sdlclkp_1 merge992 (.CLK(clknet_4_12_0_clk),
    .GATE(net903),
    .SCE(net832),
    .GCLK(net984));
 sky130_fd_sc_hd__sdlclkp_2 merge993 (.CLK(clknet_4_11_0_clk),
    .GATE(net861),
    .SCE(net828),
    .GCLK(net985));
 sky130_fd_sc_hd__dlclkp_2 s1000 (.CLK(clknet_4_3_0_clk),
    .GATE(net693),
    .GCLK(net993));
 sky130_fd_sc_hd__dlclkp_4 s1001 (.CLK(clknet_4_5_0_clk),
    .GATE(net841),
    .GCLK(net994));
 sky130_fd_sc_hd__dfxbp_1 s994 (.CLK(clknet_4_11_0_clk),
    .D(net82),
    .Q(net987),
    .Q_N(net986));
 sky130_fd_sc_hd__dfxbp_1 s995 (.CLK(clknet_4_8_0_clk),
    .D(net246),
    .Q(net989),
    .Q_N(net988));
 sky130_fd_sc_hd__dfxtp_1 s996 (.CLK(clknet_4_13_0_clk),
    .D(net314),
    .Q(net990));
 sky130_fd_sc_hd__dfxtp_1 s997 (.CLK(clknet_4_3_0_clk),
    .D(net427),
    .Q(net991));
 sky130_fd_sc_hd__dfxtp_1 s998 (.CLK(clknet_4_7_0_clk),
    .D(net604),
    .Q(net992));
 sky130_fd_sc_hd__dlclkp_1 s999 (.CLK(clknet_4_5_0_clk),
    .GATE(net629),
    .GCLK(net1020));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Right_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Right_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Right_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Right_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Right_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Right_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Right_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Right_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Right_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Right_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Right_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Right_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Right_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Right_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Right_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Right_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Right_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Right_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Right_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Right_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Right_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_161 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_162 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_163 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_164 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_165 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_166 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_167 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_168 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_169 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_170 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_171 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_172 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_173 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_174 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_175 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_176 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_177 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_178 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_179 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_180 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_181 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_182 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Left_183 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Left_184 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Left_185 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Left_186 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Left_187 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Left_188 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Left_189 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Left_190 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Left_191 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Left_192 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Left_193 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Left_194 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Left_195 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Left_196 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Left_197 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Left_198 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Left_199 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Left_200 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Left_201 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Left_202 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Left_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1347 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(in0),
    .X(net556));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(in1),
    .X(net628));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(in10),
    .X(net759));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(in11),
    .X(net995));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(in12),
    .X(net996));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(in13),
    .X(net997));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(in14),
    .X(net998));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(in15),
    .X(net999));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(in16),
    .X(net1000));
 sky130_fd_sc_hd__buf_1 input10 (.A(in17),
    .X(net1001));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(in19),
    .X(net1002));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(in2),
    .X(net1003));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(in20),
    .X(net1004));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(in21),
    .X(net1005));
 sky130_fd_sc_hd__clkbuf_4 input15 (.A(in22),
    .X(net1006));
 sky130_fd_sc_hd__buf_1 input16 (.A(in23),
    .X(net1007));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(in24),
    .X(net1008));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(in3),
    .X(net1009));
 sky130_fd_sc_hd__clkbuf_1 input19 (.A(in4),
    .X(net1010));
 sky130_fd_sc_hd__clkbuf_1 input20 (.A(in5),
    .X(net1011));
 sky130_fd_sc_hd__buf_1 input21 (.A(in6),
    .X(net1012));
 sky130_fd_sc_hd__buf_1 input22 (.A(in7),
    .X(net1013));
 sky130_fd_sc_hd__clkbuf_1 input23 (.A(in8),
    .X(net1014));
 sky130_fd_sc_hd__clkbuf_1 input24 (.A(in9),
    .X(net1015));
 sky130_fd_sc_hd__buf_2 output25 (.A(net1016),
    .X(out0));
 sky130_fd_sc_hd__buf_2 output26 (.A(net1017),
    .X(out1));
 sky130_fd_sc_hd__clkbuf_1 output27 (.A(net1018),
    .X(out12));
 sky130_fd_sc_hd__buf_2 output28 (.A(net1019),
    .X(out13));
 sky130_fd_sc_hd__clkbuf_1 output29 (.A(clknet_1_0__leaf_net1020),
    .X(out14));
 sky130_fd_sc_hd__buf_2 output30 (.A(net1021),
    .X(out16));
 sky130_fd_sc_hd__buf_2 output31 (.A(net1022),
    .X(out19));
 sky130_fd_sc_hd__buf_2 output32 (.A(net1023),
    .X(out21));
 sky130_fd_sc_hd__buf_2 output33 (.A(net1024),
    .X(out22));
 sky130_fd_sc_hd__buf_2 output34 (.A(net1025),
    .X(out23));
 sky130_fd_sc_hd__buf_2 output35 (.A(net1026),
    .X(out24));
 sky130_fd_sc_hd__buf_2 output36 (.A(net1027),
    .X(out4));
 sky130_fd_sc_hd__buf_2 output37 (.A(net1028),
    .X(out5));
 sky130_fd_sc_hd__buf_2 output38 (.A(net1029),
    .X(out7));
 sky130_fd_sc_hd__buf_2 output39 (.A(net1030),
    .X(out9));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net1020 (.A(net1020),
    .X(clknet_0_net1020));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net1020 (.A(clknet_0_net1020),
    .X(clknet_1_0__leaf_net1020));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net1020 (.A(clknet_0_net1020),
    .X(clknet_1_1__leaf_net1020));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net994 (.A(net994),
    .X(clknet_0_net994));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net994 (.A(clknet_0_net994),
    .X(clknet_1_0__leaf_net994));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net994 (.A(clknet_0_net994),
    .X(clknet_1_1__leaf_net994));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net558 (.A(net558),
    .X(clknet_0_net558));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net558 (.A(clknet_0_net558),
    .X(clknet_1_0__leaf_net558));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net558 (.A(clknet_0_net558),
    .X(clknet_1_1__leaf_net558));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net563 (.A(net563),
    .X(clknet_0_net563));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net563 (.A(clknet_0_net563),
    .X(clknet_1_0__leaf_net563));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net563 (.A(clknet_0_net563),
    .X(clknet_1_1__leaf_net563));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net993 (.A(net993),
    .X(clknet_0_net993));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net993 (.A(clknet_0_net993),
    .X(clknet_1_0__leaf_net993));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net993 (.A(clknet_0_net993),
    .X(clknet_1_1__leaf_net993));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net694 (.A(net694),
    .X(clknet_0_net694));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net694 (.A(clknet_0_net694),
    .X(clknet_1_0__leaf_net694));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net694 (.A(clknet_0_net694),
    .X(clknet_1_1__leaf_net694));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net949 (.A(net949),
    .X(clknet_0_net949));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net949 (.A(clknet_0_net949),
    .X(clknet_1_0__leaf_net949));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net949 (.A(clknet_0_net949),
    .X(clknet_1_1__leaf_net949));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net710 (.A(net710),
    .X(clknet_0_net710));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net710 (.A(clknet_0_net710),
    .X(clknet_1_0__leaf_net710));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net710 (.A(clknet_0_net710),
    .X(clknet_1_1__leaf_net710));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net717 (.A(net717),
    .X(clknet_0_net717));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net717 (.A(clknet_0_net717),
    .X(clknet_1_0__leaf_net717));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net717 (.A(clknet_0_net717),
    .X(clknet_1_1__leaf_net717));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net719 (.A(net719),
    .X(clknet_0_net719));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net719 (.A(clknet_0_net719),
    .X(clknet_1_0__leaf_net719));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net719 (.A(clknet_0_net719),
    .X(clknet_1_1__leaf_net719));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net712 (.A(net712),
    .X(clknet_0_net712));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net712 (.A(clknet_0_net712),
    .X(clknet_1_0__leaf_net712));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net712 (.A(clknet_0_net712),
    .X(clknet_1_1__leaf_net712));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net442 (.A(net442),
    .X(clknet_0_net442));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net442 (.A(clknet_0_net442),
    .X(clknet_1_0__leaf_net442));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net442 (.A(clknet_0_net442),
    .X(clknet_1_1__leaf_net442));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net447 (.A(net447),
    .X(clknet_0_net447));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net447 (.A(clknet_0_net447),
    .X(clknet_1_0__leaf_net447));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net447 (.A(clknet_0_net447),
    .X(clknet_1_1__leaf_net447));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net914 (.A(net914),
    .X(clknet_0_net914));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net914 (.A(clknet_0_net914),
    .X(clknet_1_0__leaf_net914));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net914 (.A(clknet_0_net914),
    .X(clknet_1_1__leaf_net914));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net985 (.A(net985),
    .X(clknet_0_net985));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net985 (.A(clknet_0_net985),
    .X(clknet_1_0__leaf_net985));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net985 (.A(clknet_0_net985),
    .X(clknet_1_1__leaf_net985));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net984 (.A(net984),
    .X(clknet_0_net984));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net984 (.A(clknet_0_net984),
    .X(clknet_1_0__leaf_net984));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net984 (.A(clknet_0_net984),
    .X(clknet_1_1__leaf_net984));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net498 (.A(net498),
    .X(clknet_0_net498));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net498 (.A(clknet_0_net498),
    .X(clknet_1_0__leaf_net498));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net498 (.A(clknet_0_net498),
    .X(clknet_1_1__leaf_net498));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net357 (.A(net357),
    .X(clknet_0_net357));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net357 (.A(clknet_0_net357),
    .X(clknet_1_0__leaf_net357));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net357 (.A(clknet_0_net357),
    .X(clknet_1_1__leaf_net357));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net197 (.A(net197),
    .X(clknet_0_net197));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net197 (.A(clknet_0_net197),
    .X(clknet_1_0__leaf_net197));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net197 (.A(clknet_0_net197),
    .X(clknet_1_1__leaf_net197));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net201 (.A(net201),
    .X(clknet_0_net201));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net201 (.A(clknet_0_net201),
    .X(clknet_1_0__leaf_net201));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net201 (.A(clknet_0_net201),
    .X(clknet_1_1__leaf_net201));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net85 (.A(net85),
    .X(clknet_0_net85));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net85 (.A(clknet_0_net85),
    .X(clknet_1_0__leaf_net85));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net85 (.A(clknet_0_net85),
    .X(clknet_1_1__leaf_net85));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net205 (.A(net205),
    .X(clknet_0_net205));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net205 (.A(clknet_0_net205),
    .X(clknet_1_0__leaf_net205));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net205 (.A(clknet_0_net205),
    .X(clknet_1_1__leaf_net205));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net208 (.A(net208),
    .X(clknet_0_net208));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net208 (.A(clknet_0_net208),
    .X(clknet_1_0__leaf_net208));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net208 (.A(clknet_0_net208),
    .X(clknet_1_1__leaf_net208));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net226 (.A(net226),
    .X(clknet_0_net226));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net226 (.A(clknet_0_net226),
    .X(clknet_1_0__leaf_net226));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net226 (.A(clknet_0_net226),
    .X(clknet_1_1__leaf_net226));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net210 (.A(net210),
    .X(clknet_0_net210));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net210 (.A(clknet_0_net210),
    .X(clknet_1_0__leaf_net210));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net210 (.A(clknet_0_net210),
    .X(clknet_1_1__leaf_net210));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net207 (.A(net207),
    .X(clknet_0_net207));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net207 (.A(clknet_0_net207),
    .X(clknet_1_0__leaf_net207));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net207 (.A(clknet_0_net207),
    .X(clknet_1_1__leaf_net207));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net213 (.A(net213),
    .X(clknet_0_net213));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net213 (.A(clknet_0_net213),
    .X(clknet_1_0__leaf_net213));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net213 (.A(clknet_0_net213),
    .X(clknet_1_1__leaf_net213));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net87 (.A(net87),
    .X(clknet_0_net87));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net87 (.A(clknet_0_net87),
    .X(clknet_1_0__leaf_net87));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net87 (.A(clknet_0_net87),
    .X(clknet_1_1__leaf_net87));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net91 (.A(net91),
    .X(clknet_0_net91));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net91 (.A(clknet_0_net91),
    .X(clknet_1_0__leaf_net91));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net91 (.A(clknet_0_net91),
    .X(clknet_1_1__leaf_net91));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net89 (.A(net89),
    .X(clknet_0_net89));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net89 (.A(clknet_0_net89),
    .X(clknet_1_0__leaf_net89));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net89 (.A(clknet_0_net89),
    .X(clknet_1_1__leaf_net89));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net88 (.A(net88),
    .X(clknet_0_net88));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net88 (.A(clknet_0_net88),
    .X(clknet_1_0__leaf_net88));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net88 (.A(clknet_0_net88),
    .X(clknet_1_1__leaf_net88));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net95 (.A(net95),
    .X(clknet_0_net95));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net95 (.A(clknet_0_net95),
    .X(clknet_1_0__leaf_net95));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net95 (.A(clknet_0_net95),
    .X(clknet_1_1__leaf_net95));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net79 (.A(net79),
    .X(clknet_0_net79));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net79 (.A(clknet_0_net79),
    .X(clknet_1_0__leaf_net79));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net79 (.A(clknet_0_net79),
    .X(clknet_1_1__leaf_net79));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net81 (.A(net81),
    .X(clknet_0_net81));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net81 (.A(clknet_0_net81),
    .X(clknet_1_0__leaf_net81));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net81 (.A(clknet_0_net81),
    .X(clknet_1_1__leaf_net81));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net951 (.A(net951),
    .X(clknet_0_net951));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net951 (.A(clknet_0_net951),
    .X(clknet_1_0__leaf_net951));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net951 (.A(clknet_0_net951),
    .X(clknet_1_1__leaf_net951));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net42 (.A(net42),
    .X(clknet_0_net42));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net42 (.A(clknet_0_net42),
    .X(clknet_1_0__leaf_net42));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net42 (.A(clknet_0_net42),
    .X(clknet_1_1__leaf_net42));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net29 (.A(net29),
    .X(clknet_0_net29));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net29 (.A(clknet_0_net29),
    .X(clknet_1_0__leaf_net29));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net29 (.A(clknet_0_net29),
    .X(clknet_1_1__leaf_net29));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net912 (.A(net912),
    .X(clknet_0_net912));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net912 (.A(clknet_0_net912),
    .X(clknet_1_0__leaf_net912));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net912 (.A(clknet_0_net912),
    .X(clknet_1_1__leaf_net912));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net26 (.A(net26),
    .X(clknet_0_net26));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net26 (.A(clknet_0_net26),
    .X(clknet_1_0__leaf_net26));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net26 (.A(clknet_0_net26),
    .X(clknet_1_1__leaf_net26));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net21 (.A(net21),
    .X(clknet_0_net21));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net21 (.A(clknet_0_net21),
    .X(clknet_1_0__leaf_net21));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net21 (.A(clknet_0_net21),
    .X(clknet_1_1__leaf_net21));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net24 (.A(net24),
    .X(clknet_0_net24));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net24 (.A(clknet_0_net24),
    .X(clknet_1_0__leaf_net24));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net24 (.A(clknet_0_net24),
    .X(clknet_1_1__leaf_net24));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net20 (.A(net20),
    .X(clknet_0_net20));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net20 (.A(clknet_0_net20),
    .X(clknet_1_0__leaf_net20));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net20 (.A(clknet_0_net20),
    .X(clknet_1_1__leaf_net20));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net25 (.A(net25),
    .X(clknet_0_net25));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net25 (.A(clknet_0_net25),
    .X(clknet_1_0__leaf_net25));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net25 (.A(clknet_0_net25),
    .X(clknet_1_1__leaf_net25));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net23 (.A(net23),
    .X(clknet_0_net23));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net23 (.A(clknet_0_net23),
    .X(clknet_1_0__leaf_net23));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net23 (.A(clknet_0_net23),
    .X(clknet_1_1__leaf_net23));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net34 (.A(net34),
    .X(clknet_0_net34));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net34 (.A(clknet_0_net34),
    .X(clknet_1_0__leaf_net34));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net34 (.A(clknet_0_net34),
    .X(clknet_1_1__leaf_net34));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net161 (.A(net161),
    .X(clknet_0_net161));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net161 (.A(clknet_0_net161),
    .X(clknet_1_0__leaf_net161));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net161 (.A(clknet_0_net161),
    .X(clknet_1_1__leaf_net161));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net163 (.A(net163),
    .X(clknet_0_net163));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net163 (.A(clknet_0_net163),
    .X(clknet_1_0__leaf_net163));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net163 (.A(clknet_0_net163),
    .X(clknet_1_1__leaf_net163));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net168 (.A(net168),
    .X(clknet_0_net168));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net168 (.A(clknet_0_net168),
    .X(clknet_1_0__leaf_net168));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net168 (.A(clknet_0_net168),
    .X(clknet_1_1__leaf_net168));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net162 (.A(net162),
    .X(clknet_0_net162));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net162 (.A(clknet_0_net162),
    .X(clknet_1_0__leaf_net162));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net162 (.A(clknet_0_net162),
    .X(clknet_1_1__leaf_net162));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net27 (.A(net27),
    .X(clknet_0_net27));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net27 (.A(clknet_0_net27),
    .X(clknet_1_0__leaf_net27));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net27 (.A(clknet_0_net27),
    .X(clknet_1_1__leaf_net27));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net22 (.A(net22),
    .X(clknet_0_net22));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net22 (.A(clknet_0_net22),
    .X(clknet_1_0__leaf_net22));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net22 (.A(clknet_0_net22),
    .X(clknet_1_1__leaf_net22));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net352 (.A(net352),
    .X(clknet_0_net352));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net352 (.A(clknet_0_net352),
    .X(clknet_1_0__leaf_net352));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net352 (.A(clknet_0_net352),
    .X(clknet_1_1__leaf_net352));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net353 (.A(net353),
    .X(clknet_0_net353));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net353 (.A(clknet_0_net353),
    .X(clknet_1_0__leaf_net353));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net353 (.A(clknet_0_net353),
    .X(clknet_1_1__leaf_net353));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net950 (.A(net950),
    .X(clknet_0_net950));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net950 (.A(clknet_0_net950),
    .X(clknet_1_0__leaf_net950));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net950 (.A(clknet_0_net950),
    .X(clknet_1_1__leaf_net950));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net764 (.A(net764),
    .X(clknet_0_net764));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net764 (.A(clknet_0_net764),
    .X(clknet_1_0__leaf_net764));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net764 (.A(clknet_0_net764),
    .X(clknet_1_1__leaf_net764));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net482 (.A(net482),
    .X(clknet_0_net482));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net482 (.A(clknet_0_net482),
    .X(clknet_1_0__leaf_net482));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net482 (.A(clknet_0_net482),
    .X(clknet_1_1__leaf_net482));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net479 (.A(net479),
    .X(clknet_0_net479));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net479 (.A(clknet_0_net479),
    .X(clknet_1_0__leaf_net479));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net479 (.A(clknet_0_net479),
    .X(clknet_1_1__leaf_net479));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net491 (.A(net491),
    .X(clknet_0_net491));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net491 (.A(clknet_0_net491),
    .X(clknet_1_0__leaf_net491));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net491 (.A(clknet_0_net491),
    .X(clknet_1_1__leaf_net491));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net496 (.A(net496),
    .X(clknet_0_net496));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net496 (.A(clknet_0_net496),
    .X(clknet_1_0__leaf_net496));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net496 (.A(clknet_0_net496),
    .X(clknet_1_1__leaf_net496));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net493 (.A(net493),
    .X(clknet_0_net493));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net493 (.A(clknet_0_net493),
    .X(clknet_1_0__leaf_net493));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net493 (.A(clknet_0_net493),
    .X(clknet_1_1__leaf_net493));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net747 (.A(net747),
    .X(clknet_0_net747));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net747 (.A(clknet_0_net747),
    .X(clknet_1_0__leaf_net747));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net747 (.A(clknet_0_net747),
    .X(clknet_1_1__leaf_net747));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net318 (.A(net318),
    .X(clknet_0_net318));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net318 (.A(clknet_0_net318),
    .X(clknet_1_0__leaf_net318));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net318 (.A(clknet_0_net318),
    .X(clknet_1_1__leaf_net318));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net325 (.A(net325),
    .X(clknet_0_net325));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net325 (.A(clknet_0_net325),
    .X(clknet_1_0__leaf_net325));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net325 (.A(clknet_0_net325),
    .X(clknet_1_1__leaf_net325));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net320 (.A(net320),
    .X(clknet_0_net320));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net320 (.A(clknet_0_net320),
    .X(clknet_1_0__leaf_net320));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net320 (.A(clknet_0_net320),
    .X(clknet_1_1__leaf_net320));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net321 (.A(net321),
    .X(clknet_0_net321));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net321 (.A(clknet_0_net321),
    .X(clknet_1_0__leaf_net321));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net321 (.A(clknet_0_net321),
    .X(clknet_1_1__leaf_net321));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net317 (.A(net317),
    .X(clknet_0_net317));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net317 (.A(clknet_0_net317),
    .X(clknet_1_0__leaf_net317));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net317 (.A(clknet_0_net317),
    .X(clknet_1_1__leaf_net317));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net324 (.A(net324),
    .X(clknet_0_net324));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net324 (.A(clknet_0_net324),
    .X(clknet_1_0__leaf_net324));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net324 (.A(clknet_0_net324),
    .X(clknet_1_1__leaf_net324));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net329 (.A(net329),
    .X(clknet_0_net329));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net329 (.A(clknet_0_net329),
    .X(clknet_1_0__leaf_net329));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net329 (.A(clknet_0_net329),
    .X(clknet_1_1__leaf_net329));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net326 (.A(net326),
    .X(clknet_0_net326));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net326 (.A(clknet_0_net326),
    .X(clknet_1_0__leaf_net326));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net326 (.A(clknet_0_net326),
    .X(clknet_1_1__leaf_net326));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net330 (.A(net330),
    .X(clknet_0_net330));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net330 (.A(clknet_0_net330),
    .X(clknet_1_0__leaf_net330));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net330 (.A(clknet_0_net330),
    .X(clknet_1_1__leaf_net330));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net328 (.A(net328),
    .X(clknet_0_net328));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net328 (.A(clknet_0_net328),
    .X(clknet_1_0__leaf_net328));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net328 (.A(clknet_0_net328),
    .X(clknet_1_1__leaf_net328));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net915 (.A(net915),
    .X(clknet_0_net915));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net915 (.A(clknet_0_net915),
    .X(clknet_1_0__leaf_net915));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net915 (.A(clknet_0_net915),
    .X(clknet_1_1__leaf_net915));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net160 (.A(net160),
    .X(clknet_0_net160));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net160 (.A(clknet_0_net160),
    .X(clknet_1_0__leaf_net160));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net160 (.A(clknet_0_net160),
    .X(clknet_1_1__leaf_net160));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net144 (.A(net144),
    .X(clknet_0_net144));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net144 (.A(clknet_0_net144),
    .X(clknet_1_0__leaf_net144));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net144 (.A(clknet_0_net144),
    .X(clknet_1_1__leaf_net144));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net147 (.A(net147),
    .X(clknet_0_net147));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net147 (.A(clknet_0_net147),
    .X(clknet_1_0__leaf_net147));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net147 (.A(clknet_0_net147),
    .X(clknet_1_1__leaf_net147));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net145 (.A(net145),
    .X(clknet_0_net145));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net145 (.A(clknet_0_net145),
    .X(clknet_1_0__leaf_net145));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net145 (.A(clknet_0_net145),
    .X(clknet_1_1__leaf_net145));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net272 (.A(net272),
    .X(clknet_0_net272));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net272 (.A(clknet_0_net272),
    .X(clknet_1_0__leaf_net272));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net272 (.A(clknet_0_net272),
    .X(clknet_1_1__leaf_net272));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net126 (.A(net126),
    .X(clknet_0_net126));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net126 (.A(clknet_0_net126),
    .X(clknet_1_0__leaf_net126));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net126 (.A(clknet_0_net126),
    .X(clknet_1_1__leaf_net126));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net129 (.A(net129),
    .X(clknet_0_net129));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net129 (.A(clknet_0_net129),
    .X(clknet_1_0__leaf_net129));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net129 (.A(clknet_0_net129),
    .X(clknet_1_1__leaf_net129));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net127 (.A(net127),
    .X(clknet_0_net127));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net127 (.A(clknet_0_net127),
    .X(clknet_1_0__leaf_net127));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net127 (.A(clknet_0_net127),
    .X(clknet_1_1__leaf_net127));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer1 (.A(net902),
    .X(net1031));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer2 (.A(net1031),
    .X(net1032));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer3 (.A(net33),
    .X(net1033));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(net102),
    .X(net1034));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(net530),
    .X(net1035));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(net536),
    .X(net1036));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(net873),
    .X(net1037));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(net969),
    .X(net1038));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(net824),
    .X(net1039));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(net980),
    .X(net1040));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(net114),
    .X(net1041));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(net962),
    .X(net1042));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(net16),
    .X(net1043));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(net228),
    .X(net1044));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(net222),
    .X(net1045));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(net792),
    .X(net1046));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(net843),
    .X(net1047));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(net952),
    .X(net1048));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(net807),
    .X(net1049));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(net648),
    .X(net1050));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(net235),
    .X(net1051));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(net992),
    .X(net1052));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(net607),
    .X(net1053));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(net818),
    .X(net1054));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(net99),
    .X(net1055));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(net105),
    .X(net1056));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(net1021),
    .X(net1057));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(net280),
    .X(net1058));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(net871),
    .X(net1059));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(net555),
    .X(net1060));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(net924),
    .X(net1061));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(net539),
    .X(net1062));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(net889),
    .X(net1063));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(net891),
    .X(net1064));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(net229),
    .X(net1065));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(net986),
    .X(net1066));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(net578),
    .X(net1067));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(net380),
    .X(net1068));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(net802),
    .X(net1069));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(net451),
    .X(net1070));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_A (.DIODE(clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(in0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(in1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(in10));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(in11));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(in12));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(in13));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(in14));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(in15));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(in16));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(in17));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_A (.DIODE(in18));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(in19));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(in2));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(in20));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(in21));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(in22));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(in23));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(in24));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(in3));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(in4));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(in5));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(in6));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_A (.DIODE(in7));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_A (.DIODE(in8));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_A (.DIODE(in9));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge872_S0 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge785_A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_c134_X (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge874_A3 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge872_S1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c140_X (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge860_C_N (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge808_C (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge794_D_N (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge782_S1 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c59_SCD (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c42_A2 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c41_A3 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c38_D_N (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c37_X (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_S0 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge883_S1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge874_S1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge872_A3 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_S0 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_A2 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_X (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge880_S1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge865_A3 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge818_C_N (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge793_B (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_A3 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_SET_B (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_X (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_A (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_B (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_Q (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge884_A1 (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge840_B (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge824_B (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge822_B (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_S1 (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA_c323_S0 (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_X (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge868_A2 (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge833_A (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_D_N (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_A (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_C (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_X (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_C_N (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_B (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_A (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA_c373_X (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge881_A2 (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge870_S0 (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge861_DE (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge841_A (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA_c395_S1 (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA_c392_C1 (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA_c385_C_N (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA_c383_A (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA_c375_X (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge871_A1 (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge870_S1 (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge862_A2 (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge841_B (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA_c385_B (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA_c378_X (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge814_A2 (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA_c507_B (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA_c394_Q_N (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA_c513_B (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA_c511_A (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA_c395_A3 (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA_c394_Q (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA_c404_B (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA_c403_A (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA_c397_A (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_X (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA_c563_C (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_A (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA_c416_X (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge792_D (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_X (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_A3 (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_C (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA_c431_A (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_B (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_B (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_B (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_B (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_A (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_X (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge883_A1 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_A1 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_B (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_B (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_B (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_C_N (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_B (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_A (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_X (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge859_D_N (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge858_SCD (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge855_B (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_A1 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_X (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge853_SCD (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_C (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_A (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_S0 (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_S0 (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_X (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge867_A1 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_c88_A (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_c70_B (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_c67_A (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_c66_X (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_A (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_c107_A2 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_c105_S1 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge810_B (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_A (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA_c482_C (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_S0 (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_D1 (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_A3 (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_B (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_X (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge926_A (.DIODE(net494));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_X (.DIODE(net494));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge882_A1 (.DIODE(net509));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge869_A3 (.DIODE(net509));
 sky130_fd_sc_hd__diode_2 ANTENNA_c525_B (.DIODE(net509));
 sky130_fd_sc_hd__diode_2 ANTENNA_c523_B (.DIODE(net509));
 sky130_fd_sc_hd__diode_2 ANTENNA_c522_C (.DIODE(net509));
 sky130_fd_sc_hd__diode_2 ANTENNA_c521_A (.DIODE(net509));
 sky130_fd_sc_hd__diode_2 ANTENNA_c519_X (.DIODE(net509));
 sky130_fd_sc_hd__diode_2 ANTENNA_c657_S1 (.DIODE(net510));
 sky130_fd_sc_hd__diode_2 ANTENNA_c655_A (.DIODE(net510));
 sky130_fd_sc_hd__diode_2 ANTENNA_c654_C_N (.DIODE(net510));
 sky130_fd_sc_hd__diode_2 ANTENNA_c527_C (.DIODE(net510));
 sky130_fd_sc_hd__diode_2 ANTENNA_c524_B (.DIODE(net510));
 sky130_fd_sc_hd__diode_2 ANTENNA_c521_C (.DIODE(net510));
 sky130_fd_sc_hd__diode_2 ANTENNA_c520_X (.DIODE(net510));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge829_SCD (.DIODE(net523));
 sky130_fd_sc_hd__diode_2 ANTENNA_c541_A (.DIODE(net523));
 sky130_fd_sc_hd__diode_2 ANTENNA_c533_X (.DIODE(net523));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge829_D (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA_c543_A2 (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA_c538_D (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA_c534_X (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge807_SCD (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA_c564_B (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA_c556_A (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA_c555_B (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA_c544_B (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA_c540_C (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA_c539_SCD (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA_c535_X (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net563_A (.DIODE(net563));
 sky130_fd_sc_hd__diode_2 ANTENNA_c571_X (.DIODE(net563));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge879_A2 (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_B1 (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_B1 (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_C (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_A (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_B (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_A (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_X (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge887_A2 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge846_B (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge803_C (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_c87_B1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_c86_D_N (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_c80_X (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_c101_A (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge814_A0 (.DIODE(net589));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_B (.DIODE(net589));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_SCD (.DIODE(net589));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_X (.DIODE(net589));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge817_A (.DIODE(net601));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_X (.DIODE(net601));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge863_A (.DIODE(net669));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_C_N (.DIODE(net669));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_B (.DIODE(net669));
 sky130_fd_sc_hd__diode_2 ANTENNA_c698_C (.DIODE(net669));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_X (.DIODE(net669));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge872_A0 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge851_A (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge846_D_N (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge804_B (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA_c90_X (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA_c106_D_N (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA_c100_B (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge880_A2 (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge830_B (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA_c747_A3 (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA_c742_RESET_B (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_A (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_S0 (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_B (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_B (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_B (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_X (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A (.DIODE(net720));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_A (.DIODE(net720));
 sky130_fd_sc_hd__diode_2 ANTENNA_c747_A2 (.DIODE(net720));
 sky130_fd_sc_hd__diode_2 ANTENNA_c746_X (.DIODE(net720));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge935_D (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge857_X (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge989_RESET_B (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge881_X (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge959_D (.DIODE(net853));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge887_X (.DIODE(net853));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge971_D (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge927_X (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge946_Q (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge869_S0 (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_A (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_A (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold31_A (.DIODE(net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge948_Q (.DIODE(net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge852_D_N (.DIODE(net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_c703_D_N (.DIODE(net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge951_Q (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge799_A (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c42_C1 (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c41_S1 (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_A (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge959_Q (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c85_A (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c82_A (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_A (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_A (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge960_Q (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c513_C (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c240_C (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_A (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_A (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge961_Q (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge849_D1 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c586_A (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_D_N (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_A (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge962_Q (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge815_A (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_c526_A (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_A (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_A (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge964_Q (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c194_A (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_A (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge972_Q (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_A (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_B (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_S1 (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_A (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge973_Q (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge869_S1 (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge805_A (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c525_D_N (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_A (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge976_Q (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge862_D1 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c101_C (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge977_Q (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c744_A (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_A (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c693_A (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c582_A (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge984_Q (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_A (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_D1 (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c159_A (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_A (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge986_Q (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_B (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_B (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_D1 (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_S1 (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge988_Q (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge867_S1 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c62_D1 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_D1 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_C (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold10_A (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge989_Q (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge809_A (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c382_A (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_A (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge991_Q (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c746_A (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c384_A (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c369_A (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_B (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_s996_Q (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge884_S1 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_B (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_D_N (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_D_N (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_s997_Q (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge801_C (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_B (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_A (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_X (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge808_B (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c56_C1 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c42_B1 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c37_C (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c34_SCE (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c32_D_N (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c27_B (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c25_B (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_A (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_X (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge880_A3 (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_output35_A (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c514_X (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_15_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_14_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_13_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_12_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_11_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_10_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_9_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_8_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_7_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_6_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_5_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_4_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_3_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_2_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_1_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_0_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_X (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c767_CLK_N (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge932_GATE_N (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge937_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge944_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge969_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge975_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge977_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge981_GATE_N (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_1_0_clk_X (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c656_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge900_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge905_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge914_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge945_CLK_N (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge961_GATE (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge982_GATE (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_4_0_clk_X (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_CLK_N (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c494_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c518_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge946_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge954_GATE_N (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge959_GATE_N (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge973_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge978_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_6_0_clk_X (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c610_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge902_CLK_N (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge920_GATE (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge935_GATE (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge941_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge957_GATE (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge964_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge979_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge984_GATE_N (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge986_GATE_N (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s998_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_7_0_clk_X (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c394_CLK_N (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge861_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge938_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge947_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge950_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge953_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge955_GATE_N (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge991_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_9_0_clk_X (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c237_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c34_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge816_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge909_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge928_GATE (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge951_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge952_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge965_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge968_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge976_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_14_0_clk_X (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge825_SCD (.DIODE(clknet_1_0__leaf_net563));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge836_B (.DIODE(clknet_1_0__leaf_net563));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net563_X (.DIODE(clknet_1_0__leaf_net563));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge797_SCD (.DIODE(clknet_1_1__leaf_net563));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge852_C_N (.DIODE(clknet_1_1__leaf_net563));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge879_A1 (.DIODE(clknet_1_1__leaf_net563));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net563_X (.DIODE(clknet_1_1__leaf_net563));
 sky130_fd_sc_hd__diode_2 ANTENNA_c369_B (.DIODE(clknet_1_0__leaf_net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c508_B (.DIODE(clknet_1_0__leaf_net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net984_X (.DIODE(clknet_1_0__leaf_net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c286_B (.DIODE(clknet_1_0__leaf_net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge880_S0 (.DIODE(clknet_1_0__leaf_net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net145_X (.DIODE(clknet_1_0__leaf_net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(net575));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_439 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_355 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_466 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_441 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_199 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_497 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_400 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_497 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_359 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_544 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_540 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_484 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_468 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_494 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_359 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_522 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_534 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_542 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_282 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_598 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_608 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_593 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_588 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_487 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_508 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_563 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_301 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_522 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_565 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_552 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_273 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_522 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_441 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_574 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_582 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_283 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_462 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_413 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_327 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_357 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_568 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_576 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_384 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_454 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_252 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_280 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_410 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_547 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_584 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_592 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_256 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_594 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_588 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_612 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_407 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_301 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_284 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_539 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_328 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_535 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_536 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_518 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_274 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_510 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_518 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_245 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_546 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_282 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_552 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_490 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_518 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_273 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_338 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_196 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_413 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_459 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_617 ();
endmodule
