module netlist_0 (clk,
    in0,
    in1,
    in10,
    in11,
    in12,
    in13,
    in14,
    in15,
    in16,
    in17,
    in18,
    in19,
    in2,
    in20,
    in21,
    in22,
    in23,
    in24,
    in25,
    in26,
    in27,
    in28,
    in29,
    in3,
    in30,
    in31,
    in32,
    in33,
    in34,
    in35,
    in36,
    in37,
    in38,
    in39,
    in4,
    in40,
    in41,
    in42,
    in43,
    in44,
    in45,
    in46,
    in47,
    in48,
    in49,
    in5,
    in50,
    in51,
    in52,
    in53,
    in54,
    in55,
    in56,
    in57,
    in58,
    in59,
    in6,
    in60,
    in61,
    in62,
    in63,
    in64,
    in65,
    in66,
    in67,
    in68,
    in69,
    in7,
    in70,
    in71,
    in72,
    in73,
    in74,
    in75,
    in76,
    in77,
    in78,
    in79,
    in8,
    in80,
    in81,
    in82,
    in83,
    in84,
    in85,
    in86,
    in87,
    in88,
    in89,
    in9,
    in90,
    in91,
    in92,
    in93,
    in94,
    in95,
    in96,
    in97,
    in98,
    in99,
    out0,
    out1,
    out10,
    out11,
    out12,
    out13,
    out14,
    out15,
    out16,
    out17,
    out18,
    out19,
    out2,
    out20,
    out21,
    out22,
    out23,
    out24,
    out25,
    out26,
    out27,
    out28,
    out29,
    out3,
    out30,
    out31,
    out32,
    out33,
    out34,
    out35,
    out36,
    out37,
    out38,
    out39,
    out4,
    out40,
    out41,
    out42,
    out43,
    out44,
    out45,
    out46,
    out47,
    out48,
    out49,
    out5,
    out50,
    out51,
    out52,
    out53,
    out54,
    out55,
    out56,
    out57,
    out58,
    out59,
    out6,
    out60,
    out61,
    out62,
    out63,
    out64,
    out65,
    out66,
    out67,
    out68,
    out69,
    out7,
    out70,
    out71,
    out72,
    out73,
    out74,
    out75,
    out76,
    out77,
    out78,
    out79,
    out8,
    out80,
    out81,
    out82,
    out83,
    out84,
    out85,
    out86,
    out87,
    out88,
    out89,
    out9,
    out90,
    out91,
    out92,
    out93,
    out94,
    out95,
    out96,
    out97,
    out98,
    out99,
    rst);
 input clk;
 input in0;
 input in1;
 input in10;
 input in11;
 input in12;
 input in13;
 input in14;
 input in15;
 input in16;
 input in17;
 input in18;
 input in19;
 input in2;
 input in20;
 input in21;
 input in22;
 input in23;
 input in24;
 input in25;
 input in26;
 input in27;
 input in28;
 input in29;
 input in3;
 input in30;
 input in31;
 input in32;
 input in33;
 input in34;
 input in35;
 input in36;
 input in37;
 input in38;
 input in39;
 input in4;
 input in40;
 input in41;
 input in42;
 input in43;
 input in44;
 input in45;
 input in46;
 input in47;
 input in48;
 input in49;
 input in5;
 input in50;
 input in51;
 input in52;
 input in53;
 input in54;
 input in55;
 input in56;
 input in57;
 input in58;
 input in59;
 input in6;
 input in60;
 input in61;
 input in62;
 input in63;
 input in64;
 input in65;
 input in66;
 input in67;
 input in68;
 input in69;
 input in7;
 input in70;
 input in71;
 input in72;
 input in73;
 input in74;
 input in75;
 input in76;
 input in77;
 input in78;
 input in79;
 input in8;
 input in80;
 input in81;
 input in82;
 input in83;
 input in84;
 input in85;
 input in86;
 input in87;
 input in88;
 input in89;
 input in9;
 input in90;
 input in91;
 input in92;
 input in93;
 input in94;
 input in95;
 input in96;
 input in97;
 input in98;
 input in99;
 output out0;
 output out1;
 output out10;
 output out11;
 output out12;
 output out13;
 output out14;
 output out15;
 output out16;
 output out17;
 output out18;
 output out19;
 output out2;
 output out20;
 output out21;
 output out22;
 output out23;
 output out24;
 output out25;
 output out26;
 output out27;
 output out28;
 output out29;
 output out3;
 output out30;
 output out31;
 output out32;
 output out33;
 output out34;
 output out35;
 output out36;
 output out37;
 output out38;
 output out39;
 output out4;
 output out40;
 output out41;
 output out42;
 output out43;
 output out44;
 output out45;
 output out46;
 output out47;
 output out48;
 output out49;
 output out5;
 output out50;
 output out51;
 output out52;
 output out53;
 output out54;
 output out55;
 output out56;
 output out57;
 output out58;
 output out59;
 output out6;
 output out60;
 output out61;
 output out62;
 output out63;
 output out64;
 output out65;
 output out66;
 output out67;
 output out68;
 output out69;
 output out7;
 output out70;
 output out71;
 output out72;
 output out73;
 output out74;
 output out75;
 output out76;
 output out77;
 output out78;
 output out79;
 output out8;
 output out80;
 output out81;
 output out82;
 output out83;
 output out84;
 output out85;
 output out86;
 output out87;
 output out88;
 output out89;
 output out9;
 output out90;
 output out91;
 output out92;
 output out93;
 output out94;
 output out95;
 output out96;
 output out97;
 output out98;
 output out99;
 input rst;

 wire net0;
 wire net1;
 wire net10;
 wire net100;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net63;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net64;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net65;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net66;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net67;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net68;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net69;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net7;
 wire net70;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net71;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net72;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net101;
 wire net192;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_0_net713;
 wire clknet_1_0__leaf_net713;
 wire clknet_1_1__leaf_net713;
 wire clknet_0_net712;
 wire clknet_1_0__leaf_net712;
 wire clknet_1_1__leaf_net712;
 wire clknet_0_net711;
 wire clknet_1_0__leaf_net711;
 wire clknet_1_1__leaf_net711;
 wire clknet_0_net458;
 wire clknet_1_0__leaf_net458;
 wire clknet_1_1__leaf_net458;
 wire clknet_0_net482;
 wire clknet_1_0__leaf_net482;
 wire clknet_1_1__leaf_net482;
 wire clknet_0_net609;
 wire clknet_1_0__leaf_net609;
 wire clknet_1_1__leaf_net609;
 wire clknet_0_net483;
 wire clknet_1_0__leaf_net483;
 wire clknet_1_1__leaf_net483;
 wire clknet_0_net452;
 wire clknet_1_0__leaf_net452;
 wire clknet_1_1__leaf_net452;
 wire clknet_0_net457;
 wire clknet_1_0__leaf_net457;
 wire clknet_1_1__leaf_net457;
 wire clknet_0_net437;
 wire clknet_1_0__leaf_net437;
 wire clknet_1_1__leaf_net437;
 wire clknet_0_net454;
 wire clknet_1_0__leaf_net454;
 wire clknet_1_1__leaf_net454;
 wire clknet_0_net450;
 wire clknet_1_0__leaf_net450;
 wire clknet_1_1__leaf_net450;
 wire clknet_0_net444;
 wire clknet_1_0__leaf_net444;
 wire clknet_1_1__leaf_net444;
 wire clknet_0_net435;
 wire clknet_1_0__leaf_net435;
 wire clknet_1_1__leaf_net435;
 wire clknet_0_net451;
 wire clknet_1_0__leaf_net451;
 wire clknet_1_1__leaf_net451;
 wire clknet_0_net693;
 wire clknet_1_0__leaf_net693;
 wire clknet_1_1__leaf_net693;
 wire clknet_0_net345;
 wire clknet_1_0__leaf_net345;
 wire clknet_1_1__leaf_net345;
 wire clknet_0_net577;
 wire clknet_1_0__leaf_net577;
 wire clknet_1_1__leaf_net577;
 wire clknet_0_net466;
 wire clknet_1_0__leaf_net466;
 wire clknet_1_1__leaf_net466;
 wire clknet_0_net338;
 wire clknet_1_0__leaf_net338;
 wire clknet_1_1__leaf_net338;
 wire clknet_0_net343;
 wire clknet_1_0__leaf_net343;
 wire clknet_1_1__leaf_net343;
 wire clknet_0_net692;
 wire clknet_1_0__leaf_net692;
 wire clknet_1_1__leaf_net692;
 wire clknet_0_net691;
 wire clknet_1_0__leaf_net691;
 wire clknet_1_1__leaf_net691;
 wire clknet_0_net673;
 wire clknet_1_0__leaf_net673;
 wire clknet_1_1__leaf_net673;
 wire clknet_0_net463;
 wire clknet_1_0__leaf_net463;
 wire clknet_1_1__leaf_net463;
 wire clknet_0_net426;
 wire clknet_1_0__leaf_net426;
 wire clknet_1_1__leaf_net426;
 wire clknet_0_net428;
 wire clknet_1_0__leaf_net428;
 wire clknet_1_1__leaf_net428;
 wire clknet_0_net429;
 wire clknet_1_0__leaf_net429;
 wire clknet_1_1__leaf_net429;
 wire clknet_0_net316;
 wire clknet_1_0__leaf_net316;
 wire clknet_1_1__leaf_net316;
 wire clknet_0_net448;
 wire clknet_1_0__leaf_net448;
 wire clknet_1_1__leaf_net448;
 wire clknet_0_net610;
 wire clknet_1_0__leaf_net610;
 wire clknet_1_1__leaf_net610;
 wire clknet_0_net318;
 wire clknet_1_0__leaf_net318;
 wire clknet_1_1__leaf_net318;
 wire clknet_0_net440;
 wire clknet_1_0__leaf_net440;
 wire clknet_1_1__leaf_net440;
 wire clknet_0_net321;
 wire clknet_1_0__leaf_net321;
 wire clknet_1_1__leaf_net321;
 wire clknet_0_net315;
 wire clknet_1_0__leaf_net315;
 wire clknet_1_1__leaf_net315;
 wire clknet_0_net400;
 wire clknet_1_0__leaf_net400;
 wire clknet_1_1__leaf_net400;
 wire clknet_0_net349;
 wire clknet_1_0__leaf_net349;
 wire clknet_1_1__leaf_net349;
 wire clknet_0_net317;
 wire clknet_1_0__leaf_net317;
 wire clknet_1_1__leaf_net317;
 wire clknet_0_net367;
 wire clknet_1_0__leaf_net367;
 wire clknet_1_1__leaf_net367;
 wire clknet_0_net492;
 wire clknet_1_0__leaf_net492;
 wire clknet_1_1__leaf_net492;
 wire clknet_0_net672;
 wire clknet_1_0__leaf_net672;
 wire clknet_1_1__leaf_net672;
 wire clknet_0_net290;
 wire clknet_1_0__leaf_net290;
 wire clknet_1_1__leaf_net290;
 wire clknet_0_net671;
 wire clknet_1_0__leaf_net671;
 wire clknet_1_1__leaf_net671;
 wire clknet_0_net276;
 wire clknet_1_0__leaf_net276;
 wire clknet_1_1__leaf_net276;
 wire clknet_0_net653;
 wire clknet_1_0__leaf_net653;
 wire clknet_1_1__leaf_net653;
 wire clknet_0_net296;
 wire clknet_1_0__leaf_net296;
 wire clknet_1_1__leaf_net296;
 wire clknet_0_net292;
 wire clknet_1_0__leaf_net292;
 wire clknet_1_1__leaf_net292;
 wire clknet_0_net652;
 wire clknet_1_0__leaf_net652;
 wire clknet_1_1__leaf_net652;
 wire clknet_0_net866;
 wire clknet_1_0__leaf_net866;
 wire clknet_1_1__leaf_net866;
 wire clknet_0_net860;
 wire clknet_1_0__leaf_net860;
 wire clknet_1_1__leaf_net860;
 wire clknet_0_net853;
 wire clknet_1_0__leaf_net853;
 wire clknet_1_1__leaf_net853;
 wire clknet_0_net651;
 wire clknet_1_0__leaf_net651;
 wire clknet_1_1__leaf_net651;
 wire clknet_0_net177;
 wire clknet_1_0__leaf_net177;
 wire clknet_1_1__leaf_net177;
 wire clknet_0_net385;
 wire clknet_1_0__leaf_net385;
 wire clknet_1_1__leaf_net385;
 wire clknet_0_net176;
 wire clknet_1_0__leaf_net176;
 wire clknet_1_1__leaf_net176;
 wire clknet_0_net836;
 wire clknet_1_0__leaf_net836;
 wire clknet_1_1__leaf_net836;
 wire clknet_0_net281;
 wire clknet_1_0__leaf_net281;
 wire clknet_1_1__leaf_net281;
 wire clknet_0_net174;
 wire clknet_1_0__leaf_net174;
 wire clknet_1_1__leaf_net174;
 wire clknet_0_net371;
 wire clknet_1_0__leaf_net371;
 wire clknet_1_1__leaf_net371;
 wire clknet_0_net386;
 wire clknet_1_0__leaf_net386;
 wire clknet_1_1__leaf_net386;
 wire clknet_0_net173;
 wire clknet_1_0__leaf_net173;
 wire clknet_1_1__leaf_net173;
 wire clknet_0_net571;
 wire clknet_1_0__leaf_net571;
 wire clknet_1_1__leaf_net571;
 wire clknet_0_net189;
 wire clknet_1_0__leaf_net189;
 wire clknet_1_1__leaf_net189;
 wire clknet_0_net180;
 wire clknet_1_0__leaf_net180;
 wire clknet_1_1__leaf_net180;
 wire clknet_0_net155;
 wire clknet_1_0__leaf_net155;
 wire clknet_1_1__leaf_net155;
 wire clknet_0_net459;
 wire clknet_1_0__leaf_net459;
 wire clknet_1_1__leaf_net459;
 wire clknet_0_net250;
 wire clknet_1_0__leaf_net250;
 wire clknet_1_1__leaf_net250;
 wire clknet_0_net359;
 wire clknet_1_0__leaf_net359;
 wire clknet_1_1__leaf_net359;
 wire clknet_0_net355;
 wire clknet_1_0__leaf_net355;
 wire clknet_1_1__leaf_net355;
 wire clknet_0_net855;
 wire clknet_1_0__leaf_net855;
 wire clknet_1_1__leaf_net855;
 wire clknet_0_net632;
 wire clknet_1_0__leaf_net632;
 wire clknet_1_1__leaf_net632;
 wire clknet_0_net96;
 wire clknet_1_0__leaf_net96;
 wire clknet_1_1__leaf_net96;
 wire clknet_0_net868;
 wire clknet_1_0__leaf_net868;
 wire clknet_1_1__leaf_net868;
 wire clknet_0_net631;
 wire clknet_1_0__leaf_net631;
 wire clknet_1_1__leaf_net631;
 wire clknet_0_net875;
 wire clknet_1_0__leaf_net875;
 wire clknet_1_1__leaf_net875;
 wire clknet_0_net851;
 wire clknet_1_0__leaf_net851;
 wire clknet_1_1__leaf_net851;
 wire clknet_0_net84;
 wire clknet_1_0__leaf_net84;
 wire clknet_1_1__leaf_net84;
 wire clknet_0_net183;
 wire clknet_1_0__leaf_net183;
 wire clknet_1_1__leaf_net183;
 wire clknet_0_net834;
 wire clknet_1_0__leaf_net834;
 wire clknet_1_1__leaf_net834;
 wire clknet_0_net86;
 wire clknet_1_0__leaf_net86;
 wire clknet_1_1__leaf_net86;
 wire clknet_0_net78;
 wire clknet_1_0__leaf_net78;
 wire clknet_1_1__leaf_net78;
 wire clknet_0_net93;
 wire clknet_1_0__leaf_net93;
 wire clknet_1_1__leaf_net93;
 wire clknet_0_net630;
 wire clknet_1_0__leaf_net630;
 wire clknet_1_1__leaf_net630;
 wire clknet_0_net389;
 wire clknet_1_0__leaf_net389;
 wire clknet_1_1__leaf_net389;
 wire clknet_0_net844;
 wire clknet_1_0__leaf_net844;
 wire clknet_1_1__leaf_net844;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;

 sky130_fd_sc_hd__mux4_1 c100 (.A0(net740),
    .A1(net812),
    .A2(net818),
    .A3(net820),
    .S0(net821),
    .S1(net813),
    .X(net0));
 sky130_fd_sc_hd__mux4_2 c101 (.A0(net783),
    .A1(net810),
    .A2(net819),
    .A3(net814),
    .S0(net797),
    .S1(net792),
    .X(net863));
 sky130_fd_sc_hd__mux4_2 c102 (.A0(net815),
    .A1(net746),
    .A2(net820),
    .A3(net819),
    .S0(net972),
    .S1(net775),
    .X(net1));
 sky130_fd_sc_hd__mux4_2 c103 (.A0(net819),
    .A1(net802),
    .A2(net1023),
    .A3(net820),
    .S0(net863),
    .S1(net817),
    .X(net2));
 sky130_fd_sc_hd__mux4_2 c104 (.A0(net820),
    .A1(net815),
    .A2(net821),
    .A3(net818),
    .S0(net1),
    .S1(net2),
    .X(net3));
 sky130_fd_sc_hd__mux4_1 c105 (.A0(net2),
    .A1(net819),
    .A2(net1),
    .A3(net818),
    .S0(net813),
    .S1(net812),
    .X(net4));
 sky130_fd_sc_hd__mux4_1 c106 (.A0(net803),
    .A1(net809),
    .A2(net795),
    .A3(net802),
    .S0(net819),
    .S1(net1),
    .X(net882));
 sky130_fd_sc_hd__mux4_2 c107 (.A0(net816),
    .A1(net802),
    .A2(net818),
    .A3(net815),
    .S0(net956),
    .S1(net950),
    .X(net879));
 sky130_fd_sc_hd__mux4_1 c108 (.A0(net882),
    .A1(net980),
    .A2(net4),
    .A3(net958),
    .S0(net2),
    .S1(net820),
    .X(net876));
 sky130_fd_sc_hd__mux4_2 c109 (.A0(net766),
    .A1(net2),
    .A2(net783),
    .A3(net876),
    .S0(net814),
    .S1(net785),
    .X(net887));
 sky130_fd_sc_hd__mux4_1 c122 (.A0(net806),
    .A1(net785),
    .A2(net771),
    .A3(net765),
    .S0(net950),
    .S1(net887),
    .X(net840));
 sky130_fd_sc_hd__mux4_1 c123 (.A0(net727),
    .A1(net819),
    .A2(net802),
    .A3(net768),
    .S0(net821),
    .S1(net882),
    .X(net886));
 sky130_fd_sc_hd__mux4_1 c124 (.A0(net758),
    .A1(net765),
    .A2(net1041),
    .A3(net780),
    .S0(net776),
    .S1(net950),
    .X(net877));
 sky130_fd_sc_hd__mux4_1 c125 (.A0(net2),
    .A1(net887),
    .A2(net863),
    .A3(net806),
    .S0(net879),
    .S1(net968),
    .X(net885));
 sky130_fd_sc_hd__mux4_2 c126 (.A0(net819),
    .A1(net877),
    .A2(net820),
    .A3(net808),
    .S0(net787),
    .S1(net950),
    .X(net854));
 sky130_fd_sc_hd__mux4_1 c127 (.A0(net771),
    .A1(net840),
    .A2(net854),
    .A3(net885),
    .S0(net768),
    .S1(net2),
    .X(net5));
 sky130_fd_sc_hd__mux4_1 c128 (.A0(net820),
    .A1(net854),
    .A2(net785),
    .A3(net5),
    .S0(net809),
    .S1(net819),
    .X(net883));
 sky130_fd_sc_hd__mux4_1 c129 (.A0(net751),
    .A1(net749),
    .A2(net883),
    .A3(net806),
    .S0(net780),
    .S1(net854),
    .X(net878));
 sky130_fd_sc_hd__mux4_1 c130 (.A0(net5),
    .A1(net727),
    .A2(net878),
    .A3(net785),
    .S0(net854),
    .S1(net885),
    .X(net823));
 sky130_fd_sc_hd__mux4_1 c131 (.A0(net768),
    .A1(net820),
    .A2(net854),
    .A3(net823),
    .S0(net808),
    .S1(net776),
    .X(net870));
 sky130_fd_sc_hd__a41o_4 c132 (.A1(net977),
    .A2(net974),
    .A3(net959),
    .A4(net967),
    .B1(net727),
    .X(net6));
 sky130_fd_sc_hd__a41o_4 c133 (.A1(net948),
    .A2(net1041),
    .A3(net1023),
    .A4(net1022),
    .B1(net1021),
    .X(net7));
 sky130_fd_sc_hd__a41o_4 c134 (.A1(net7),
    .A2(net959),
    .A3(net6),
    .A4(net965),
    .B1(net735),
    .X(net8));
 sky130_fd_sc_hd__a41o_4 c135 (.A1(net937),
    .A2(net952),
    .A3(net1041),
    .A4(net7),
    .B1(net968),
    .X(net822));
 sky130_fd_sc_hd__mux4_2 c136 (.A0(net1042),
    .A1(net745),
    .A2(net1021),
    .A3(net979),
    .S0(net7),
    .S1(net1023),
    .X(net9));
 sky130_fd_sc_hd__a41o_2 c137 (.A1(net932),
    .A2(net971),
    .A3(net1042),
    .A4(net965),
    .B1(net1021),
    .X(net10));
 sky130_fd_sc_hd__a41o_1 c138 (.A1(net964),
    .A2(net937),
    .A3(net1021),
    .A4(net1022),
    .B1(net952),
    .X(net11));
 sky130_fd_sc_hd__a41o_4 c139 (.A1(net979),
    .A2(net7),
    .A3(net961),
    .A4(net965),
    .B1(net952),
    .X(net12));
 sky130_fd_sc_hd__a41o_4 c140 (.A1(net932),
    .A2(net972),
    .A3(net1022),
    .A4(net965),
    .B1(net974),
    .X(net872));
 sky130_fd_sc_hd__a41o_4 c141 (.A1(net930),
    .A2(net11),
    .A3(net980),
    .A4(net1022),
    .B1(net1021),
    .X(net13));
 sky130_fd_sc_hd__a41o_4 c142 (.A1(net927),
    .A2(net932),
    .A3(net930),
    .A4(net1021),
    .B1(net979),
    .X(net14));
 sky130_fd_sc_hd__a41o_2 c143 (.A1(net930),
    .A2(net11),
    .A3(net965),
    .A4(net6),
    .B1(net12),
    .X(net15));
 sky130_fd_sc_hd__mux4_2 c144 (.A0(net11),
    .A1(net996),
    .A2(net927),
    .A3(net1042),
    .S0(net968),
    .S1(net1021),
    .X(net16));
 sky130_fd_sc_hd__mux4_2 c145 (.A0(net952),
    .A1(net9),
    .A2(net1022),
    .A3(net735),
    .S0(net955),
    .S1(net930),
    .X(net17));
 sky130_fd_sc_hd__a41o_4 c146 (.A1(net924),
    .A2(net12),
    .A3(net930),
    .A4(net745),
    .B1(net1020),
    .X(net18));
 sky130_fd_sc_hd__a41o_4 c147 (.A1(net920),
    .A2(net15),
    .A3(net1020),
    .A4(net1042),
    .B1(net12),
    .X(net19));
 sky130_fd_sc_hd__a41o_4 c148 (.A1(net12),
    .A2(net924),
    .A3(net1020),
    .A4(net15),
    .B1(net920),
    .X(net871));
 sky130_fd_sc_hd__a41o_4 c149 (.A1(net19),
    .A2(net725),
    .A3(net925),
    .A4(net871),
    .B1(net920),
    .X(net20));
 sky130_fd_sc_hd__a41o_4 c150 (.A1(net915),
    .A2(net725),
    .A3(net1020),
    .A4(net871),
    .B1(net920),
    .X(net21));
 sky130_fd_sc_hd__mux4_2 c151 (.A0(net1085),
    .A1(net15),
    .A2(net924),
    .A3(net1020),
    .S0(net1016),
    .S1(net908),
    .X(net22));
 sky130_fd_sc_hd__mux4_2 c152 (.A0(net871),
    .A1(net1020),
    .A2(net905),
    .A3(net915),
    .S0(net6),
    .S1(net725),
    .X(net23));
 sky130_fd_sc_hd__mux4_2 c153 (.A0(net1023),
    .A1(net23),
    .A2(net12),
    .A3(net905),
    .S0(net19),
    .S1(net1018),
    .X(net24));
 sky130_fd_sc_hd__a41o_2 c154 (.A1(net996),
    .A2(net737),
    .A3(net1041),
    .A4(net952),
    .B1(net746),
    .X(net25));
 sky130_fd_sc_hd__a41o_4 c155 (.A1(net741),
    .A2(net755),
    .A3(net742),
    .A4(net12),
    .B1(net952),
    .X(net26));
 sky130_fd_sc_hd__a41o_1 c156 (.A1(net9),
    .A2(net970),
    .A3(net740),
    .A4(net26),
    .B1(net743),
    .X(net27));
 sky130_fd_sc_hd__a41o_4 c157 (.A1(net955),
    .A2(net929),
    .A3(net750),
    .A4(net743),
    .B1(net970),
    .X(net28));
 sky130_fd_sc_hd__a41o_4 c158 (.A1(net24),
    .A2(net759),
    .A3(net752),
    .A4(net929),
    .B1(net1041),
    .X(net29));
 sky130_fd_sc_hd__a41o_1 c159 (.A1(net923),
    .A2(net29),
    .A3(net929),
    .A4(net744),
    .B1(net954),
    .X(net843));
 sky130_fd_sc_hd__a41o_2 c160 (.A1(net902),
    .A2(net743),
    .A3(net1018),
    .A4(net23),
    .B1(net929),
    .X(net30));
 sky130_fd_sc_hd__mux4_2 c161 (.A0(net749),
    .A1(net24),
    .A2(net750),
    .A3(net29),
    .S0(net936),
    .S1(net1018),
    .X(net31));
 sky130_fd_sc_hd__a41o_2 c162 (.A1(net28),
    .A2(net747),
    .A3(net901),
    .A4(net972),
    .B1(net902),
    .X(net32));
 sky130_fd_sc_hd__mux4_2 c163 (.A0(net929),
    .A1(net902),
    .A2(net908),
    .A3(net1016),
    .S0(net757),
    .S1(net950),
    .X(net33));
 sky130_fd_sc_hd__a41o_1 c164 (.A1(net32),
    .A2(net751),
    .A3(net33),
    .A4(net903),
    .B1(net929),
    .X(net34));
 sky130_fd_sc_hd__a41o_4 c165 (.A1(net936),
    .A2(net9),
    .A3(net32),
    .A4(net24),
    .B1(net27),
    .X(net842));
 sky130_fd_sc_hd__mux4_2 c166 (.A0(net33),
    .A1(net28),
    .A2(net955),
    .A3(net971),
    .S0(net754),
    .S1(net743),
    .X(net35));
 sky130_fd_sc_hd__a41o_2 c167 (.A1(net896),
    .A2(net971),
    .A3(net32),
    .A4(net748),
    .B1(net29),
    .X(net881));
 sky130_fd_sc_hd__mux4_2 c168 (.A0(net881),
    .A1(net929),
    .A2(net970),
    .A3(net936),
    .S0(net757),
    .S1(net901),
    .X(net36));
 sky130_fd_sc_hd__mux4_2 c169 (.A0(net901),
    .A1(net747),
    .A2(net758),
    .A3(net898),
    .S0(net1023),
    .S1(net896),
    .X(net37));
 sky130_fd_sc_hd__mux4_2 c170 (.A0(net971),
    .A1(net881),
    .A2(net9),
    .A3(net1020),
    .S0(net37),
    .S1(net842),
    .X(net874));
 sky130_fd_sc_hd__mux4_2 c171 (.A0(net36),
    .A1(net29),
    .A2(net898),
    .A3(net1011),
    .S0(net1046),
    .S1(net896),
    .X(net38));
 sky130_fd_sc_hd__mux4_1 c172 (.A0(net1045),
    .A1(net38),
    .A2(net975),
    .A3(net903),
    .S0(net1076),
    .S1(net896),
    .X(net39));
 sky130_fd_sc_hd__mux4_1 c173 (.A0(net1075),
    .A1(net38),
    .A2(net929),
    .A3(net12),
    .S0(net1044),
    .S1(net624),
    .X(net40));
 sky130_fd_sc_hd__mux4_1 c174 (.A0(net26),
    .A1(net36),
    .A2(net38),
    .A3(net937),
    .S0(net881),
    .S1(net623),
    .X(net41));
 sky130_fd_sc_hd__mux4_1 c175 (.A0(net1071),
    .A1(net26),
    .A2(net38),
    .A3(net1075),
    .S1(net623),
    .X(net42));
 sky130_fd_sc_hd__a41o_2 c176 (.A1(net727),
    .A2(net747),
    .A3(net35),
    .A4(net26),
    .B1(net775),
    .X(net43));
 sky130_fd_sc_hd__mux4_2 c177 (.A0(net961),
    .A1(net762),
    .A2(net963),
    .A3(net782),
    .S0(net903),
    .S1(net19),
    .X(net44));
 sky130_fd_sc_hd__a41o_4 c178 (.A1(net950),
    .A2(net36),
    .A3(net747),
    .A4(net779),
    .B1(net555),
    .X(net45));
 sky130_fd_sc_hd__a41o_4 c179 (.A1(net770),
    .A2(net19),
    .A3(net765),
    .A4(net740),
    .B1(net908),
    .X(net46));
 sky130_fd_sc_hd__mux4_2 c180 (.A0(net46),
    .A1(net750),
    .A2(net757),
    .A3(net956),
    .S0(net727),
    .S1(net948),
    .X(net47));
 sky130_fd_sc_hd__mux4_1 c181 (.A0(net12),
    .A1(net8),
    .A2(net762),
    .A3(net961),
    .S0(net45),
    .S1(net1009),
    .X(net48));
 sky130_fd_sc_hd__mux4_2 c182 (.A0(net44),
    .A1(net753),
    .A2(net772),
    .A3(net904),
    .S0(net763),
    .S1(net770),
    .X(net49));
 sky130_fd_sc_hd__mux4_2 c183 (.A0(net1009),
    .A1(net1047),
    .A2(net904),
    .A3(net743),
    .S0(net771),
    .S1(net764),
    .X(net50));
 sky130_fd_sc_hd__mux4_1 c184 (.A0(net45),
    .A1(net771),
    .A2(net43),
    .A3(net782),
    .S0(net904),
    .S1(net50),
    .X(net51));
 sky130_fd_sc_hd__a41o_1 c185 (.A1(net781),
    .A2(net874),
    .A3(net775),
    .A4(net780),
    .B1(net49),
    .X(net52));
 sky130_fd_sc_hd__mux4_2 c186 (.A0(net743),
    .A1(net871),
    .A2(net776),
    .A3(net781),
    .S0(net761),
    .S1(net773),
    .X(net53));
 sky130_fd_sc_hd__mux4_2 c187 (.A0(net968),
    .A1(net781),
    .A2(net921),
    .A3(net771),
    .S0(net904),
    .S1(net952),
    .X(net54));
 sky130_fd_sc_hd__mux4_1 c188 (.A0(net1074),
    .A1(net32),
    .A2(net53),
    .A3(net26),
    .S0(net50),
    .S1(net944),
    .X(net55));
 sky130_fd_sc_hd__mux4_2 c189 (.A0(net782),
    .A1(net762),
    .A2(net932),
    .A3(net538),
    .S0(net559),
    .S1(net624),
    .X(net839));
 sky130_fd_sc_hd__mux4_2 c190 (.A0(net782),
    .A1(net776),
    .A2(net993),
    .A3(net770),
    .S0(net44),
    .S1(net625),
    .X(net56));
 sky130_fd_sc_hd__mux4_2 c191 (.A0(net747),
    .A1(net759),
    .A2(net772),
    .A3(net6),
    .S0(net56),
    .S1(net538),
    .X(net57));
 sky130_fd_sc_hd__mux4_1 c192 (.A0(net928),
    .A1(net749),
    .A2(net45),
    .A3(net57),
    .S0(net740),
    .S1(net757),
    .X(net58));
 sky130_fd_sc_hd__mux4_2 c193 (.A0(net54),
    .A1(net752),
    .A2(net53),
    .A3(net904),
    .S0(net776),
    .S1(net37),
    .X(net59));
 sky130_fd_sc_hd__mux4_2 c194 (.A0(net904),
    .A1(net59),
    .A2(net761),
    .A3(net56),
    .S0(net928),
    .S1(net881),
    .X(net60));
 sky130_fd_sc_hd__a41o_1 c195 (.A1(net53),
    .A2(net52),
    .A3(net57),
    .A4(net765),
    .B1(net59),
    .X(net61));
 sky130_fd_sc_hd__mux4_1 c196 (.A0(net50),
    .A1(net60),
    .A2(net59),
    .A3(net54),
    .S0(net1040),
    .S1(net626),
    .X(net62));
 sky130_fd_sc_hd__mux4_1 c197 (.A0(net60),
    .A1(net56),
    .A2(net59),
    .A3(net959),
    .S0(net537),
    .S1(net559),
    .X(net63));
 sky130_fd_sc_hd__mux4_2 c198 (.A0(net807),
    .A1(net874),
    .A2(net784),
    .A3(net737),
    .S0(net1070),
    .S1(net537),
    .X(net64));
 sky130_fd_sc_hd__mux4_2 c199 (.A0(net936),
    .A1(net786),
    .A2(net977),
    .A3(net763),
    .S0(net921),
    .S1(net625),
    .X(net858));
 sky130_fd_sc_hd__a41o_1 c200 (.A1(net793),
    .A2(net60),
    .A3(net804),
    .A4(net54),
    .B1(net744),
    .X(net65));
 sky130_fd_sc_hd__mux4_2 c201 (.A0(net784),
    .A1(net928),
    .A2(net56),
    .A3(net785),
    .S0(net790),
    .S1(net944),
    .X(net66));
 sky130_fd_sc_hd__a41o_2 c202 (.A1(net796),
    .A2(net776),
    .A3(net858),
    .A4(net43),
    .B1(net627),
    .X(net67));
 sky130_fd_sc_hd__mux4_2 c203 (.A0(net760),
    .A1(net796),
    .A2(net769),
    .A3(net908),
    .S0(net871),
    .S1(net543),
    .X(net68));
 sky130_fd_sc_hd__a41o_2 c204 (.A1(net67),
    .A2(net858),
    .A3(net784),
    .A4(net874),
    .B1(net764),
    .X(net69));
 sky130_fd_sc_hd__mux4_2 c205 (.A0(net987),
    .A1(net752),
    .A2(net751),
    .A3(net749),
    .S0(net902),
    .S1(net943),
    .X(net70));
 sky130_fd_sc_hd__mux4_2 c206 (.A0(net786),
    .A1(net775),
    .A2(net771),
    .A3(net798),
    .S0(net944),
    .S1(net628),
    .X(net71));
 sky130_fd_sc_hd__mux4_1 c207 (.A0(net956),
    .A1(net64),
    .A2(net958),
    .A3(net1016),
    .S0(net60),
    .S1(net997),
    .X(net72));
 sky130_fd_sc_hd__mux4_1 c208 (.A0(net69),
    .A1(net727),
    .A2(net1015),
    .A3(net793),
    .S0(net807),
    .S1(net71),
    .X(net73));
 sky130_fd_sc_hd__mux4_1 c209 (.A0(net66),
    .A1(net842),
    .A2(net52),
    .A3(net952),
    .S0(net629),
    .S1(clknet_1_0__leaf_net630),
    .X(net74));
 sky130_fd_sc_hd__mux4_2 c210 (.A0(net763),
    .A1(net788),
    .A2(net881),
    .A3(net972),
    .S0(net970),
    .S1(net880),
    .X(net75));
 sky130_fd_sc_hd__a41o_1 c211 (.A1(net52),
    .A2(net68),
    .A3(net70),
    .A4(net961),
    .B1(net75),
    .X(net76));
 sky130_fd_sc_hd__mux4_1 c212 (.A0(net798),
    .A1(net958),
    .A2(net52),
    .A3(net727),
    .S0(net970),
    .S1(net880),
    .X(net77));
 sky130_fd_sc_hd__a41o_2 c213 (.A1(net70),
    .A2(net842),
    .A3(net738),
    .A4(net746),
    .B1(net802),
    .X(net849));
 sky130_fd_sc_hd__mux4_1 c214 (.A0(net937),
    .A1(net958),
    .A2(net997),
    .A3(net67),
    .S0(clknet_1_1__leaf_net868),
    .S1(clknet_1_0__leaf_net630),
    .X(net78));
 sky130_fd_sc_hd__mux4_2 c215 (.A0(net71),
    .A1(net849),
    .A2(net748),
    .A3(net796),
    .S0(net974),
    .S1(net795),
    .X(net79));
 sky130_fd_sc_hd__mux4_1 c216 (.A0(net68),
    .A1(net849),
    .A2(net801),
    .A3(clknet_1_0__leaf_net78),
    .S0(clknet_1_1__leaf_net868),
    .S1(net629),
    .X(net80));
 sky130_fd_sc_hd__mux4_1 c217 (.A0(net79),
    .A1(net68),
    .A2(net801),
    .A3(net881),
    .S0(net623),
    .S1(clknet_1_0__leaf_net630),
    .X(net844));
 sky130_fd_sc_hd__mux4_1 c218 (.A0(net1016),
    .A1(clknet_1_0__leaf_net78),
    .A2(net70),
    .A3(net943),
    .S0(net880),
    .S1(clknet_1_1__leaf_net631),
    .X(net81));
 sky130_fd_sc_hd__mux4_1 c219 (.A0(net64),
    .A1(net904),
    .A2(net798),
    .A3(net880),
    .S0(net605),
    .S1(clknet_1_1__leaf_net631),
    .X(net82));
 sky130_fd_sc_hd__mux4_1 c220 (.A0(net879),
    .A1(net60),
    .A2(net876),
    .A3(net794),
    .S0(net943),
    .S1(net625),
    .X(net83));
 sky130_fd_sc_hd__mux4_1 c221 (.A0(net4),
    .A1(net849),
    .A2(net808),
    .A3(net555),
    .S0(net943),
    .S1(clknet_1_0__leaf_net631),
    .X(net84));
 sky130_fd_sc_hd__mux4_2 c222 (.A0(net810),
    .A1(net902),
    .A2(net879),
    .A3(net761),
    .S0(net43),
    .S1(net873),
    .X(net859));
 sky130_fd_sc_hd__mux4_1 c223 (.A0(net4),
    .A1(net0),
    .A2(net902),
    .A3(net738),
    .S0(net761),
    .S1(net627),
    .X(net85));
 sky130_fd_sc_hd__mux4_1 c224 (.A0(net816),
    .A1(net859),
    .A2(clknet_1_0__leaf_net84),
    .A3(net85),
    .S0(net963),
    .S1(net943),
    .X(net86));
 sky130_fd_sc_hd__mux4_2 c225 (.A0(net727),
    .A1(net1023),
    .A2(net997),
    .A3(net1013),
    .S0(net943),
    .S1(net880),
    .X(net87));
 sky130_fd_sc_hd__mux4_2 c226 (.A0(net812),
    .A1(net816),
    .A2(net0),
    .A3(net928),
    .S0(net625),
    .S1(net627),
    .X(net88));
 sky130_fd_sc_hd__mux4_2 c227 (.A0(net0),
    .A1(net740),
    .A2(net974),
    .A3(net1013),
    .S0(net743),
    .S1(net928),
    .X(net89));
 sky130_fd_sc_hd__mux4_1 c228 (.A0(net775),
    .A1(net60),
    .A2(net1016),
    .A3(net760),
    .S0(net70),
    .S1(net89),
    .X(net90));
 sky130_fd_sc_hd__mux4_1 c229 (.A0(net88),
    .A1(net89),
    .A2(net810),
    .A3(net1017),
    .S0(clknet_1_0__leaf_net86),
    .S1(net943),
    .X(net91));
 sky130_fd_sc_hd__mux4_2 c230 (.A0(net974),
    .A1(net752),
    .A2(net958),
    .A3(net871),
    .S0(net867),
    .S1(net943),
    .X(net92));
 sky130_fd_sc_hd__mux4_1 c231 (.A0(net754),
    .A1(clknet_1_0__leaf_net84),
    .A2(net804),
    .A3(net816),
    .S0(net873),
    .S1(net627),
    .X(net834));
 sky130_fd_sc_hd__mux4_1 c232 (.A0(net904),
    .A1(net92),
    .A2(net957),
    .A3(net867),
    .S0(net943),
    .S1(clknet_1_0__leaf_net632),
    .X(net93));
 sky130_fd_sc_hd__mux4_1 c233 (.A0(net85),
    .A1(clknet_1_0__leaf_net834),
    .A2(net89),
    .A3(clknet_1_0__leaf_net86),
    .S0(net958),
    .S1(net88),
    .X(net94));
 sky130_fd_sc_hd__mux4_1 c234 (.A0(net89),
    .A1(net997),
    .A2(clknet_1_0__leaf_net84),
    .A3(net749),
    .S0(net543),
    .S1(clknet_1_0__leaf_net631),
    .X(net875));
 sky130_fd_sc_hd__mux4_1 c235 (.A0(clknet_1_1__leaf_net93),
    .A1(net979),
    .A2(net3),
    .A3(net737),
    .S0(clknet_1_0__leaf_net834),
    .S1(net943),
    .X(net95));
 sky130_fd_sc_hd__mux4_1 c236 (.A0(net785),
    .A1(net859),
    .A2(net624),
    .A3(clknet_1_0__leaf_net631),
    .S0(clknet_1_0__leaf_net632),
    .S1(net634),
    .X(net96));
 sky130_fd_sc_hd__mux4_1 c237 (.A0(net43),
    .A1(clknet_1_1__leaf_net875),
    .A2(net871),
    .A3(net3),
    .S0(net849),
    .S1(net633),
    .X(net97));
 sky130_fd_sc_hd__mux4_1 c238 (.A0(clknet_1_1__leaf_net86),
    .A1(net88),
    .A2(net75),
    .A3(clknet_1_0__leaf_net93),
    .S0(net794),
    .S1(clknet_1_0__leaf_net868),
    .X(net98));
 sky130_fd_sc_hd__mux4_1 c239 (.A0(net795),
    .A1(net89),
    .A2(clknet_1_0__leaf_net875),
    .A3(clknet_1_0__leaf_net96),
    .S0(net634),
    .S1(net635),
    .X(net99));
 sky130_fd_sc_hd__mux4_1 c240 (.A0(clknet_1_1__leaf_net96),
    .A1(net88),
    .A2(net43),
    .A3(net867),
    .S0(clknet_1_0__leaf_net851),
    .S1(net628),
    .X(net100));
 sky130_fd_sc_hd__mux4_1 c241 (.A0(clknet_1_1__leaf_net86),
    .A1(net43),
    .A2(net85),
    .S0(net629),
    .S1(net635),
    .X(net851));
 sky130_fd_sc_hd__a41o_2 c264 (.A1(net924),
    .A2(net948),
    .A3(net965),
    .A4(net1041),
    .B1(net11),
    .X(net102));
 sky130_fd_sc_hd__a41o_1 c265 (.A1(net966),
    .A2(net725),
    .A3(net7),
    .A4(net1022),
    .B1(net954),
    .X(net103));
 sky130_fd_sc_hd__a41o_1 c266 (.A1(net724),
    .A2(net1042),
    .A3(net975),
    .A4(net9),
    .B1(net920),
    .X(net862));
 sky130_fd_sc_hd__a41o_2 c267 (.A1(net745),
    .A2(net918),
    .A3(net923),
    .A4(net724),
    .B1(net966),
    .X(net104));
 sky130_fd_sc_hd__mux4_2 c268 (.A0(net916),
    .A1(net9),
    .A2(net934),
    .A3(net959),
    .S0(net954),
    .S1(net1021),
    .X(net105));
 sky130_fd_sc_hd__a41o_2 c269 (.A1(net11),
    .A2(net1042),
    .A3(net934),
    .A4(net916),
    .B1(net914),
    .X(net106));
 sky130_fd_sc_hd__mux4_1 c270 (.A0(net15),
    .A1(net102),
    .A2(net916),
    .A3(net964),
    .S0(net966),
    .S1(net954),
    .X(net107));
 sky130_fd_sc_hd__a41o_4 c271 (.A1(net1022),
    .A2(net910),
    .A3(net724),
    .A4(net914),
    .B1(net917),
    .X(net108));
 sky130_fd_sc_hd__a41o_4 c272 (.A1(net108),
    .A2(net23),
    .A3(net934),
    .A4(net910),
    .B1(net916),
    .X(net109));
 sky130_fd_sc_hd__a41o_2 c273 (.A1(net109),
    .A2(net914),
    .A3(net916),
    .A4(net910),
    .B1(net1042),
    .X(net110));
 sky130_fd_sc_hd__a41o_2 c274 (.A1(net934),
    .A2(net914),
    .A3(net910),
    .A4(net917),
    .B1(net977),
    .X(net111));
 sky130_fd_sc_hd__a41o_2 c275 (.A1(net110),
    .A2(net905),
    .A3(net919),
    .A4(net923),
    .B1(net911),
    .X(net841));
 sky130_fd_sc_hd__a41o_4 c276 (.A1(net934),
    .A2(net110),
    .A3(net111),
    .A4(net910),
    .B1(net916),
    .X(net112));
 sky130_fd_sc_hd__mux4_2 c277 (.A0(net911),
    .A1(net111),
    .A2(net899),
    .A3(net916),
    .S0(net1022),
    .S1(net110),
    .X(net113));
 sky130_fd_sc_hd__mux4_2 c278 (.A0(net971),
    .A1(net899),
    .A2(net113),
    .A3(net9),
    .S0(net111),
    .S1(net910),
    .X(net833));
 sky130_fd_sc_hd__mux4_2 c279 (.A0(net113),
    .A1(net899),
    .A2(net959),
    .A3(net111),
    .S0(net910),
    .S1(net917),
    .X(net114));
 sky130_fd_sc_hd__mux4_2 c280 (.A0(net102),
    .A1(net113),
    .A2(net110),
    .A3(net899),
    .S0(net910),
    .S1(net916),
    .X(net852));
 sky130_fd_sc_hd__mux4_2 c281 (.A0(net106),
    .A1(net914),
    .A2(net111),
    .A3(net917),
    .S0(net964),
    .S1(net852),
    .X(net115));
 sky130_fd_sc_hd__mux4_2 c282 (.A0(net852),
    .A1(net115),
    .A2(net106),
    .A3(net113),
    .S0(net899),
    .S1(net917),
    .X(net116));
 sky130_fd_sc_hd__mux4_2 c283 (.A0(net15),
    .A1(net852),
    .A2(net116),
    .A3(net923),
    .S0(net115),
    .S1(net899),
    .X(net117));
 sky130_fd_sc_hd__mux4_2 c284 (.A0(net116),
    .A1(net833),
    .A2(net1053),
    .A3(net108),
    .S0(net104),
    .S1(net899),
    .X(net118));
 sky130_fd_sc_hd__mux4_1 c285 (.A0(net111),
    .A1(net118),
    .A2(net899),
    .A3(net910),
    .S0(net105),
    .S1(net895),
    .X(net119));
 sky130_fd_sc_hd__a41o_2 c286 (.A1(net751),
    .A2(net970),
    .A3(net735),
    .A4(net28),
    .B1(net555),
    .X(net120));
 sky130_fd_sc_hd__a41o_2 c287 (.A1(net746),
    .A2(net106),
    .A3(net924),
    .A4(net28),
    .B1(net749),
    .X(net121));
 sky130_fd_sc_hd__a41o_4 c288 (.A1(net121),
    .A2(net105),
    .A3(net923),
    .A4(net950),
    .B1(net1021),
    .X(net122));
 sky130_fd_sc_hd__a41o_2 c289 (.A1(net740),
    .A2(net121),
    .A3(net965),
    .A4(net911),
    .B1(net725),
    .X(net123));
 sky130_fd_sc_hd__mux4_2 c290 (.A0(net113),
    .A1(net923),
    .A2(net738),
    .A3(net122),
    .S0(net748),
    .S1(net921),
    .X(net124));
 sky130_fd_sc_hd__a41o_2 c291 (.A1(net1021),
    .A2(net929),
    .A3(net896),
    .A4(net121),
    .B1(net555),
    .X(net125));
 sky130_fd_sc_hd__a41o_2 c292 (.A1(net29),
    .A2(net956),
    .A3(net110),
    .A4(net122),
    .B1(net555),
    .X(net864));
 sky130_fd_sc_hd__a41o_2 c293 (.A1(net122),
    .A2(net841),
    .A3(net1018),
    .A4(net725),
    .B1(net749),
    .X(net126));
 sky130_fd_sc_hd__a41o_4 c294 (.A1(net26),
    .A2(net916),
    .A3(net896),
    .A4(net990),
    .B1(net944),
    .X(net127));
 sky130_fd_sc_hd__mux4_2 c295 (.A0(net124),
    .A1(net109),
    .A2(net125),
    .A3(net898),
    .S0(net741),
    .S1(net991),
    .X(net128));
 sky130_fd_sc_hd__a41o_2 c296 (.A1(net127),
    .A2(net897),
    .A3(net975),
    .A4(net1020),
    .B1(net916),
    .X(net129));
 sky130_fd_sc_hd__a41o_2 c297 (.A1(net125),
    .A2(net124),
    .A3(net29),
    .A4(net898),
    .B1(net965),
    .X(net826));
 sky130_fd_sc_hd__mux4_2 c298 (.A0(net120),
    .A1(net758),
    .A2(net127),
    .A3(net121),
    .S0(net892),
    .S1(net129),
    .X(net130));
 sky130_fd_sc_hd__a41o_1 c299 (.A1(net892),
    .A2(net130),
    .A3(net1009),
    .A4(net897),
    .B1(net993),
    .X(net131));
 sky130_fd_sc_hd__mux4_2 c300 (.A0(net123),
    .A1(net892),
    .A2(net897),
    .A3(net970),
    .S0(net945),
    .S1(net555),
    .X(net132));
 sky130_fd_sc_hd__mux4_2 c301 (.A0(net961),
    .A1(net748),
    .A2(net26),
    .A3(net892),
    .S0(net125),
    .S1(net945),
    .X(net133));
 sky130_fd_sc_hd__a41o_1 c302 (.A1(net897),
    .A2(net130),
    .A3(net892),
    .A4(net133),
    .B1(net128),
    .X(net134));
 sky130_fd_sc_hd__mux4_1 c303 (.A0(net133),
    .A1(net896),
    .A2(net123),
    .A3(net128),
    .S0(net892),
    .S1(net130),
    .X(net135));
 sky130_fd_sc_hd__mux4_1 c304 (.A0(net127),
    .A1(net29),
    .A2(net892),
    .A3(net38),
    .S0(net132),
    .S1(net942),
    .X(net136));
 sky130_fd_sc_hd__mux4_1 c305 (.A0(net992),
    .A1(net133),
    .A2(net129),
    .A3(net893),
    .S0(net942),
    .S1(net940),
    .X(net137));
 sky130_fd_sc_hd__mux4_1 c306 (.A0(net864),
    .A1(net746),
    .A2(net133),
    .A3(net129),
    .S0(net945),
    .S1(net942),
    .X(net138));
 sky130_fd_sc_hd__mux4_1 c307 (.A0(net864),
    .A1(net125),
    .A2(net102),
    .A3(net132),
    .S0(net945),
    .S1(net940),
    .X(net139));
 sky130_fd_sc_hd__mux4_1 c308 (.A0(net132),
    .A1(net913),
    .A2(net993),
    .A3(net965),
    .S0(net538),
    .S1(net1024),
    .X(net140));
 sky130_fd_sc_hd__mux4_1 c309 (.A0(net125),
    .A1(net737),
    .A2(net54),
    .A3(net49),
    .S0(net977),
    .S1(net921),
    .X(net141));
 sky130_fd_sc_hd__mux4_2 c310 (.A0(net769),
    .A1(net129),
    .A2(net759),
    .A3(net750),
    .S0(net26),
    .S1(net627),
    .X(net846));
 sky130_fd_sc_hd__mux4_1 c311 (.A0(net929),
    .A1(net744),
    .A2(net45),
    .A3(net952),
    .S0(net102),
    .S1(net628),
    .X(net142));
 sky130_fd_sc_hd__mux4_2 c312 (.A0(net779),
    .A1(net120),
    .A2(net915),
    .A3(net963),
    .S0(net942),
    .S1(net641),
    .X(net143));
 sky130_fd_sc_hd__mux4_1 c313 (.A0(net111),
    .A1(net26),
    .A2(net132),
    .A3(net753),
    .S0(net934),
    .S1(net977),
    .X(net144));
 sky130_fd_sc_hd__mux4_2 c314 (.A0(net141),
    .A1(net914),
    .A2(net773),
    .A3(net892),
    .S0(net46),
    .S1(net527),
    .X(net145));
 sky130_fd_sc_hd__mux4_2 c315 (.A0(net44),
    .A1(net931),
    .A2(net903),
    .A3(net914),
    .S0(net56),
    .S1(net141),
    .X(net146));
 sky130_fd_sc_hd__mux4_1 c316 (.A0(net146),
    .A1(net771),
    .A2(net913),
    .A3(net935),
    .S0(net750),
    .S1(net46),
    .X(net147));
 sky130_fd_sc_hd__mux4_1 c317 (.A0(net45),
    .A1(net127),
    .A2(net59),
    .A3(net122),
    .S0(net53),
    .S1(net919),
    .X(net148));
 sky130_fd_sc_hd__mux4_1 c318 (.A0(net102),
    .A1(net132),
    .A2(net111),
    .A3(net740),
    .S0(net127),
    .S1(net737),
    .X(net149));
 sky130_fd_sc_hd__mux4_1 c319 (.A0(net914),
    .A1(net122),
    .A2(net127),
    .A3(net527),
    .S0(net944),
    .S1(net645),
    .X(net150));
 sky130_fd_sc_hd__mux4_1 c320 (.A0(net145),
    .A1(net45),
    .A2(net1011),
    .A3(net742),
    .S0(net890),
    .S1(net643),
    .X(net151));
 sky130_fd_sc_hd__mux4_1 c321 (.A0(net32),
    .A1(net931),
    .A2(net890),
    .A3(net130),
    .S0(net897),
    .S1(net643),
    .X(net152));
 sky130_fd_sc_hd__mux4_2 c322 (.A0(net773),
    .A1(net890),
    .A2(net124),
    .A3(net748),
    .S0(net638),
    .S1(net646),
    .X(net153));
 sky130_fd_sc_hd__mux4_1 c323 (.A0(net26),
    .A1(net145),
    .A2(net153),
    .A3(net44),
    .S0(net644),
    .S1(net646),
    .X(net154));
 sky130_fd_sc_hd__a41o_1 c324 (.A1(net970),
    .A2(net779),
    .A3(clknet_1_1__leaf_net571),
    .A4(net865),
    .B1(net646),
    .X(net155));
 sky130_fd_sc_hd__mux4_2 c325 (.A0(net751),
    .A1(net890),
    .A2(net974),
    .A3(net538),
    .S0(net551),
    .S1(net646),
    .X(net156));
 sky130_fd_sc_hd__mux4_1 c326 (.A0(net890),
    .A1(net153),
    .A2(net750),
    .A3(net32),
    .S0(net156),
    .S1(net865),
    .X(net157));
 sky130_fd_sc_hd__mux4_1 c327 (.A0(net156),
    .A1(net146),
    .A2(net890),
    .A3(net779),
    .S0(clknet_1_0__leaf_net155),
    .S1(net865),
    .X(net158));
 sky130_fd_sc_hd__mux4_1 c328 (.A0(net49),
    .A1(net846),
    .A2(clknet_1_0__leaf_net155),
    .A3(net156),
    .S0(net645),
    .S1(net648),
    .X(net159));
 sky130_fd_sc_hd__mux4_1 c329 (.A0(net153),
    .A1(net891),
    .A2(net141),
    .A3(net551),
    .S0(net865),
    .S1(net649),
    .X(net160));
 sky130_fd_sc_hd__mux4_1 c330 (.A0(clknet_1_1__leaf_net78),
    .A1(net70),
    .A2(net75),
    .A3(net744),
    .S0(net890),
    .S1(net67),
    .X(net161));
 sky130_fd_sc_hd__mux4_1 c331 (.A0(net36),
    .A1(net788),
    .A2(net75),
    .A3(net955),
    .S0(net948),
    .S1(net890),
    .X(net162));
 sky130_fd_sc_hd__mux4_2 c332 (.A0(net790),
    .A1(net776),
    .A2(net901),
    .A3(net71),
    .S0(net555),
    .S1(net641),
    .X(net163));
 sky130_fd_sc_hd__mux4_2 c333 (.A0(net121),
    .A1(net790),
    .A2(net761),
    .A3(net902),
    .S0(net163),
    .S1(net963),
    .X(net164));
 sky130_fd_sc_hd__mux4_1 c334 (.A0(net130),
    .A1(net71),
    .A2(net64),
    .A3(net936),
    .S0(net1036),
    .S1(net1030),
    .X(net165));
 sky130_fd_sc_hd__mux4_1 c335 (.A0(net162),
    .A1(net738),
    .A2(net1017),
    .A3(net1015),
    .S0(net998),
    .S1(net641),
    .X(net166));
 sky130_fd_sc_hd__mux4_1 c336 (.A0(net64),
    .A1(net60),
    .A2(net936),
    .A3(net904),
    .S0(net914),
    .S1(net940),
    .X(net167));
 sky130_fd_sc_hd__mux4_2 c337 (.A0(net54),
    .A1(net1041),
    .A2(net143),
    .A3(net586),
    .S0(net643),
    .S1(net650),
    .X(net828));
 sky130_fd_sc_hd__mux4_1 c338 (.A0(net841),
    .A1(net898),
    .A2(net892),
    .A3(net968),
    .S0(net538),
    .S1(net585),
    .X(net168));
 sky130_fd_sc_hd__mux4_1 c339 (.A0(net164),
    .A1(net162),
    .A2(clknet_1_1__leaf_net844),
    .A3(net740),
    .S0(net1023),
    .S1(net585),
    .X(net169));
 sky130_fd_sc_hd__mux4_2 c340 (.A0(net163),
    .A1(net805),
    .A2(net828),
    .A3(net164),
    .S0(net754),
    .S1(net890),
    .X(net170));
 sky130_fd_sc_hd__mux4_2 c341 (.A0(net1041),
    .A1(net801),
    .A2(net143),
    .A3(net952),
    .S0(net942),
    .S1(net623),
    .X(net832));
 sky130_fd_sc_hd__mux4_1 c342 (.A0(net771),
    .A1(net168),
    .A2(net143),
    .A3(net902),
    .S0(net623),
    .S1(net650),
    .X(net171));
 sky130_fd_sc_hd__mux4_1 c343 (.A0(net66),
    .A1(net832),
    .A2(net979),
    .A3(net898),
    .S0(net629),
    .S1(clknet_1_1__leaf_net651),
    .X(net855));
 sky130_fd_sc_hd__mux4_1 c344 (.A0(net50),
    .A1(net168),
    .A2(net120),
    .A3(net890),
    .S0(net801),
    .S1(clknet_1_1__leaf_net651),
    .X(net172));
 sky130_fd_sc_hd__mux4_1 c345 (.A0(net832),
    .A1(net543),
    .A2(clknet_1_1__leaf_net571),
    .A3(net835),
    .S0(net650),
    .S1(clknet_1_1__leaf_net651),
    .X(net173));
 sky130_fd_sc_hd__mux4_1 c346 (.A0(net164),
    .A1(clknet_1_0__leaf_net173),
    .A2(net771),
    .A3(net585),
    .S0(net650),
    .S1(clknet_1_1__leaf_net651),
    .X(net174));
 sky130_fd_sc_hd__mux4_1 c347 (.A0(net170),
    .A1(net780),
    .A2(clknet_1_0__leaf_net174),
    .A3(net543),
    .S0(net641),
    .S1(clknet_1_1__leaf_net651),
    .X(net175));
 sky130_fd_sc_hd__mux4_1 c348 (.A0(clknet_1_0__leaf_net173),
    .A1(clknet_1_0__leaf_net174),
    .A2(net835),
    .A3(net625),
    .S0(net650),
    .S1(clknet_1_0__leaf_net651),
    .X(net836));
 sky130_fd_sc_hd__mux4_1 c349 (.A0(net828),
    .A1(clknet_1_0__leaf_net173),
    .A2(net143),
    .A3(net835),
    .S0(net650),
    .S1(clknet_1_0__leaf_net651),
    .X(net176));
 sky130_fd_sc_hd__mux4_1 c350 (.A0(clknet_1_1__leaf_net173),
    .A1(clknet_1_0__leaf_net174),
    .A2(net828),
    .A3(net864),
    .S0(net835),
    .S1(clknet_1_0__leaf_net651),
    .X(net177));
 sky130_fd_sc_hd__mux4_1 c351 (.A0(net117),
    .A1(clknet_1_0__leaf_net177),
    .A2(clknet_1_0__leaf_net174),
    .A3(net68),
    .S0(clknet_1_1__leaf_net173),
    .S1(net835),
    .X(net178));
 sky130_fd_sc_hd__mux4_1 c352 (.A0(clknet_1_1__leaf_net844),
    .A1(net3),
    .A2(net873),
    .A3(net628),
    .S0(net634),
    .S1(clknet_1_0__leaf_net652),
    .X(net179));
 sky130_fd_sc_hd__mux4_1 c353 (.A0(net1008),
    .A1(net928),
    .A2(clknet_1_0__leaf_net855),
    .A3(net555),
    .S0(net628),
    .S1(net633),
    .X(net861));
 sky130_fd_sc_hd__mux4_1 c354 (.A0(net1023),
    .A1(clknet_1_1__leaf_net84),
    .A2(net3),
    .A3(net962),
    .S0(net1),
    .S1(clknet_1_0__leaf_net571),
    .X(net180));
 sky130_fd_sc_hd__mux4_1 c355 (.A0(net958),
    .A1(net75),
    .A2(net802),
    .A3(net817),
    .S0(net757),
    .S1(clknet_1_0__leaf_net571),
    .X(net857));
 sky130_fd_sc_hd__mux4_1 c356 (.A0(net156),
    .A1(clknet_1_0__leaf_net173),
    .A2(net1),
    .A3(net68),
    .S0(net555),
    .S1(net643),
    .X(net181));
 sky130_fd_sc_hd__mux4_2 c357 (.A0(net817),
    .A1(net937),
    .A2(net128),
    .A3(net88),
    .S0(net627),
    .S1(net643),
    .X(net182));
 sky130_fd_sc_hd__mux4_1 c358 (.A0(net749),
    .A1(net128),
    .A2(clknet_1_1__leaf_net84),
    .A3(net864),
    .S0(net590),
    .S1(net627),
    .X(net183));
 sky130_fd_sc_hd__mux4_1 c359 (.A0(net802),
    .A1(net863),
    .A2(net864),
    .A3(clknet_1_0__leaf_net834),
    .S0(net636),
    .S1(clknet_1_0__leaf_net651),
    .X(net184));
 sky130_fd_sc_hd__mux4_1 c360 (.A0(net802),
    .A1(net87),
    .A2(clknet_1_1__leaf_net183),
    .A3(net552),
    .S0(net873),
    .S1(net606),
    .X(net185));
 sky130_fd_sc_hd__mux4_1 c361 (.A0(net1008),
    .A1(net70),
    .A2(net780),
    .A3(net958),
    .S0(net590),
    .S1(clknet_1_0__leaf_net652),
    .X(net866));
 sky130_fd_sc_hd__mux4_1 c362 (.A0(net818),
    .A1(net813),
    .A2(clknet_1_0__leaf_net177),
    .A3(clknet_1_1__leaf_net866),
    .S0(clknet_1_0__leaf_net868),
    .S1(net606),
    .X(net186));
 sky130_fd_sc_hd__mux4_1 c363 (.A0(net738),
    .A1(net852),
    .A2(net813),
    .A3(clknet_1_1__leaf_net84),
    .S0(net590),
    .S1(net629),
    .X(net850));
 sky130_fd_sc_hd__mux4_1 c364 (.A0(clknet_1_1__leaf_net866),
    .A1(net858),
    .A2(net846),
    .A3(clknet_1_0__leaf_net177),
    .S0(clknet_1_1__leaf_net571),
    .S1(clknet_1_1__leaf_net868),
    .X(net187));
 sky130_fd_sc_hd__mux4_1 c365 (.A0(clknet_1_1__leaf_net180),
    .A1(net815),
    .A2(net122),
    .A3(net859),
    .S0(clknet_1_0__leaf_net183),
    .S1(net636),
    .X(net188));
 sky130_fd_sc_hd__mux4_1 c366 (.A0(clknet_1_1__leaf_net855),
    .A1(net746),
    .A2(net1011),
    .A3(clknet_1_1__leaf_net851),
    .S0(clknet_1_0__leaf_net571),
    .S1(net590),
    .X(net189));
 sky130_fd_sc_hd__mux4_1 c367 (.A0(clknet_1_1__leaf_net84),
    .A1(clknet_1_1__leaf_net189),
    .A2(net928),
    .A3(net904),
    .S0(net979),
    .S1(net650),
    .X(net190));
 sky130_fd_sc_hd__mux4_1 c368 (.A0(net914),
    .A1(net957),
    .A2(net771),
    .A3(net813),
    .S0(net552),
    .S1(net606),
    .X(net856));
 sky130_fd_sc_hd__mux4_1 c369 (.A0(clknet_1_0__leaf_net844),
    .A1(net833),
    .A2(net842),
    .A3(net1),
    .S0(clknet_1_0__leaf_net180),
    .S1(net873),
    .X(net191));
 sky130_fd_sc_hd__mux4_1 c370 (.A0(clknet_1_0__leaf_net183),
    .A1(net87),
    .A2(net849),
    .S0(net628),
    .S1(clknet_1_0__leaf_net651),
    .X(net853));
 sky130_fd_sc_hd__mux4_1 c371 (.A0(net856),
    .A1(net128),
    .A2(clknet_1_0__leaf_net866),
    .A3(net758),
    .S0(net552),
    .S1(net590),
    .X(net860));
 sky130_fd_sc_hd__mux4_1 c372 (.A0(net186),
    .A1(clknet_1_1__leaf_net189),
    .A2(net821),
    .A3(net902),
    .S0(net828),
    .S1(net543),
    .X(net193));
 sky130_fd_sc_hd__mux4_1 c373 (.A0(net813),
    .A1(clknet_1_0__leaf_net860),
    .A2(net814),
    .A3(clknet_1_0__leaf_net189),
    .S0(net579),
    .S1(net636),
    .X(net194));
 sky130_fd_sc_hd__a41o_4 c396 (.A1(net735),
    .A2(net833),
    .A3(net953),
    .A4(net115),
    .B1(net637),
    .X(net195));
 sky130_fd_sc_hd__a41o_2 c397 (.A1(net931),
    .A2(net934),
    .A3(net115),
    .A4(net972),
    .B1(net195),
    .X(net196));
 sky130_fd_sc_hd__mux4_2 c398 (.A0(net980),
    .A1(net735),
    .A2(net955),
    .A3(net918),
    .S0(net1041),
    .S1(net1010),
    .X(net197));
 sky130_fd_sc_hd__a41o_2 c399 (.A1(net1023),
    .A2(net915),
    .A3(net996),
    .A4(net1022),
    .B1(net934),
    .X(net198));
 sky130_fd_sc_hd__sdfbbn_1 c400 (.CLK_N(clknet_4_14_0_clk),
    .D(net195),
    .RESET_B(net745),
    .SCD(net118),
    .SCE(net933),
    .SET_B(net198),
    .Q(net200),
    .Q_N(net199));
 sky130_fd_sc_hd__a41o_2 c401 (.A1(net725),
    .A2(net906),
    .A3(net899),
    .A4(net946),
    .B1(net951),
    .X(net201));
 sky130_fd_sc_hd__a41o_1 c402 (.A1(net201),
    .A2(net115),
    .A3(net947),
    .A4(net195),
    .B1(net906),
    .X(net202));
 sky130_fd_sc_hd__a41o_2 c403 (.A1(net955),
    .A2(net745),
    .A3(net947),
    .A4(net906),
    .B1(net201),
    .X(net203));
 sky130_fd_sc_hd__mux4_1 c404 (.A0(net202),
    .A1(net906),
    .A2(net946),
    .A3(net203),
    .S0(net911),
    .S1(net637),
    .X(net204));
 sky130_fd_sc_hd__mux4_2 c405 (.A0(net947),
    .A1(net735),
    .A2(net927),
    .A3(net971),
    .S0(net203),
    .S1(net906),
    .X(net205));
 sky130_fd_sc_hd__mux4_1 c406 (.A0(net197),
    .A1(net203),
    .A2(net946),
    .A3(net196),
    .S0(net894),
    .S1(net906),
    .X(net206));
 sky130_fd_sc_hd__mux4_1 c407 (.A0(net203),
    .A1(net202),
    .A2(net955),
    .A3(net910),
    .S0(net899),
    .S1(net544),
    .X(net207));
 sky130_fd_sc_hd__mux4_2 c408 (.A0(net971),
    .A1(net996),
    .A2(net203),
    .A3(net921),
    .S0(net1022),
    .S1(net657),
    .X(net208));
 sky130_fd_sc_hd__mux4_2 c409 (.A0(net197),
    .A1(net894),
    .A2(net203),
    .A3(net544),
    .S0(net654),
    .S1(net656),
    .X(net209));
 sky130_fd_sc_hd__mux4_1 c410 (.A0(net209),
    .A1(net918),
    .A2(net947),
    .A3(net115),
    .S0(net202),
    .S1(net894),
    .X(net210));
 sky130_fd_sc_hd__mux4_2 c411 (.A0(net208),
    .A1(net918),
    .A2(net833),
    .A3(net946),
    .S0(net544),
    .S1(net654),
    .X(net211));
 sky130_fd_sc_hd__mux4_2 c412 (.A0(net104),
    .A1(net906),
    .A2(net946),
    .A3(net654),
    .S0(net656),
    .S1(net659),
    .X(net212));
 sky130_fd_sc_hd__mux4_2 c413 (.A0(net725),
    .A1(net208),
    .A2(net894),
    .A3(net906),
    .S0(net654),
    .S1(net658),
    .X(net213));
 sky130_fd_sc_hd__mux4_2 c414 (.A0(net203),
    .A1(net1009),
    .A2(net212),
    .A3(net894),
    .S0(net655),
    .S1(net659),
    .X(net214));
 sky130_fd_sc_hd__mux4_2 c415 (.A0(net214),
    .A1(net213),
    .A2(net211),
    .A3(net203),
    .S0(net947),
    .S1(net209),
    .X(net215));
 sky130_fd_sc_hd__mux4_1 c416 (.A0(net212),
    .A1(net215),
    .A2(net197),
    .A3(net214),
    .S0(net211),
    .S1(net213),
    .X(net216));
 sky130_fd_sc_hd__a41o_1 c417 (.A1(net213),
    .A2(net215),
    .A3(net209),
    .A4(net214),
    .B1(net1034),
    .X(net217));
 sky130_fd_sc_hd__a41o_2 c418 (.A1(net964),
    .A2(net896),
    .A3(net933),
    .A4(net942),
    .B1(net940),
    .X(net218));
 sky130_fd_sc_hd__a41o_1 c419 (.A1(net898),
    .A2(net750),
    .A3(net742),
    .A4(net894),
    .B1(net725),
    .X(net219));
 sky130_fd_sc_hd__mux4_2 c420 (.A0(net735),
    .A1(net742),
    .A2(net923),
    .A3(net897),
    .S0(net724),
    .S1(net942),
    .X(net220));
 sky130_fd_sc_hd__mux4_2 c421 (.A0(net748),
    .A1(net744),
    .A2(net218),
    .A3(net933),
    .S0(net1020),
    .S1(net640),
    .X(net221));
 sky130_fd_sc_hd__mux4_2 c422 (.A0(net214),
    .A1(net123),
    .A2(net946),
    .A3(net760),
    .S0(net221),
    .S1(net964),
    .X(net222));
 sky130_fd_sc_hd__mux4_2 c423 (.A0(net212),
    .A1(net218),
    .A2(net221),
    .A3(net965),
    .S0(net906),
    .S1(net908),
    .X(net223));
 sky130_fd_sc_hd__mux4_1 c424 (.A0(net211),
    .A1(net750),
    .A2(net223),
    .A3(net1077),
    .S0(net220),
    .S1(net893),
    .X(net224));
 sky130_fd_sc_hd__a41o_2 c425 (.A1(net9),
    .A2(net894),
    .A3(net950),
    .A4(net896),
    .B1(net945),
    .X(net225));
 sky130_fd_sc_hd__mux4_1 c426 (.A0(net759),
    .A1(net221),
    .A2(net222),
    .A3(net919),
    .S0(net942),
    .S1(net640),
    .X(net226));
 sky130_fd_sc_hd__mux4_2 c427 (.A0(net218),
    .A1(net901),
    .A2(net9),
    .A3(net564),
    .S0(net640),
    .S1(net660),
    .X(net227));
 sky130_fd_sc_hd__mux4_1 c428 (.A0(net725),
    .A1(net211),
    .A2(net117),
    .A3(net999),
    .S0(net196),
    .S1(net847),
    .X(net228));
 sky130_fd_sc_hd__a41o_1 c429 (.A1(net227),
    .A2(net219),
    .A3(net220),
    .A4(net555),
    .B1(net660),
    .X(net229));
 sky130_fd_sc_hd__a41o_2 c430 (.A1(net221),
    .A2(net742),
    .A3(net936),
    .A4(net225),
    .B1(net660),
    .X(net230));
 sky130_fd_sc_hd__sdfbbn_2 c431 (.CLK_N(clknet_4_9_0_clk),
    .D(net230),
    .RESET_B(net1023),
    .SCD(net744),
    .SCE(net223),
    .SET_B(net1027),
    .Q(net884),
    .Q_N(net231));
 sky130_fd_sc_hd__mux4_1 c432 (.A0(net230),
    .A1(net993),
    .A2(net128),
    .A3(net129),
    .S0(net221),
    .S1(net661),
    .X(net232));
 sky130_fd_sc_hd__mux4_2 c433 (.A0(net227),
    .A1(net106),
    .A2(net884),
    .A3(net128),
    .S0(net225),
    .S1(net657),
    .X(net233));
 sky130_fd_sc_hd__mux4_1 c434 (.A0(net223),
    .A1(net230),
    .A2(net231),
    .A3(net229),
    .S0(net847),
    .S1(net1027),
    .X(net234));
 sky130_fd_sc_hd__mux4_1 c435 (.A0(net38),
    .A1(net884),
    .A2(net222),
    .A3(net225),
    .S0(net212),
    .S1(net663),
    .X(net235));
 sky130_fd_sc_hd__mux4_1 c436 (.A0(net110),
    .A1(net980),
    .A2(net923),
    .A3(net233),
    .S0(net1037),
    .S1(net1029),
    .X(net236));
 sky130_fd_sc_hd__mux4_1 c437 (.A0(net202),
    .A1(net229),
    .A2(net28),
    .A3(net536),
    .S0(net847),
    .S1(net662),
    .X(net237));
 sky130_fd_sc_hd__mux4_2 c438 (.A0(net959),
    .A1(net897),
    .A2(net735),
    .A3(net896),
    .S0(net971),
    .S1(net661),
    .X(net238));
 sky130_fd_sc_hd__mux4_1 c439 (.A0(net28),
    .A1(net230),
    .A2(net233),
    .A3(net535),
    .S0(net847),
    .S1(net665),
    .X(net239));
 sky130_fd_sc_hd__mux4_2 c440 (.A0(net59),
    .A1(net993),
    .A2(net192),
    .A3(net907),
    .S0(net945),
    .S1(net661),
    .X(net240));
 sky130_fd_sc_hd__mux4_2 c441 (.A0(net106),
    .A1(net28),
    .A2(net755),
    .A3(net772),
    .S0(net944),
    .S1(net660),
    .X(net848));
 sky130_fd_sc_hd__mux4_2 c442 (.A0(net772),
    .A1(net201),
    .A2(net109),
    .A3(net956),
    .S0(net195),
    .S1(net962),
    .X(net241));
 sky130_fd_sc_hd__mux4_1 c443 (.A0(net153),
    .A1(net968),
    .A2(net942),
    .A3(net865),
    .S0(net640),
    .S1(net938),
    .X(net242));
 sky130_fd_sc_hd__mux4_2 c444 (.A0(net109),
    .A1(net761),
    .A2(net962),
    .A3(net892),
    .S0(net46),
    .S1(net971),
    .X(net243));
 sky130_fd_sc_hd__mux4_2 c445 (.A0(net759),
    .A1(net59),
    .A2(net738),
    .A3(net238),
    .S0(net116),
    .S1(net741),
    .X(net830));
 sky130_fd_sc_hd__mux4_1 c446 (.A0(net47),
    .A1(clknet_1_0__leaf_net155),
    .A2(net830),
    .A3(net977),
    .S0(net865),
    .S1(net667),
    .X(net244));
 sky130_fd_sc_hd__mux4_1 c447 (.A0(net220),
    .A1(net830),
    .A2(net209),
    .A3(net956),
    .S0(net564),
    .S1(net628),
    .X(net245));
 sky130_fd_sc_hd__mux4_1 c448 (.A0(net19),
    .A1(net963),
    .A2(net106),
    .A3(net640),
    .S0(net648),
    .S1(net938),
    .X(net246));
 sky130_fd_sc_hd__mux4_1 c449 (.A0(net209),
    .A1(net839),
    .A2(net243),
    .A3(net961),
    .S0(net1039),
    .S1(net1026),
    .X(net247));
 sky130_fd_sc_hd__mux4_1 c450 (.A0(net243),
    .A1(net56),
    .A2(net776),
    .A3(net539),
    .S0(net551),
    .S1(net666),
    .X(net248));
 sky130_fd_sc_hd__mux4_2 c451 (.A0(net738),
    .A1(net212),
    .A2(net231),
    .A3(net527),
    .S0(net646),
    .S1(net668),
    .X(net249));
 sky130_fd_sc_hd__mux4_1 c452 (.A0(net246),
    .A1(clknet_1_0__leaf_net155),
    .A2(net753),
    .A3(net249),
    .S0(net539),
    .S1(net847),
    .X(net250));
 sky130_fd_sc_hd__mux4_1 c453 (.A0(net28),
    .A1(net60),
    .A2(clknet_1_0__leaf_net155),
    .A3(net243),
    .S0(net846),
    .S1(net668),
    .X(net251));
 sky130_fd_sc_hd__mux4_2 c454 (.A0(net212),
    .A1(net249),
    .A2(net919),
    .A3(net628),
    .S0(net661),
    .S1(net667),
    .X(net252));
 sky130_fd_sc_hd__mux4_1 c455 (.A0(net252),
    .A1(net45),
    .A2(net249),
    .A3(net907),
    .S0(net589),
    .X(net253));
 sky130_fd_sc_hd__mux4_1 c456 (.A0(net249),
    .A1(net243),
    .A2(net539),
    .A3(net589),
    .S0(net608),
    .S1(net647),
    .X(net254));
 sky130_fd_sc_hd__mux4_1 c457 (.A0(net249),
    .A1(net891),
    .A2(net830),
    .A3(net536),
    .S0(net666),
    .S1(net668),
    .X(net255));
 sky130_fd_sc_hd__mux4_1 c458 (.A0(net750),
    .A1(net243),
    .A2(net1000),
    .A3(clknet_1_0__leaf_net250),
    .S0(net865),
    .S1(net670),
    .X(net256));
 sky130_fd_sc_hd__mux4_1 c459 (.A0(net153),
    .A1(net830),
    .A2(net220),
    .A3(net907),
    .S0(net608),
    .S1(net667),
    .X(net257));
 sky130_fd_sc_hd__mux4_1 c460 (.A0(clknet_1_0__leaf_net155),
    .A1(net219),
    .A2(net240),
    .A3(net249),
    .S0(net596),
    .S1(net670),
    .X(net258));
 sky130_fd_sc_hd__a31o_1 c461 (.A1(net608),
    .A2(net649),
    .A3(net669),
    .B1(net670),
    .X(net259));
 sky130_fd_sc_hd__mux4_2 c462 (.A0(net143),
    .A1(net259),
    .A2(net164),
    .A3(net907),
    .S0(net754),
    .S1(net801),
    .X(net260));
 sky130_fd_sc_hd__mux4_2 c463 (.A0(net225),
    .A1(net754),
    .A2(net963),
    .A3(net967),
    .S0(net983),
    .S1(net629),
    .X(net829));
 sky130_fd_sc_hd__mux4_1 c464 (.A0(net764),
    .A1(net769),
    .A2(net1006),
    .A3(net839),
    .S0(net68),
    .S1(net958),
    .X(net261));
 sky130_fd_sc_hd__mux4_2 c465 (.A0(net238),
    .A1(net848),
    .A2(net1008),
    .A3(net957),
    .S0(net898),
    .S1(net605),
    .X(net262));
 sky130_fd_sc_hd__mux4_1 c466 (.A0(net788),
    .A1(net1007),
    .A2(net829),
    .A3(net741),
    .S0(net261),
    .S1(clknet_1_1__leaf_net630),
    .X(net263));
 sky130_fd_sc_hd__mux4_1 c467 (.A0(net238),
    .A1(net1014),
    .A2(net848),
    .A3(net617),
    .S0(net642),
    .S1(net648),
    .X(net264));
 sky130_fd_sc_hd__mux4_1 c468 (.A0(net170),
    .A1(net264),
    .A2(net829),
    .A3(net1014),
    .S0(net584),
    .S1(clknet_1_1__leaf_net651),
    .X(net265));
 sky130_fd_sc_hd__mux4_1 c469 (.A0(clknet_1_1__leaf_net174),
    .A1(net841),
    .A2(net980),
    .A3(clknet_1_0__leaf_net177),
    .S0(net553),
    .S1(net641),
    .X(net266));
 sky130_fd_sc_hd__mux4_1 c470 (.A0(net805),
    .A1(clknet_1_0__leaf_net176),
    .A2(net984),
    .A3(net828),
    .S0(net170),
    .S1(clknet_1_0__leaf_net652),
    .X(net267));
 sky130_fd_sc_hd__mux4_2 c471 (.A0(net129),
    .A1(net805),
    .A2(net764),
    .A3(net227),
    .S0(net617),
    .S1(net649),
    .X(net268));
 sky130_fd_sc_hd__mux4_1 c472 (.A0(net56),
    .A1(clknet_1_1__leaf_net177),
    .A2(net829),
    .A3(net801),
    .S0(net953),
    .S1(net553),
    .X(net269));
 sky130_fd_sc_hd__mux4_2 c473 (.A0(net828),
    .A1(net262),
    .A2(net983),
    .A3(net238),
    .S0(net835),
    .S1(net641),
    .X(net270));
 sky130_fd_sc_hd__mux4_1 c474 (.A0(net270),
    .A1(net260),
    .A2(net243),
    .A3(net268),
    .S0(net539),
    .S1(net605),
    .X(net271));
 sky130_fd_sc_hd__mux4_1 c475 (.A0(net776),
    .A1(net947),
    .A2(net984),
    .A3(net852),
    .S0(net584),
    .S1(net615),
    .X(net272));
 sky130_fd_sc_hd__mux4_1 c476 (.A0(net264),
    .A1(net958),
    .A2(clknet_1_1__leaf_net174),
    .A3(net1002),
    .S0(net596),
    .S1(net617),
    .X(net273));
 sky130_fd_sc_hd__mux4_1 c477 (.A0(net273),
    .A1(net221),
    .A2(net272),
    .A3(net1017),
    .S0(net79),
    .S1(net593),
    .X(net274));
 sky130_fd_sc_hd__mux4_2 c478 (.A0(net986),
    .A1(net841),
    .A2(net956),
    .A3(net527),
    .S0(net942),
    .S1(net608),
    .X(net275));
 sky130_fd_sc_hd__mux4_1 c479 (.A0(net261),
    .A1(net272),
    .A2(net791),
    .A3(net275),
    .S0(net944),
    .S1(clknet_1_0__leaf_net671),
    .X(net276));
 sky130_fd_sc_hd__mux4_1 c480 (.A0(net266),
    .A1(net156),
    .A2(net275),
    .A3(clknet_1_0__leaf_net276),
    .S0(net791),
    .S1(net830),
    .X(net277));
 sky130_fd_sc_hd__mux4_1 c481 (.A0(net829),
    .A1(net268),
    .A2(clknet_1_1__leaf_net276),
    .A3(net275),
    .S0(net527),
    .S1(clknet_1_0__leaf_net671),
    .X(net278));
 sky130_fd_sc_hd__mux4_1 c482 (.A0(net240),
    .A1(net275),
    .A2(net985),
    .A3(clknet_1_1__leaf_net836),
    .S0(net880),
    .S1(net617),
    .X(net279));
 sky130_fd_sc_hd__mux4_1 c483 (.A0(clknet_1_0__leaf_net276),
    .A1(net275),
    .A2(net270),
    .A3(net613),
    .S0(clknet_1_1__leaf_net651),
    .S1(clknet_1_0__leaf_net652),
    .X(net280));
 sky130_fd_sc_hd__mux4_1 c484 (.A0(net87),
    .A1(net977),
    .A2(clknet_1_1__leaf_net836),
    .A3(net962),
    .S0(net785),
    .S1(net606),
    .X(net281));
 sky130_fd_sc_hd__mux4_1 c485 (.A0(net761),
    .A1(net974),
    .A2(net1011),
    .A3(net753),
    .S0(net1),
    .S1(net817),
    .X(net282));
 sky130_fd_sc_hd__mux4_1 c486 (.A0(net757),
    .A1(net738),
    .A2(net928),
    .A3(net1),
    .S0(net586),
    .S1(net648),
    .X(net283));
 sky130_fd_sc_hd__mux4_1 c487 (.A0(net1),
    .A1(net1008),
    .A2(net902),
    .A3(net963),
    .S0(net3),
    .S1(net660),
    .X(net284));
 sky130_fd_sc_hd__mux4_1 c488 (.A0(net268),
    .A1(net951),
    .A2(net87),
    .A3(net817),
    .S0(net615),
    .S1(clknet_1_1__leaf_net632),
    .X(net285));
 sky130_fd_sc_hd__mux4_1 c489 (.A0(net859),
    .A1(net182),
    .A2(clknet_1_1__leaf_net177),
    .A3(net555),
    .S0(net614),
    .S1(clknet_1_1__leaf_net632),
    .X(net286));
 sky130_fd_sc_hd__mux4_1 c490 (.A0(clknet_1_1__leaf_net281),
    .A1(net88),
    .A2(net268),
    .A3(net835),
    .S0(net614),
    .S1(clknet_1_0__leaf_net653),
    .X(net287));
 sky130_fd_sc_hd__mux4_1 c491 (.A0(net182),
    .A1(net859),
    .A2(net1),
    .A3(net757),
    .S0(net586),
    .S1(clknet_1_0__leaf_net672),
    .X(net288));
 sky130_fd_sc_hd__mux4_1 c492 (.A0(net128),
    .A1(net1017),
    .A2(net957),
    .A3(net156),
    .S0(net829),
    .S1(net87),
    .X(net289));
 sky130_fd_sc_hd__mux4_1 c493 (.A0(net814),
    .A1(net761),
    .A2(net838),
    .A3(net628),
    .S0(net660),
    .S1(clknet_1_0__leaf_net672),
    .X(net290));
 sky130_fd_sc_hd__mux4_1 c494 (.A0(net68),
    .A1(net809),
    .A2(net947),
    .A3(clknet_1_0__leaf_net189),
    .S0(clknet_1_1__leaf_net834),
    .S1(net838),
    .X(net291));
 sky130_fd_sc_hd__mux4_1 c495 (.A0(net785),
    .A1(clknet_1_1__leaf_net853),
    .A2(net590),
    .A3(net605),
    .S0(clknet_1_0__leaf_net653),
    .S1(net667),
    .X(net292));
 sky130_fd_sc_hd__mux4_1 c496 (.A0(net284),
    .A1(net89),
    .A2(clknet_1_0__leaf_net836),
    .A3(net968),
    .S0(clknet_1_1__leaf_net632),
    .S1(net648),
    .X(net293));
 sky130_fd_sc_hd__mux4_1 c497 (.A0(clknet_1_1__leaf_net189),
    .A1(net776),
    .A2(net968),
    .A3(clknet_1_1__leaf_net834),
    .S0(net607),
    .S1(net624),
    .X(net294));
 sky130_fd_sc_hd__mux4_1 c498 (.A0(net3),
    .A1(net928),
    .A2(net89),
    .A3(net182),
    .S0(net846),
    .S1(net666),
    .X(net295));
 sky130_fd_sc_hd__mux4_1 c499 (.A0(net859),
    .A1(clknet_1_0__leaf_net177),
    .A2(net617),
    .A3(net629),
    .S0(clknet_1_0__leaf_net652),
    .S1(clknet_1_0__leaf_net653),
    .X(net296));
 sky130_fd_sc_hd__mux4_1 c500 (.A0(net814),
    .A1(net284),
    .A2(clknet_1_0__leaf_net296),
    .A3(net761),
    .S0(net543),
    .S1(net607),
    .X(net297));
 sky130_fd_sc_hd__mux4_1 c501 (.A0(net221),
    .A1(net70),
    .A2(net1017),
    .A3(net87),
    .S0(net846),
    .S1(clknet_1_0__leaf_net296),
    .X(net298));
 sky130_fd_sc_hd__mux4_1 c502 (.A0(net738),
    .A1(clknet_1_1__leaf_net292),
    .A2(clknet_1_1__leaf_net296),
    .A3(clknet_1_1__leaf_net834),
    .S0(net838),
    .S1(net615),
    .X(net299));
 sky130_fd_sc_hd__mux4_1 c503 (.A0(net282),
    .A1(net791),
    .A2(clknet_1_1__leaf_net296),
    .A3(net869),
    .S0(clknet_1_0__leaf_net651),
    .S1(clknet_1_0__leaf_net672),
    .X(net300));
 sky130_fd_sc_hd__mux4_1 c504 (.A0(clknet_1_0__leaf_net292),
    .A1(net293),
    .A2(net849),
    .A3(clknet_1_0__leaf_net281),
    .S0(clknet_1_0__leaf_net296),
    .S1(net607),
    .X(net301));
 sky130_fd_sc_hd__mux4_1 c505 (.A0(clknet_1_1__leaf_net296),
    .A1(net182),
    .A2(net951),
    .A3(net837),
    .S0(net590),
    .S1(net607),
    .X(net302));
 sky130_fd_sc_hd__a41o_2 c528 (.A1(net933),
    .A2(net1042),
    .A3(net966),
    .A4(net912),
    .B1(net637),
    .X(net303));
 sky130_fd_sc_hd__a41o_1 c529 (.A1(net735),
    .A2(net116),
    .A3(net971),
    .A4(net951),
    .B1(net656),
    .X(net304));
 sky130_fd_sc_hd__mux4_1 c530 (.A0(net975),
    .A1(net102),
    .A2(net951),
    .A3(net889),
    .S0(net1042),
    .S1(net658),
    .X(net305));
 sky130_fd_sc_hd__mux4_1 c531 (.A0(net203),
    .A1(net926),
    .A2(net998),
    .A3(net889),
    .S0(net953),
    .S1(net654),
    .X(net306));
 sky130_fd_sc_hd__mux4_2 c532 (.A0(net1010),
    .A1(net205),
    .A2(net208),
    .A3(net964),
    .S0(net659),
    .S1(net674),
    .X(net307));
 sky130_fd_sc_hd__sdfbbp_1 c533 (.CLK(clknet_4_11_0_clk),
    .D(net108),
    .RESET_B(net198),
    .SCD(net889),
    .SCE(net303),
    .SET_B(net1025),
    .Q(net309),
    .Q_N(net308));
 sky130_fd_sc_hd__mux4_1 c534 (.A0(net215),
    .A1(net953),
    .A2(net116),
    .A3(net203),
    .S0(net303),
    .S1(net926),
    .X(net310));
 sky130_fd_sc_hd__mux4_1 c535 (.A0(net996),
    .A1(net894),
    .A2(net934),
    .A3(net972),
    .S0(net966),
    .S1(net889),
    .X(net311));
 sky130_fd_sc_hd__mux4_1 c536 (.A0(net108),
    .A1(net115),
    .A2(net1054),
    .A3(net889),
    .S0(net674),
    .S1(net677),
    .X(net312));
 sky130_fd_sc_hd__sdfbbn_1 c537 (.CLK_N(clknet_4_11_0_clk),
    .D(net953),
    .RESET_B(net889),
    .SCD(net934),
    .SCE(net972),
    .SET_B(clknet_1_1__leaf_net673),
    .Q(net314),
    .Q_N(net313));
 sky130_fd_sc_hd__mux4_2 c538 (.A0(net303),
    .A1(net926),
    .A2(net529),
    .A3(net941),
    .S0(clknet_1_1__leaf_net673),
    .S1(net675),
    .X(net315));
 sky130_fd_sc_hd__mux4_1 c539 (.A0(net313),
    .A1(clknet_1_1__leaf_net315),
    .A2(net308),
    .A3(net303),
    .S0(net529),
    .S1(clknet_1_1__leaf_net673),
    .X(net316));
 sky130_fd_sc_hd__mux4_1 c540 (.A0(clknet_1_1__leaf_net315),
    .A1(net975),
    .A2(net199),
    .A3(net933),
    .S0(net545),
    .S1(net678),
    .X(net317));
 sky130_fd_sc_hd__mux4_1 c541 (.A0(net756),
    .A1(clknet_1_1__leaf_net316),
    .A2(clknet_1_1__leaf_net317),
    .A3(net894),
    .S0(net108),
    .S1(net674),
    .X(net318));
 sky130_fd_sc_hd__mux4_1 c542 (.A0(clknet_1_1__leaf_net316),
    .A1(clknet_1_0__leaf_net317),
    .A2(net104),
    .A3(net196),
    .S0(net888),
    .S1(net567),
    .X(net319));
 sky130_fd_sc_hd__mux4_1 c543 (.A0(clknet_1_1__leaf_net317),
    .A1(net313),
    .A2(net745),
    .A3(net889),
    .S0(clknet_1_1__leaf_net673),
    .S1(net679),
    .X(net320));
 sky130_fd_sc_hd__mux4_1 c544 (.A0(net208),
    .A1(clknet_1_1__leaf_net318),
    .A2(net314),
    .A3(net109),
    .S0(net677),
    .S1(net680),
    .X(net321));
 sky130_fd_sc_hd__mux4_1 c545 (.A0(net889),
    .A1(clknet_1_1__leaf_net318),
    .A2(clknet_1_1__leaf_net321),
    .A3(net307),
    .S0(net529),
    .S1(clknet_1_1__leaf_net673),
    .X(net322));
 sky130_fd_sc_hd__mux4_1 c546 (.A0(clknet_1_1__leaf_net321),
    .A1(net895),
    .A2(net307),
    .A3(net108),
    .S0(net681),
    .S1(net682),
    .X(net323));
 sky130_fd_sc_hd__mux4_1 c547 (.A0(clknet_1_0__leaf_net321),
    .A1(net951),
    .A2(net975),
    .A3(net676),
    .S0(net679),
    .S1(net681),
    .X(net324));
 sky130_fd_sc_hd__mux4_1 c548 (.A0(net215),
    .A1(net980),
    .A2(clknet_1_1__leaf_net318),
    .A3(net676),
    .S0(net682),
    .S1(net683),
    .X(net325));
 sky130_fd_sc_hd__mux4_2 c549 (.A0(net205),
    .A1(net1041),
    .A2(net529),
    .A3(net675),
    .S0(net681),
    .S1(net684),
    .X(net326));
 sky130_fd_sc_hd__mux4_2 c550 (.A0(net303),
    .A1(net918),
    .A2(net970),
    .A3(net926),
    .S0(net945),
    .S1(net940),
    .X(net327));
 sky130_fd_sc_hd__mux4_1 c551 (.A0(net213),
    .A1(net307),
    .A2(net115),
    .A3(net230),
    .S0(net955),
    .S1(net663),
    .X(net328));
 sky130_fd_sc_hd__mux4_1 c552 (.A0(net34),
    .A1(net923),
    .A2(net229),
    .A3(net737),
    .S0(net654),
    .S1(net657),
    .X(net329));
 sky130_fd_sc_hd__mux4_1 c553 (.A0(net230),
    .A1(net972),
    .A2(net1066),
    .A3(net661),
    .S0(net664),
    .S1(net1035),
    .X(net330));
 sky130_fd_sc_hd__mux4_1 c554 (.A0(net327),
    .A1(net118),
    .A2(net946),
    .A3(clknet_1_0__leaf_net577),
    .S0(net663),
    .S1(net687),
    .X(net331));
 sky130_fd_sc_hd__mux4_1 c555 (.A0(net115),
    .A1(net218),
    .A2(net308),
    .A3(net980),
    .S0(net931),
    .S1(net912),
    .X(net332));
 sky130_fd_sc_hd__mux4_2 c556 (.A0(net332),
    .A1(net964),
    .A2(net966),
    .A3(net327),
    .S0(net945),
    .S1(net683),
    .X(net333));
 sky130_fd_sc_hd__mux4_1 c557 (.A0(net222),
    .A1(net117),
    .A2(net327),
    .A3(net737),
    .S0(net945),
    .S1(net845),
    .X(net334));
 sky130_fd_sc_hd__mux4_1 c558 (.A0(net122),
    .A1(net907),
    .A2(net303),
    .A3(net309),
    .S0(net737),
    .S1(net688),
    .X(net335));
 sky130_fd_sc_hd__mux4_1 c559 (.A0(net332),
    .A1(net133),
    .A2(net535),
    .A3(clknet_1_0__leaf_net577),
    .S0(net688),
    .S1(net690),
    .X(net336));
 sky130_fd_sc_hd__mux4_1 c560 (.A0(net229),
    .A1(net104),
    .A2(net332),
    .A3(net685),
    .S0(net690),
    .S1(net831),
    .X(net337));
 sky130_fd_sc_hd__mux4_1 c561 (.A0(net926),
    .A1(net897),
    .A2(net945),
    .A3(clknet_1_0__leaf_net577),
    .S0(net662),
    .S1(net690),
    .X(net338));
 sky130_fd_sc_hd__mux4_2 c562 (.A0(net1075),
    .A1(net205),
    .A2(net955),
    .A3(net115),
    .S0(net680),
    .S1(net687),
    .X(net339));
 sky130_fd_sc_hd__mux4_1 c563 (.A0(net335),
    .A1(net326),
    .A2(net567),
    .A3(net689),
    .S0(net690),
    .S1(net831),
    .X(net340));
 sky130_fd_sc_hd__mux4_1 c564 (.A0(net894),
    .A1(net340),
    .A2(clknet_1_1__leaf_net338),
    .A3(net197),
    .S0(net940),
    .S1(net831),
    .X(net341));
 sky130_fd_sc_hd__mux4_1 c565 (.A0(net340),
    .A1(net219),
    .A2(net339),
    .A3(net567),
    .S0(net690),
    .S1(clknet_1_1__leaf_net692),
    .X(net342));
 sky130_fd_sc_hd__mux4_1 c566 (.A0(clknet_1_0__leaf_net338),
    .A1(net760),
    .A2(net335),
    .A3(net529),
    .S0(net831),
    .S1(clknet_1_0__leaf_net693),
    .X(net343));
 sky130_fd_sc_hd__mux4_1 c567 (.A0(net335),
    .A1(net333),
    .A2(net327),
    .A3(net664),
    .S0(net831),
    .S1(clknet_1_1__leaf_net693),
    .X(net344));
 sky130_fd_sc_hd__mux4_1 c568 (.A0(clknet_1_0__leaf_net343),
    .A1(net197),
    .A2(net893),
    .A3(net535),
    .S0(net663),
    .S1(clknet_1_0__leaf_net693),
    .X(net345));
 sky130_fd_sc_hd__mux4_1 c569 (.A0(net222),
    .A1(net936),
    .A2(net127),
    .A3(clknet_1_0__leaf_net343),
    .S0(net340),
    .S1(clknet_1_1__leaf_net692),
    .X(net346));
 sky130_fd_sc_hd__mux4_1 c570 (.A0(net333),
    .A1(clknet_1_1__leaf_net343),
    .A2(net229),
    .A3(net664),
    .S0(clknet_1_1__leaf_net692),
    .S1(clknet_1_1__leaf_net693),
    .X(net347));
 sky130_fd_sc_hd__mux4_1 c571 (.A0(net229),
    .A1(net309),
    .A2(net326),
    .S0(net831),
    .S1(clknet_1_1__leaf_net692),
    .X(net348));
 sky130_fd_sc_hd__mux4_1 c572 (.A0(net307),
    .A1(clknet_1_0__leaf_net315),
    .A2(net57),
    .A3(net521),
    .S0(net647),
    .S1(net685),
    .X(net349));
 sky130_fd_sc_hd__mux4_1 c573 (.A0(net45),
    .A1(net936),
    .A2(net196),
    .A3(net755),
    .S0(net1019),
    .S1(net647),
    .X(net350));
 sky130_fd_sc_hd__mux4_1 c574 (.A0(net104),
    .A1(net223),
    .A2(net961),
    .A3(net962),
    .S0(net1033),
    .S1(net681),
    .X(net351));
 sky130_fd_sc_hd__mux4_1 c575 (.A0(net246),
    .A1(net974),
    .A2(clknet_1_0__leaf_net250),
    .A3(net243),
    .S0(net252),
    .S1(net956),
    .X(net352));
 sky130_fd_sc_hd__mux4_2 c576 (.A0(net122),
    .A1(net915),
    .A2(net655),
    .A3(net667),
    .S0(net669),
    .S1(net690),
    .X(net353));
 sky130_fd_sc_hd__mux4_1 c577 (.A0(net219),
    .A1(net243),
    .A2(net884),
    .A3(net53),
    .S0(net936),
    .S1(net1028),
    .X(net354));
 sky130_fd_sc_hd__mux4_1 c578 (.A0(clknet_1_0__leaf_net250),
    .A1(net769),
    .A2(net753),
    .A3(net893),
    .S0(net621),
    .S1(net665),
    .X(net355));
 sky130_fd_sc_hd__mux4_1 c579 (.A0(net196),
    .A1(net249),
    .A2(net760),
    .A3(clknet_1_1__leaf_net155),
    .S0(net845),
    .S1(net597),
    .X(net356));
 sky130_fd_sc_hd__mux4_1 c580 (.A0(net252),
    .A1(net241),
    .A2(net895),
    .A3(net259),
    .S0(net649),
    .S1(net655),
    .X(net357));
 sky130_fd_sc_hd__mux4_1 c581 (.A0(net1066),
    .A1(net145),
    .A2(net241),
    .A3(net209),
    .S0(net972),
    .S1(net695),
    .X(net358));
 sky130_fd_sc_hd__mux4_1 c582 (.A0(net1009),
    .A1(clknet_1_0__leaf_net250),
    .A2(net621),
    .A3(net686),
    .S0(net690),
    .S1(net698),
    .X(net359));
 sky130_fd_sc_hd__mux4_1 c583 (.A0(net309),
    .A1(clknet_1_1__leaf_net349),
    .A2(net891),
    .A3(net1001),
    .S0(net647),
    .S1(net698),
    .X(net360));
 sky130_fd_sc_hd__mux4_1 c584 (.A0(net249),
    .A1(net227),
    .A2(net895),
    .A3(net252),
    .S0(net907),
    .S1(net699),
    .X(net361));
 sky130_fd_sc_hd__mux4_1 c585 (.A0(net49),
    .A1(net201),
    .A2(net978),
    .A3(net200),
    .S0(net563),
    .S1(net621),
    .X(net362));
 sky130_fd_sc_hd__mux4_1 c586 (.A0(net361),
    .A1(net931),
    .A2(net20),
    .A3(net597),
    .S0(net655),
    .S1(net670),
    .X(net363));
 sky130_fd_sc_hd__mux4_1 c587 (.A0(net962),
    .A1(net57),
    .A2(net124),
    .A3(net741),
    .S0(net588),
    .S1(net649),
    .X(net364));
 sky130_fd_sc_hd__mux4_1 c588 (.A0(net967),
    .A1(net57),
    .A2(net45),
    .A3(net644),
    .S0(net697),
    .S1(net699),
    .X(net365));
 sky130_fd_sc_hd__mux4_1 c589 (.A0(clknet_1_1__leaf_net349),
    .A1(net748),
    .A2(net1005),
    .A3(net895),
    .S0(net362),
    .S1(net697),
    .X(net366));
 sky130_fd_sc_hd__mux4_1 c590 (.A0(clknet_1_1__leaf_net359),
    .A1(clknet_1_0__leaf_net317),
    .A2(clknet_1_1__leaf_net250),
    .A3(net654),
    .S0(net674),
    .S1(net700),
    .X(net367));
 sky130_fd_sc_hd__mux4_1 c591 (.A0(net1066),
    .A1(net897),
    .A2(net963),
    .A3(net120),
    .S0(net536),
    .S1(net827),
    .X(net368));
 sky130_fd_sc_hd__mux4_1 c592 (.A0(clknet_1_0__leaf_net359),
    .A1(net361),
    .A2(net589),
    .A3(net666),
    .S0(net696),
    .S1(net827),
    .X(net369));
 sky130_fd_sc_hd__mux4_1 c593 (.A0(net146),
    .A1(net1077),
    .A2(clknet_1_1__leaf_net355),
    .A3(clknet_1_1__leaf_net155),
    .S0(net529),
    .S1(net700),
    .X(net370));
 sky130_fd_sc_hd__mux4_1 c594 (.A0(clknet_1_1__leaf_net174),
    .A1(net120),
    .A2(net757),
    .A3(net959),
    .S0(net963),
    .S1(net831),
    .X(net371));
 sky130_fd_sc_hd__mux4_1 c595 (.A0(net922),
    .A1(net1067),
    .A2(net801),
    .A3(net907),
    .S0(net69),
    .S1(net587),
    .X(net372));
 sky130_fd_sc_hd__mux4_1 c596 (.A0(clknet_1_0__leaf_net176),
    .A1(clknet_1_0__leaf_net355),
    .A2(net36),
    .A3(net231),
    .S0(net837),
    .S1(clknet_1_0__leaf_net671),
    .X(net373));
 sky130_fd_sc_hd__mux4_1 c597 (.A0(net744),
    .A1(clknet_1_0__leaf_net345),
    .A2(net117),
    .A3(net801),
    .S0(net880),
    .S1(clknet_1_1__leaf_net652),
    .X(net374));
 sky130_fd_sc_hd__mux4_1 c598 (.A0(net196),
    .A1(net1003),
    .A2(net801),
    .A3(clknet_1_0__leaf_net345),
    .S0(net825),
    .S1(net702),
    .X(net375));
 sky130_fd_sc_hd__mux4_1 c599 (.A0(net67),
    .A1(net1001),
    .A2(net769),
    .A3(net741),
    .S0(net120),
    .S1(net675),
    .X(net376));
 sky130_fd_sc_hd__mux4_1 c600 (.A0(net762),
    .A1(net243),
    .A2(net53),
    .A3(clknet_1_1__leaf_net174),
    .S0(net832),
    .S1(net957),
    .X(net377));
 sky130_fd_sc_hd__mux4_1 c601 (.A0(net36),
    .A1(net196),
    .A2(net1069),
    .A3(net604),
    .S0(net940),
    .S1(clknet_1_0__leaf_net692),
    .X(net378));
 sky130_fd_sc_hd__mux4_1 c602 (.A0(net270),
    .A1(net117),
    .A2(net231),
    .A3(net75),
    .S0(net681),
    .S1(net683),
    .X(net379));
 sky130_fd_sc_hd__mux4_1 c603 (.A0(net968),
    .A1(clknet_1_0__leaf_net315),
    .A2(net829),
    .A3(clknet_1_1__leaf_net355),
    .S0(net600),
    .S1(net669),
    .X(net380));
 sky130_fd_sc_hd__mux4_2 c604 (.A0(net260),
    .A1(net353),
    .A2(net919),
    .A3(net1002),
    .S0(clknet_1_1__leaf_net630),
    .S1(net703),
    .X(net381));
 sky130_fd_sc_hd__mux4_1 c605 (.A0(net1068),
    .A1(net69),
    .A2(net120),
    .A3(clknet_1_0__leaf_net349),
    .S0(net603),
    .S1(net619),
    .X(net382));
 sky130_fd_sc_hd__mux4_1 c606 (.A0(net801),
    .A1(clknet_1_0__leaf_net349),
    .A2(net79),
    .A3(net832),
    .S0(net601),
    .S1(net703),
    .X(net383));
 sky130_fd_sc_hd__mux4_1 c607 (.A0(clknet_1_1__leaf_net345),
    .A1(net109),
    .A2(net968),
    .A3(net619),
    .S0(net683),
    .S1(net703),
    .X(net384));
 sky130_fd_sc_hd__mux4_1 c608 (.A0(net116),
    .A1(clknet_1_0__leaf_net371),
    .A2(clknet_1_1__leaf_net177),
    .A3(net961),
    .S0(net938),
    .S1(net669),
    .X(net385));
 sky130_fd_sc_hd__mux4_1 c609 (.A0(net79),
    .A1(clknet_1_1__leaf_net371),
    .A2(net754),
    .A3(net593),
    .S0(net603),
    .S1(net677),
    .X(net386));
 sky130_fd_sc_hd__mux4_1 c610 (.A0(clknet_1_1__leaf_net386),
    .A1(net195),
    .A2(net959),
    .A3(net262),
    .S0(net587),
    .S1(net649),
    .X(net387));
 sky130_fd_sc_hd__mux4_1 c611 (.A0(net333),
    .A1(net1014),
    .A2(clknet_1_0__leaf_net386),
    .A3(net959),
    .S0(net603),
    .S1(net703),
    .X(net388));
 sky130_fd_sc_hd__mux4_2 c612 (.A0(net381),
    .A1(net972),
    .A2(net957),
    .A3(net25),
    .S0(net940),
    .S1(net681),
    .X(net389));
 sky130_fd_sc_hd__mux4_1 c613 (.A0(net999),
    .A1(net988),
    .A2(clknet_1_1__leaf_net389),
    .A3(clknet_1_1__leaf_net176),
    .S0(net595),
    .S1(net603),
    .X(net390));
 sky130_fd_sc_hd__mux4_2 c614 (.A0(clknet_1_1__leaf_net389),
    .A1(net953),
    .A2(clknet_1_0__leaf_net609),
    .A3(clknet_1_0__leaf_net610),
    .S0(net702),
    .S1(net704),
    .X(net391));
 sky130_fd_sc_hd__mux4_1 c615 (.A0(net376),
    .A1(clknet_1_0__leaf_net389),
    .A2(clknet_1_1__leaf_net177),
    .A3(net748),
    .S0(net615),
    .S1(net661),
    .X(net392));
 sky130_fd_sc_hd__mux4_1 c616 (.A0(net737),
    .A1(net283),
    .A2(net828),
    .A3(net92),
    .S0(net959),
    .S1(net831),
    .X(net393));
 sky130_fd_sc_hd__mux4_2 c617 (.A0(net755),
    .A1(net842),
    .A2(net283),
    .A3(net963),
    .S0(net957),
    .S1(net529),
    .X(net394));
 sky130_fd_sc_hd__mux4_1 c618 (.A0(net774),
    .A1(clknet_1_0__leaf_net385),
    .A2(net967),
    .A3(net997),
    .S0(net826),
    .S1(net661),
    .X(net395));
 sky130_fd_sc_hd__mux4_1 c619 (.A0(net117),
    .A1(net1015),
    .A2(clknet_1_0__leaf_net389),
    .A3(net394),
    .S0(net774),
    .S1(net676),
    .X(net396));
 sky130_fd_sc_hd__mux4_1 c620 (.A0(net980),
    .A1(net60),
    .A2(net932),
    .A3(net624),
    .S0(net661),
    .S1(net703),
    .X(net397));
 sky130_fd_sc_hd__mux4_1 c621 (.A0(clknet_1_0__leaf_net355),
    .A1(net957),
    .A2(net999),
    .A3(net944),
    .S0(net619),
    .S1(net703),
    .X(net398));
 sky130_fd_sc_hd__mux4_1 c622 (.A0(net66),
    .A1(net979),
    .A2(net980),
    .A3(net353),
    .S0(net957),
    .S1(net615),
    .X(net399));
 sky130_fd_sc_hd__mux4_1 c623 (.A0(clknet_1_0__leaf_net315),
    .A1(net909),
    .A2(net980),
    .A3(net604),
    .S0(net620),
    .S1(net677),
    .X(net400));
 sky130_fd_sc_hd__mux4_2 c624 (.A0(net757),
    .A1(net47),
    .A2(net832),
    .A3(net92),
    .S0(net974),
    .S1(net675),
    .X(net401));
 sky130_fd_sc_hd__mux4_1 c625 (.A0(clknet_1_1__leaf_net177),
    .A1(net399),
    .A2(net970),
    .A3(net967),
    .S0(net642),
    .S1(clknet_1_1__leaf_net653),
    .X(net402));
 sky130_fd_sc_hd__mux4_1 c626 (.A0(net842),
    .A1(net66),
    .A2(net760),
    .A3(net909),
    .S0(net614),
    .S1(net665),
    .X(net403));
 sky130_fd_sc_hd__mux4_1 c627 (.A0(net259),
    .A1(net60),
    .A2(net757),
    .A3(clknet_1_0__leaf_net400),
    .S0(net615),
    .S1(clknet_1_0__leaf_net672),
    .X(net404));
 sky130_fd_sc_hd__mux4_1 c628 (.A0(net957),
    .A1(net739),
    .A2(net1011),
    .A3(net830),
    .S0(clknet_1_1__leaf_net355),
    .S1(net599),
    .X(net405));
 sky130_fd_sc_hd__mux4_1 c629 (.A0(net989),
    .A1(net755),
    .A2(clknet_1_0__leaf_net367),
    .A3(net967),
    .S0(net944),
    .S1(net869),
    .X(net406));
 sky130_fd_sc_hd__mux4_1 c630 (.A0(net75),
    .A1(net403),
    .A2(net755),
    .A3(clknet_1_0__leaf_net367),
    .S0(net146),
    .S1(net979),
    .X(net407));
 sky130_fd_sc_hd__mux4_1 c631 (.A0(net406),
    .A1(clknet_1_0__leaf_net367),
    .A2(net774),
    .A3(net401),
    .S0(net590),
    .S1(net604),
    .X(net408));
 sky130_fd_sc_hd__mux4_1 c632 (.A0(clknet_1_1__leaf_net385),
    .A1(net408),
    .A2(net826),
    .A3(clknet_1_0__leaf_net290),
    .S0(net1014),
    .S1(clknet_1_1__leaf_net672),
    .X(net409));
 sky130_fd_sc_hd__mux4_1 c633 (.A0(net353),
    .A1(net92),
    .A2(net814),
    .A3(clknet_1_0__leaf_net400),
    .S0(net607),
    .S1(net661),
    .X(net410));
 sky130_fd_sc_hd__mux4_1 c634 (.A0(net402),
    .A1(net799),
    .A2(net584),
    .A3(net611),
    .S0(clknet_1_1__leaf_net671),
    .S1(net700),
    .X(net411));
 sky130_fd_sc_hd__mux4_1 c635 (.A0(net905),
    .A1(net579),
    .A2(net602),
    .A3(net604),
    .S0(net611),
    .S1(net620),
    .X(net412));
 sky130_fd_sc_hd__mux4_1 c636 (.A0(net410),
    .A1(net401),
    .A2(net832),
    .A3(clknet_1_0__leaf_net355),
    .S0(net602),
    .S1(net703),
    .X(net413));
 sky130_fd_sc_hd__mux4_1 c637 (.A0(net282),
    .A1(net974),
    .A2(net394),
    .A3(net869),
    .S0(net611),
    .S1(net620),
    .X(net414));
 sky130_fd_sc_hd__mux4_1 c660 (.A0(net998),
    .A1(net728),
    .A2(net326),
    .A3(net978),
    .S0(net953),
    .S1(net1032),
    .X(net415));
 sky130_fd_sc_hd__mux4_2 c661 (.A0(net978),
    .A1(net931),
    .A2(net22),
    .A3(net895),
    .S0(net545),
    .S1(net567),
    .X(net416));
 sky130_fd_sc_hd__mux4_2 c662 (.A0(net895),
    .A1(net953),
    .A2(net745),
    .A3(net731),
    .S0(net544),
    .S1(net682),
    .X(net417));
 sky130_fd_sc_hd__mux4_1 c663 (.A0(net964),
    .A1(net923),
    .A2(net889),
    .A3(net946),
    .S0(net931),
    .S1(net745),
    .X(net418));
 sky130_fd_sc_hd__mux4_1 c664 (.A0(net900),
    .A1(net1057),
    .A2(net909),
    .A3(net951),
    .S0(net922),
    .S1(net682),
    .X(net419));
 sky130_fd_sc_hd__mux4_1 c665 (.A0(net1057),
    .A1(net966),
    .A2(net419),
    .A3(net912),
    .S0(net657),
    .S1(net684),
    .X(net420));
 sky130_fd_sc_hd__mux4_2 c666 (.A0(net417),
    .A1(net953),
    .A2(net1057),
    .A3(net567),
    .S0(net682),
    .S1(net706),
    .X(net421));
 sky130_fd_sc_hd__mux4_1 c667 (.A0(net955),
    .A1(net964),
    .A2(net931),
    .A3(net888),
    .S0(net912),
    .S1(net707),
    .X(net422));
 sky130_fd_sc_hd__mux4_1 c668 (.A0(net745),
    .A1(net118),
    .A2(net415),
    .A3(net931),
    .S0(net951),
    .S1(net954),
    .X(net423));
 sky130_fd_sc_hd__mux4_2 c669 (.A0(net419),
    .A1(net922),
    .A2(net209),
    .A3(net999),
    .S0(net523),
    .S1(net706),
    .X(net424));
 sky130_fd_sc_hd__mux4_1 c670 (.A0(net415),
    .A1(net888),
    .A2(net421),
    .A3(net912),
    .S0(clknet_1_1__leaf_net673),
    .S1(net706),
    .X(net425));
 sky130_fd_sc_hd__mux4_1 c671 (.A0(net314),
    .A1(clknet_1_1__leaf_net316),
    .A2(net22),
    .A3(clknet_1_1__leaf_net673),
    .S0(net678),
    .S1(net707),
    .X(net426));
 sky130_fd_sc_hd__mux4_1 c672 (.A0(clknet_1_0__leaf_net426),
    .A1(net420),
    .A2(net999),
    .A3(net946),
    .S0(net622),
    .S1(net637),
    .X(net427));
 sky130_fd_sc_hd__a41o_1 c673 (.A1(net912),
    .A2(clknet_1_0__leaf_net426),
    .A3(net994),
    .A4(net954),
    .B1(net523),
    .X(net428));
 sky130_fd_sc_hd__mux4_1 c674 (.A0(clknet_1_1__leaf_net428),
    .A1(net731),
    .A2(net995),
    .A3(net946),
    .S0(net522),
    .S1(net708),
    .X(net429));
 sky130_fd_sc_hd__mux4_1 c675 (.A0(net888),
    .A1(clknet_1_0__leaf_net428),
    .A2(net417),
    .A3(clknet_1_1__leaf_net429),
    .S0(net912),
    .S1(net545),
    .X(net430));
 sky130_fd_sc_hd__mux4_1 c676 (.A0(net420),
    .A1(clknet_1_1__leaf_net426),
    .A2(net951),
    .A3(net684),
    .S0(net708),
    .S1(net709),
    .X(net431));
 sky130_fd_sc_hd__mux4_1 c677 (.A0(net16),
    .A1(net420),
    .A2(net424),
    .A3(net326),
    .S0(net415),
    .S1(net522),
    .X(net432));
 sky130_fd_sc_hd__mux4_1 c678 (.A0(net888),
    .A1(net912),
    .A2(net708),
    .A3(net709),
    .S0(net710),
    .S1(clknet_1_1__leaf_net711),
    .X(net433));
 sky130_fd_sc_hd__mux4_1 c679 (.A0(net421),
    .A1(net951),
    .A2(net888),
    .A3(net966),
    .S0(clknet_1_0__leaf_net673),
    .S1(net709),
    .X(net434));
 sky130_fd_sc_hd__mux4_2 c680 (.A0(net416),
    .A1(clknet_1_0__leaf_net428),
    .A2(net736),
    .A3(net927),
    .S0(net708),
    .S1(clknet_1_1__leaf_net711),
    .X(net435));
 sky130_fd_sc_hd__mux4_1 c681 (.A0(clknet_1_1__leaf_net429),
    .A1(net424),
    .A2(clknet_1_1__leaf_net435),
    .A3(net523),
    .S0(net709),
    .S1(clknet_1_1__leaf_net713),
    .X(net436));
 sky130_fd_sc_hd__mux4_1 c682 (.A0(net964),
    .A1(net198),
    .A2(net567),
    .A3(net655),
    .S0(net689),
    .S1(clknet_1_1__leaf_net711),
    .X(net437));
 sky130_fd_sc_hd__mux4_1 c683 (.A0(clknet_1_0__leaf_net318),
    .A1(net233),
    .A2(net118),
    .A3(net122),
    .S0(net900),
    .S1(net941),
    .X(net438));
 sky130_fd_sc_hd__mux4_1 c684 (.A0(net898),
    .A1(net900),
    .A2(net888),
    .A3(net1071),
    .S0(net637),
    .S1(net680),
    .X(net439));
 sky130_fd_sc_hd__mux4_1 c685 (.A0(net201),
    .A1(clknet_1_0__leaf_net318),
    .A2(net726),
    .A3(net622),
    .S0(net623),
    .S1(net710),
    .X(net440));
 sky130_fd_sc_hd__mux4_2 c686 (.A0(net218),
    .A1(net888),
    .A2(net954),
    .A3(net982),
    .S0(net680),
    .S1(net708),
    .X(net441));
 sky130_fd_sc_hd__mux4_1 c687 (.A0(net233),
    .A1(net419),
    .A2(net888),
    .A3(net935),
    .S0(clknet_1_1__leaf_net577),
    .S1(net940),
    .X(net442));
 sky130_fd_sc_hd__mux4_1 c688 (.A0(net742),
    .A1(net898),
    .A2(net327),
    .A3(net1071),
    .S0(net728),
    .S1(net637),
    .X(net443));
 sky130_fd_sc_hd__mux4_1 c689 (.A0(clknet_1_0__leaf_net435),
    .A1(clknet_1_1__leaf_net437),
    .A2(net227),
    .A3(net895),
    .S0(net327),
    .S1(net101),
    .X(net444));
 sky130_fd_sc_hd__mux4_1 c690 (.A0(net230),
    .A1(net326),
    .A2(net124),
    .A3(net417),
    .S0(net218),
    .S1(net567),
    .X(net445));
 sky130_fd_sc_hd__mux4_1 c691 (.A0(net1071),
    .A1(net339),
    .A2(clknet_1_1__leaf_net444),
    .A3(net900),
    .S0(net689),
    .S1(clknet_1_0__leaf_net711),
    .X(net446));
 sky130_fd_sc_hd__mux4_1 c692 (.A0(net739),
    .A1(clknet_1_0__leaf_net321),
    .A2(net218),
    .A3(net888),
    .S0(clknet_1_0__leaf_net316),
    .S1(clknet_1_1__leaf_net692),
    .X(net447));
 sky130_fd_sc_hd__mux4_1 c693 (.A0(net906),
    .A1(net931),
    .A2(clknet_1_0__leaf_net316),
    .A3(net520),
    .S0(net709),
    .S1(net716),
    .X(net448));
 sky130_fd_sc_hd__mux4_1 c694 (.A0(net133),
    .A1(net417),
    .A2(net326),
    .A3(net623),
    .S0(net656),
    .S1(net689),
    .X(net449));
 sky130_fd_sc_hd__mux4_1 c695 (.A0(net443),
    .A1(clknet_1_1__leaf_net448),
    .A2(clknet_1_1__leaf_net437),
    .A3(net227),
    .S0(net623),
    .S1(net684),
    .X(net450));
 sky130_fd_sc_hd__mux4_2 c696 (.A0(net339),
    .A1(clknet_1_0__leaf_net435),
    .A2(clknet_1_1__leaf_net448),
    .A3(net567),
    .S0(net570),
    .S1(net718),
    .X(net451));
 sky130_fd_sc_hd__mux4_1 c697 (.A0(net789),
    .A1(net616),
    .A2(net709),
    .A3(clknet_1_0__leaf_net711),
    .S0(net717),
    .S1(net719),
    .X(net452));
 sky130_fd_sc_hd__mux4_1 c698 (.A0(net421),
    .A1(net598),
    .A2(net616),
    .A3(net639),
    .S0(net689),
    .S1(net717),
    .X(net453));
 sky130_fd_sc_hd__mux4_1 c699 (.A0(clknet_1_0__leaf_net437),
    .A1(net811),
    .A2(net981),
    .A3(net961),
    .S0(net570),
    .S1(net716),
    .X(net454));
 sky130_fd_sc_hd__mux4_1 c700 (.A0(net900),
    .A1(net443),
    .A2(clknet_1_1__leaf_net452),
    .A3(clknet_1_1__leaf_net450),
    .S0(net569),
    .S1(net598),
    .X(net455));
 sky130_fd_sc_hd__mux4_1 c701 (.A0(clknet_1_0__leaf_net450),
    .A1(clknet_1_1__leaf_net448),
    .A2(net741),
    .A3(net569),
    .S0(net622),
    .S1(clknet_1_0__leaf_net713),
    .X(net456));
 sky130_fd_sc_hd__a41o_1 c702 (.A1(clknet_1_0__leaf_net452),
    .A2(clknet_1_1__leaf_net437),
    .A3(net520),
    .A4(net618),
    .B1(net684),
    .X(net457));
 sky130_fd_sc_hd__mux4_1 c703 (.A0(clknet_1_1__leaf_net577),
    .A1(net618),
    .A2(net941),
    .A3(net707),
    .S0(clknet_1_0__leaf_net711),
    .S1(net717),
    .X(net458));
 sky130_fd_sc_hd__mux4_1 c704 (.A0(net46),
    .A1(clknet_1_1__leaf_net250),
    .A2(clknet_1_1__leaf_net155),
    .A3(net940),
    .S0(net939),
    .S1(net694),
    .X(net459));
 sky130_fd_sc_hd__mux4_1 c705 (.A0(net30),
    .A1(clknet_1_1__leaf_net250),
    .A2(clknet_1_1__leaf_net577),
    .A3(net939),
    .S0(net645),
    .S1(net694),
    .X(net460));
 sky130_fd_sc_hd__mux4_1 c706 (.A0(net145),
    .A1(clknet_1_0__leaf_net451),
    .A2(clknet_1_0__leaf_net459),
    .A3(net909),
    .S0(net533),
    .S1(net695),
    .X(net461));
 sky130_fd_sc_hd__mux4_1 c707 (.A0(clknet_1_1__leaf_net458),
    .A1(net897),
    .A2(net962),
    .A3(net542),
    .S0(net708),
    .S1(net710),
    .X(net462));
 sky130_fd_sc_hd__mux4_1 c708 (.A0(net742),
    .A1(clknet_1_1__leaf_net367),
    .A2(net567),
    .A3(net644),
    .S0(clknet_1_0__leaf_net673),
    .S1(net708),
    .X(net463));
 sky130_fd_sc_hd__mux4_1 c709 (.A0(clknet_1_1__leaf_net459),
    .A1(clknet_1_0__leaf_net316),
    .A2(net101),
    .A3(clknet_1_0__leaf_net673),
    .S0(clknet_1_1__leaf_net691),
    .S1(net701),
    .X(net464));
 sky130_fd_sc_hd__mux4_1 c710 (.A0(net364),
    .A1(clknet_1_0__leaf_net316),
    .A2(net962),
    .A3(net618),
    .S0(net710),
    .S1(clknet_1_0__leaf_net712),
    .X(net465));
 sky130_fd_sc_hd__mux4_1 c711 (.A0(net460),
    .A1(clknet_1_0__leaf_net459),
    .A2(net124),
    .A3(net973),
    .S0(net588),
    .S1(clknet_1_0__leaf_net692),
    .X(net466));
 sky130_fd_sc_hd__mux4_1 c712 (.A0(net124),
    .A1(net935),
    .A2(net811),
    .A3(net542),
    .S0(net701),
    .S1(net714),
    .X(net467));
 sky130_fd_sc_hd__mux4_1 c713 (.A0(net362),
    .A1(net956),
    .A2(net739),
    .A3(net967),
    .S0(net698),
    .S1(net709),
    .X(net468));
 sky130_fd_sc_hd__mux4_1 c714 (.A0(net742),
    .A1(net905),
    .A2(net618),
    .A3(net701),
    .S0(clknet_1_1__leaf_net712),
    .S1(net718),
    .X(net469));
 sky130_fd_sc_hd__mux4_1 c715 (.A0(net467),
    .A1(net145),
    .A2(net368),
    .A3(clknet_1_1__leaf_net457),
    .S0(net913),
    .S1(clknet_1_0__leaf_net712),
    .X(net470));
 sky130_fd_sc_hd__mux4_1 c716 (.A0(net327),
    .A1(net424),
    .A2(clknet_1_1__leaf_net457),
    .A3(net941),
    .S0(net698),
    .S1(net710),
    .X(net471));
 sky130_fd_sc_hd__mux4_2 c717 (.A0(net368),
    .A1(net468),
    .A2(net326),
    .A3(net729),
    .S0(net13),
    .S1(net736),
    .X(net472));
 sky130_fd_sc_hd__mux4_1 c718 (.A0(net10),
    .A1(net127),
    .A2(clknet_1_1__leaf_net440),
    .A3(net57),
    .S0(net626),
    .S1(clknet_1_0__leaf_net673),
    .X(net473));
 sky130_fd_sc_hd__mux4_1 c719 (.A0(net57),
    .A1(net962),
    .A2(clknet_1_0__leaf_net457),
    .A3(net1072),
    .S0(net472),
    .S1(clknet_1_0__leaf_net713),
    .X(net474));
 sky130_fd_sc_hd__mux4_1 c720 (.A0(net789),
    .A1(net472),
    .A2(net1031),
    .A3(net1038),
    .S0(net701),
    .S1(net722),
    .X(net475));
 sky130_fd_sc_hd__mux4_1 c721 (.A0(net209),
    .A1(clknet_1_0__leaf_net458),
    .A2(net126),
    .A3(clknet_1_1__leaf_net466),
    .S0(clknet_1_1__leaf_net367),
    .S1(net580),
    .X(net476));
 sky130_fd_sc_hd__mux4_1 c722 (.A0(net476),
    .A1(net243),
    .A2(net744),
    .A3(net123),
    .S0(net472),
    .S1(net580),
    .X(net477));
 sky130_fd_sc_hd__mux4_1 c723 (.A0(net464),
    .A1(net909),
    .A2(net789),
    .A3(net542),
    .S0(net563),
    .S1(net612),
    .X(net478));
 sky130_fd_sc_hd__mux4_1 c724 (.A0(clknet_1_1__leaf_net451),
    .A1(net472),
    .A2(net618),
    .A3(net624),
    .S0(net720),
    .S1(net722),
    .X(net479));
 sky130_fd_sc_hd__mux4_1 c725 (.A0(net326),
    .A1(net754),
    .A2(net472),
    .A3(net241),
    .S0(net1073),
    .S1(net563),
    .X(net480));
 sky130_fd_sc_hd__mux4_1 c726 (.A0(net241),
    .A1(net118),
    .A2(net1004),
    .A3(net953),
    .S0(net956),
    .S1(net720),
    .X(net481));
 sky130_fd_sc_hd__mux4_1 c727 (.A0(net462),
    .A1(clknet_1_0__leaf_net457),
    .A2(net961),
    .A3(clknet_1_0__leaf_net437),
    .S0(net895),
    .S1(net655),
    .X(net482));
 sky130_fd_sc_hd__mux4_1 c728 (.A0(clknet_1_1__leaf_net463),
    .A1(net262),
    .A2(net741),
    .A3(clknet_1_1__leaf_net482),
    .S0(net618),
    .S1(net699),
    .X(net483));
 sky130_fd_sc_hd__mux4_1 c729 (.A0(clknet_1_0__leaf_net466),
    .A1(net748),
    .A2(net947),
    .A3(net612),
    .S0(net709),
    .S1(net715),
    .X(net484));
 sky130_fd_sc_hd__mux4_1 c730 (.A0(clknet_1_0__leaf_net444),
    .A1(net123),
    .A2(clknet_1_0__leaf_net466),
    .A3(net741),
    .S0(net613),
    .S1(net708),
    .X(net485));
 sky130_fd_sc_hd__mux4_1 c731 (.A0(net741),
    .A1(clknet_1_0__leaf_net483),
    .A2(net938),
    .A3(net665),
    .S0(clknet_1_0__leaf_net692),
    .S1(net705),
    .X(net486));
 sky130_fd_sc_hd__mux4_2 c732 (.A0(net53),
    .A1(net962),
    .A2(net760),
    .A3(net612),
    .S0(net715),
    .S1(net721),
    .X(net487));
 sky130_fd_sc_hd__mux4_1 c733 (.A0(clknet_1_1__leaf_net155),
    .A1(clknet_1_1__leaf_net483),
    .A2(net453),
    .A3(net581),
    .S0(clknet_1_1__leaf_net691),
    .S1(net721),
    .X(net488));
 sky130_fd_sc_hd__mux4_1 c734 (.A0(net478),
    .A1(clknet_1_1__leaf_net454),
    .A2(net753),
    .A3(net487),
    .S0(net53),
    .S1(clknet_1_0__leaf_net692),
    .X(net489));
 sky130_fd_sc_hd__mux4_1 c735 (.A0(clknet_1_0__leaf_net429),
    .A1(net947),
    .A2(net800),
    .A3(net53),
    .S0(net487),
    .S1(net721),
    .X(net490));
 sky130_fd_sc_hd__mux4_1 c736 (.A0(net69),
    .A1(net729),
    .A2(net728),
    .A3(clknet_1_0__leaf_net429),
    .S0(clknet_1_0__leaf_net463),
    .S1(clknet_1_0__leaf_net457),
    .X(net491));
 sky130_fd_sc_hd__mux4_1 c737 (.A0(clknet_1_1__leaf_net367),
    .A1(net754),
    .A2(net744),
    .A3(net123),
    .S0(net705),
    .S1(net709),
    .X(net492));
 sky130_fd_sc_hd__mux4_1 c738 (.A0(net891),
    .A1(net1077),
    .A2(net118),
    .A3(net973),
    .S0(net600),
    .S1(net601),
    .X(net493));
 sky130_fd_sc_hd__mux4_1 c739 (.A0(net895),
    .A1(clknet_1_0__leaf_net448),
    .A2(net241),
    .A3(clknet_1_0__leaf_net492),
    .S0(net755),
    .S1(clknet_1_1__leaf_net609),
    .X(net494));
 sky130_fd_sc_hd__mux4_1 c740 (.A0(net453),
    .A1(clknet_1_1__leaf_net492),
    .A2(net123),
    .A3(clknet_1_0__leaf_net448),
    .S0(net778),
    .S1(net723),
    .X(net495));
 sky130_fd_sc_hd__mux4_1 c741 (.A0(net744),
    .A1(net602),
    .A2(clknet_1_1__leaf_net609),
    .A3(net626),
    .S0(net938),
    .S1(net723),
    .X(net496));
 sky130_fd_sc_hd__mux4_1 c742 (.A0(net909),
    .A1(net469),
    .A2(clknet_1_1__leaf_net155),
    .A3(net748),
    .S0(net602),
    .S1(net616),
    .X(net497));
 sky130_fd_sc_hd__mux4_1 c743 (.A0(net484),
    .A1(net487),
    .A2(net262),
    .A3(net938),
    .S0(clknet_1_0__leaf_net691),
    .S1(net702),
    .X(net498));
 sky130_fd_sc_hd__mux4_1 c744 (.A0(clknet_1_0__leaf_net440),
    .A1(net732),
    .A2(net736),
    .A3(net617),
    .S0(net939),
    .S1(net723),
    .X(net499));
 sky130_fd_sc_hd__mux4_1 c745 (.A0(clknet_1_0__leaf_net437),
    .A1(net424),
    .A2(clknet_1_0__leaf_net482),
    .A3(clknet_1_1__leaf_net610),
    .S0(net613),
    .S1(net617),
    .X(net500));
 sky130_fd_sc_hd__mux4_1 c746 (.A0(net922),
    .A1(clknet_1_0__leaf_net454),
    .A2(clknet_1_1__leaf_net652),
    .A3(clknet_1_1__leaf_net671),
    .S0(clknet_1_0__leaf_net691),
    .S1(net708),
    .X(net501));
 sky130_fd_sc_hd__mux4_1 c747 (.A0(net1004),
    .A1(net489),
    .A2(clknet_1_1__leaf_net155),
    .A3(net616),
    .S0(net626),
    .S1(net720),
    .X(net502));
 sky130_fd_sc_hd__mux4_1 c748 (.A0(net967),
    .A1(net973),
    .A2(net639),
    .A3(net665),
    .S0(net699),
    .S1(net702),
    .X(net503));
 sky130_fd_sc_hd__mux4_1 c749 (.A0(clknet_1_1__leaf_net400),
    .A1(net979),
    .A2(net498),
    .A3(net973),
    .S0(net542),
    .S1(net655),
    .X(net504));
 sky130_fd_sc_hd__mux4_1 c750 (.A0(net502),
    .A1(net501),
    .A2(net739),
    .A3(clknet_1_1__leaf_net173),
    .S0(clknet_1_0__leaf_net609),
    .S1(net624),
    .X(net505));
 sky130_fd_sc_hd__mux4_1 c751 (.A0(net424),
    .A1(clknet_1_1__leaf_net290),
    .A2(net777),
    .A3(net601),
    .S0(net702),
    .S1(net719),
    .X(net506));
 sky130_fd_sc_hd__mux4_1 c752 (.A0(net465),
    .A1(net778),
    .A2(clknet_1_1__leaf_net173),
    .A3(net655),
    .S0(net702),
    .S1(net723),
    .X(net507));
 sky130_fd_sc_hd__mux4_1 c753 (.A0(net907),
    .A1(net824),
    .A2(net584),
    .A3(net616),
    .S0(net626),
    .S1(clknet_1_1__leaf_net671),
    .X(net508));
 sky130_fd_sc_hd__mux4_1 c754 (.A0(net913),
    .A1(net503),
    .A2(net800),
    .A3(net595),
    .S0(net599),
    .S1(clknet_1_0__leaf_net673),
    .X(net509));
 sky130_fd_sc_hd__mux4_1 c755 (.A0(net935),
    .A1(net472),
    .A2(net401),
    .A3(net753),
    .S0(clknet_1_1__leaf_net610),
    .S1(net639),
    .X(net510));
 sky130_fd_sc_hd__mux4_1 c756 (.A0(net195),
    .A1(net753),
    .A2(net393),
    .A3(net509),
    .S0(net778),
    .S1(net624),
    .X(net511));
 sky130_fd_sc_hd__mux4_1 c757 (.A0(net777),
    .A1(net30),
    .A2(net146),
    .A3(net998),
    .S0(net581),
    .S1(net699),
    .X(net512));
 sky130_fd_sc_hd__mux4_1 c758 (.A0(net118),
    .A1(net122),
    .A2(clknet_1_0__leaf_net482),
    .A3(net195),
    .S0(net616),
    .S1(clknet_1_1__leaf_net653),
    .X(net513));
 sky130_fd_sc_hd__mux4_1 c759 (.A0(net728),
    .A1(net800),
    .A2(net497),
    .A3(net760),
    .S0(clknet_1_0__leaf_net610),
    .S1(net719),
    .X(net514));
 sky130_fd_sc_hd__mux4_1 c760 (.A0(net92),
    .A1(net760),
    .A2(net979),
    .A3(net414),
    .S0(net508),
    .S1(net935),
    .X(net515));
 sky130_fd_sc_hd__mux4_1 c761 (.A0(net998),
    .A1(net1014),
    .A2(net514),
    .A3(net511),
    .S0(net907),
    .S1(net592),
    .X(net516));
 sky130_fd_sc_hd__mux4_1 c762 (.A0(net505),
    .A1(net973),
    .A2(net412),
    .A3(net515),
    .S0(net626),
    .S1(clknet_1_0__leaf_net673),
    .X(net517));
 sky130_fd_sc_hd__a41o_1 c763 (.A1(net947),
    .A2(net227),
    .A3(net592),
    .A4(clknet_1_1__leaf_net671),
    .B1(net722),
    .X(net518));
 sky130_fd_sc_hd__mux4_1 c764 (.A0(net490),
    .A1(net496),
    .A2(net394),
    .A3(net518),
    .S0(net601),
    .S1(net639),
    .X(net519));
 sky130_fd_sc_hd__dfrbp_1 merge765 (.CLK(clknet_4_14_0_clk),
    .D(net347),
    .Q(net348),
    .Q_N(net520));
 sky130_fd_sc_hd__dfrbp_1 merge766 (.CLK(clknet_4_15_0_clk),
    .D(net422),
    .RESET_B(net423),
    .Q(net523),
    .Q_N(net522));
 sky130_fd_sc_hd__xnor2_1 merge767 (.A(net352),
    .B(net358),
    .Y(net524));
 sky130_fd_sc_hd__xnor2_1 merge768 (.A(net519),
    .B(net504),
    .Y(net525));
 sky130_fd_sc_hd__xnor2_1 merge769 (.A(net287),
    .B(net288),
    .Y(net526));
 sky130_fd_sc_hd__dfrtn_1 merge770 (.CLK_N(clknet_4_3_0_clk),
    .D(net160),
    .RESET_B(net140),
    .Q(net527));
 sky130_fd_sc_hd__xnor2_1 merge771 (.A(net477),
    .B(net479),
    .Y(net528));
 sky130_fd_sc_hd__dfrtp_1 merge772 (.CLK(clknet_4_0_0_clk),
    .D(net91),
    .RESET_B(net94),
    .Q(net867));
 sky130_fd_sc_hd__dfrtp_4 merge773 (.CLK(clknet_4_11_0_clk),
    .D(net325),
    .RESET_B(net311),
    .Q(net529));
 sky130_fd_sc_hd__xnor2_1 merge774 (.A(net167),
    .B(net169),
    .Y(net530));
 sky130_fd_sc_hd__xnor2_1 merge775 (.A(net396),
    .B(net397),
    .Y(net531));
 sky130_fd_sc_hd__xnor2_1 merge776 (.A(net373),
    .B(net374),
    .Y(net532));
 sky130_fd_sc_hd__dfrtp_2 merge777 (.CLK(clknet_4_8_0_clk),
    .D(net137),
    .RESET_B(net131),
    .Q(net533));
 sky130_fd_sc_hd__xnor2_1 merge778 (.A(net485),
    .B(net486),
    .Y(net534));
 sky130_fd_sc_hd__dfsbp_1 merge779 (.CLK(clknet_4_9_0_clk),
    .D(net235),
    .SET_B(net236),
    .Q(net536),
    .Q_N(net535));
 sky130_fd_sc_hd__dfsbp_2 merge780 (.CLK(clknet_4_2_0_clk),
    .D(net55),
    .SET_B(net61),
    .Q(net538),
    .Q_N(net537));
 sky130_fd_sc_hd__dfstp_1 merge781 (.CLK(clknet_4_6_0_clk),
    .D(net244),
    .SET_B(net247),
    .Q(net539));
 sky130_fd_sc_hd__xnor2_1 merge782 (.A(net41),
    .B(net40),
    .Y(net540));
 sky130_fd_sc_hd__xnor2_1 merge783 (.A(net181),
    .B(net187),
    .Y(net541));
 sky130_fd_sc_hd__dfstp_1 merge784 (.CLK(clknet_4_15_0_clk),
    .D(net438),
    .SET_B(net439),
    .Q(net542));
 sky130_fd_sc_hd__dfstp_2 merge785 (.CLK(clknet_4_0_0_clk),
    .D(net82),
    .SET_B(net65),
    .Q(net543));
 sky130_fd_sc_hd__dlrbn_2 merge786 (.D(net216),
    .GATE_N(clknet_4_10_0_clk),
    .RESET_B(net204),
    .Q(net545),
    .Q_N(net544));
 sky130_fd_sc_hd__xnor2_1 merge787 (.A(net274),
    .B(net279),
    .Y(net546));
 sky130_fd_sc_hd__xnor2_1 merge788 (.A(net188),
    .B(net191),
    .Y(net547));
 sky130_fd_sc_hd__xnor2_1 merge789 (.A(net525),
    .B(net375),
    .Y(net548));
 sky130_fd_sc_hd__xnor2_1 merge790 (.A(net301),
    .B(net413),
    .Y(net549));
 sky130_fd_sc_hd__xnor2_1 merge791 (.A(net369),
    .B(net363),
    .Y(net550));
 sky130_fd_sc_hd__dlrbn_1 merge792 (.D(net157),
    .GATE_N(clknet_4_3_0_clk),
    .RESET_B(net154),
    .Q(net552),
    .Q_N(net551));
 sky130_fd_sc_hd__dlrbp_1 merge793 (.D(net265),
    .GATE(clknet_4_4_0_clk),
    .RESET_B(net280),
    .Q(net553),
    .Q_N(net825));
 sky130_fd_sc_hd__xnor2_1 merge794 (.A(net382),
    .B(net517),
    .Y(net554));
 sky130_fd_sc_hd__dlrbp_2 merge795 (.GATE(clknet_4_8_0_clk),
    .RESET_B(net540),
    .Q(net845),
    .Q_N(net42));
 sky130_fd_sc_hd__xnor2_1 merge796 (.A(net398),
    .B(net404),
    .Y(net556));
 sky130_fd_sc_hd__xnor2_1 merge797 (.A(net411),
    .B(net193),
    .Y(net557));
 sky130_fd_sc_hd__xnor2_1 merge798 (.A(net194),
    .B(net547),
    .Y(net558));
 sky130_fd_sc_hd__dlrtn_1 merge799 (.D(net51),
    .GATE_N(clknet_4_2_0_clk),
    .RESET_B(net62),
    .Q(net559));
 sky130_fd_sc_hd__xnor2_1 merge800 (.A(net248),
    .B(net258),
    .Y(net560));
 sky130_fd_sc_hd__dlrtn_4 merge801 (.D(net74),
    .GATE_N(clknet_4_0_0_clk),
    .RESET_B(net76),
    .Q(net880));
 sky130_fd_sc_hd__xnor2_1 merge802 (.A(net456),
    .B(net455),
    .Y(net561));
 sky130_fd_sc_hd__dlrtn_1 merge803 (.D(net99),
    .GATE_N(clknet_4_0_0_clk),
    .Q(net851));
 sky130_fd_sc_hd__xnor2_1 merge804 (.A(net388),
    .B(net500),
    .Y(net562));
 sky130_fd_sc_hd__dlrtp_1 merge805 (.D(net360),
    .GATE(clknet_4_13_0_clk),
    .RESET_B(net528),
    .Q(net563));
 sky130_fd_sc_hd__dlrtp_1 merge806 (.D(net134),
    .GATE(clknet_4_8_0_clk),
    .RESET_B(net135),
    .Q(net564));
 sky130_fd_sc_hd__xnor2_1 merge807 (.A(net513),
    .B(net516),
    .Y(net565));
 sky130_fd_sc_hd__xnor2_1 merge808 (.A(net299),
    .B(net289),
    .Y(net566));
 sky130_fd_sc_hd__dlrtp_2 merge809 (.D(net239),
    .GATE(clknet_4_11_0_clk),
    .RESET_B(net217),
    .Q(net567));
 sky130_fd_sc_hd__xnor2_1 merge810 (.A(net302),
    .B(net300),
    .Y(net568));
 sky130_fd_sc_hd__edfxbp_1 merge811 (.CLK(clknet_4_15_0_clk),
    .D(net449),
    .DE(net447),
    .Q(net570),
    .Q_N(net569));
 sky130_fd_sc_hd__edfxtp_1 merge812 (.CLK(clknet_4_0_0_clk),
    .D(net83),
    .DE(net97),
    .Q(net873));
 sky130_fd_sc_hd__sdlclkp_1 merge813 (.CLK(clknet_4_3_0_clk),
    .GATE(net142),
    .SCE(net172),
    .GCLK(net571));
 sky130_fd_sc_hd__xnor2_1 merge814 (.A(net387),
    .B(net512),
    .Y(net572));
 sky130_fd_sc_hd__xnor2_1 merge815 (.A(net297),
    .B(net298),
    .Y(net573));
 sky130_fd_sc_hd__xnor2_1 merge816 (.A(net383),
    .B(net384),
    .Y(net574));
 sky130_fd_sc_hd__xnor2_1 merge817 (.A(net185),
    .B(net541),
    .Y(net575));
 sky130_fd_sc_hd__xnor2_1 merge818 (.A(net493),
    .B(net499),
    .Y(net576));
 sky130_fd_sc_hd__sdlclkp_2 merge819 (.CLK(clknet_4_12_0_clk),
    .GATE(net344),
    .SCE(net330),
    .GCLK(net577));
 sky130_fd_sc_hd__sdlclkp_4 merge820 (.CLK(clknet_4_1_0_clk),
    .GATE(net100),
    .SCE(net77),
    .GCLK(net868));
 sky130_fd_sc_hd__xnor2_1 merge821 (.A(net407),
    .B(net506),
    .Y(net578));
 sky130_fd_sc_hd__dfrbp_2 merge822 (.CLK(clknet_4_5_0_clk),
    .D(net578),
    .RESET_B(net557),
    .Q(net824),
    .Q_N(net579));
 sky130_fd_sc_hd__dfrbp_1 merge823 (.CLK(clknet_4_13_0_clk),
    .D(net480),
    .RESET_B(net475),
    .Q(net581),
    .Q_N(net580));
 sky130_fd_sc_hd__dfrtn_1 merge824 (.CLK_N(clknet_4_3_0_clk),
    .D(net147),
    .RESET_B(net152),
    .Q(net865));
 sky130_fd_sc_hd__dfrtp_1 merge825 (.CLK(clknet_4_4_0_clk),
    .RESET_B(net558),
    .Q(net853));
 sky130_fd_sc_hd__xnor2_1 merge826 (.A(net565),
    .B(net507),
    .Y(net582));
 sky130_fd_sc_hd__xnor2_1 merge827 (.A(net491),
    .B(net488),
    .Y(net583));
 sky130_fd_sc_hd__dfrtp_2 merge828 (.CLK(clknet_4_5_0_clk),
    .D(net256),
    .RESET_B(net556),
    .Q(net584));
 sky130_fd_sc_hd__dfrtp_1 merge829 (.CLK(clknet_4_4_0_clk),
    .D(net546),
    .RESET_B(net568),
    .Q(net837));
 sky130_fd_sc_hd__dfsbp_2 merge830 (.CLK(clknet_4_2_0_clk),
    .D(net166),
    .SET_B(net165),
    .Q(net586),
    .Q_N(net585));
 sky130_fd_sc_hd__dfsbp_1 merge831 (.CLK(clknet_4_12_0_clk),
    .D(net550),
    .SET_B(net351),
    .Q(net588),
    .Q_N(net587));
 sky130_fd_sc_hd__dfstp_1 merge832 (.CLK(clknet_4_9_0_clk),
    .D(net251),
    .SET_B(net524),
    .Q(net589));
 sky130_fd_sc_hd__dfstp_4 merge833 (.CLK(clknet_4_1_0_clk),
    .D(net575),
    .SET_B(net190),
    .Q(net590));
 sky130_fd_sc_hd__dfstp_1 merge834 (.CLK(clknet_4_4_0_clk),
    .D(net566),
    .SET_B(net549),
    .Q(net869));
 sky130_fd_sc_hd__xnor2_1 merge835 (.A(net510),
    .B(net441),
    .Y(net591));
 sky130_fd_sc_hd__dlrbn_1 merge836 (.D(net271),
    .GATE_N(clknet_4_7_0_clk),
    .RESET_B(net582),
    .Q(net593),
    .Q_N(net592));
 sky130_fd_sc_hd__xnor2_1 merge837 (.A(net278),
    .B(net576),
    .Y(net594));
 sky130_fd_sc_hd__dlrbn_1 merge838 (.D(net257),
    .GATE_N(clknet_4_6_0_clk),
    .RESET_B(net548),
    .Q(net596),
    .Q_N(net595));
 sky130_fd_sc_hd__dlrbp_1 merge839 (.D(net442),
    .GATE(clknet_4_13_0_clk),
    .RESET_B(net350),
    .Q(net598),
    .Q_N(net597));
 sky130_fd_sc_hd__dlrbp_1 merge840 (.D(net379),
    .GATE(clknet_4_6_0_clk),
    .RESET_B(net531),
    .Q(net600),
    .Q_N(net599));
 sky130_fd_sc_hd__dlrtn_1 merge841 (.D(net554),
    .GATE_N(clknet_4_7_0_clk),
    .RESET_B(net534),
    .Q(net601));
 sky130_fd_sc_hd__dlrtn_1 merge842 (.D(net392),
    .GATE_N(clknet_4_7_0_clk),
    .RESET_B(net405),
    .Q(net602));
 sky130_fd_sc_hd__dlrtn_1 merge843 (.D(net573),
    .GATE_N(clknet_4_4_0_clk),
    .RESET_B(net526),
    .Q(net838));
 sky130_fd_sc_hd__dlrtp_1 merge844 (.D(net574),
    .GATE(clknet_4_12_0_clk),
    .RESET_B(net380),
    .Q(net603));
 sky130_fd_sc_hd__dlrtp_2 merge845 (.D(net530),
    .GATE(clknet_4_1_0_clk),
    .RESET_B(net175),
    .Q(net835));
 sky130_fd_sc_hd__dlrtp_1 merge846 (.D(net532),
    .GATE(clknet_4_5_0_clk),
    .RESET_B(net294),
    .Q(net604));
 sky130_fd_sc_hd__edfxbp_1 merge847 (.CLK(clknet_4_1_0_clk),
    .D(net179),
    .DE(net81),
    .Q(net606),
    .Q_N(net605));
 sky130_fd_sc_hd__edfxtp_1 merge848 (.CLK(clknet_4_4_0_clk),
    .D(net291),
    .DE(net295),
    .Q(net607));
 sky130_fd_sc_hd__sdlclkp_1 merge849 (.CLK(clknet_4_6_0_clk),
    .GATE(net560),
    .GCLK(net253));
 sky130_fd_sc_hd__sdlclkp_2 merge850 (.CLK(clknet_4_7_0_clk),
    .GATE(net562),
    .SCE(net583),
    .GCLK(net609));
 sky130_fd_sc_hd__sdlclkp_4 merge851 (.CLK(clknet_4_13_0_clk),
    .GATE(net572),
    .SCE(net495),
    .GCLK(net610));
 sky130_fd_sc_hd__dfrbp_2 merge852 (.CLK(clknet_4_5_0_clk),
    .D(net474),
    .RESET_B(net409),
    .Q(net612),
    .Q_N(net611));
 sky130_fd_sc_hd__dfrbp_2 merge853 (.CLK(clknet_4_4_0_clk),
    .D(net285),
    .RESET_B(net277),
    .Q(net614),
    .Q_N(net613));
 sky130_fd_sc_hd__dfrtn_1 merge854 (.CLK_N(clknet_4_6_0_clk),
    .D(net391),
    .RESET_B(net269),
    .Q(net615));
 sky130_fd_sc_hd__dfrtp_4 merge855 (.CLK(clknet_4_13_0_clk),
    .D(net591),
    .RESET_B(net481),
    .Q(net616));
 sky130_fd_sc_hd__dfrtp_4 merge856 (.CLK(clknet_4_3_0_clk),
    .D(net263),
    .RESET_B(net594),
    .Q(net617));
 sky130_fd_sc_hd__dfrtp_2 merge857 (.CLK(clknet_4_13_0_clk),
    .D(net461),
    .RESET_B(net561),
    .Q(net618));
 sky130_fd_sc_hd__dfsbp_2 merge858 (.CLK(clknet_4_5_0_clk),
    .D(net395),
    .SET_B(net378),
    .Q(net620),
    .Q_N(net619));
 sky130_fd_sc_hd__dfsbp_2 merge859 (.CLK(clknet_4_12_0_clk),
    .D(net425),
    .SET_B(net354),
    .Q(net622),
    .Q_N(net621));
 sky130_fd_sc_hd__dfxbp_2 s860 (.CLK(clknet_4_8_0_clk),
    .D(net39),
    .Q(net624),
    .Q_N(net623));
 sky130_fd_sc_hd__dfxbp_2 s861 (.CLK(clknet_4_2_0_clk),
    .D(net48),
    .Q(net626),
    .Q_N(net625));
 sky130_fd_sc_hd__dfxtp_2 s862 (.CLK(clknet_4_2_0_clk),
    .D(net58),
    .Q(net627));
 sky130_fd_sc_hd__dfxtp_4 s863 (.CLK(clknet_4_2_0_clk),
    .D(net63),
    .Q(net628));
 sky130_fd_sc_hd__dfxtp_2 s864 (.CLK(clknet_4_0_0_clk),
    .D(net72),
    .Q(net629));
 sky130_fd_sc_hd__dlclkp_1 s865 (.CLK(clknet_4_2_0_clk),
    .GATE(net73),
    .GCLK(net630));
 sky130_fd_sc_hd__dlclkp_2 s866 (.CLK(clknet_4_1_0_clk),
    .GATE(net80),
    .GCLK(net631));
 sky130_fd_sc_hd__dlclkp_4 s867 (.CLK(clknet_4_0_0_clk),
    .GATE(net90),
    .GCLK(net632));
 sky130_fd_sc_hd__dlxbn_1 s868 (.D(net95),
    .GATE_N(clknet_4_0_0_clk),
    .Q(net634),
    .Q_N(net633));
 sky130_fd_sc_hd__dlxbn_1 s869 (.D(net98),
    .GATE_N(clknet_4_0_0_clk),
    .Q(net636),
    .Q_N(net635));
 sky130_fd_sc_hd__dlxbp_1 s870 (.D(net119),
    .GATE(clknet_4_10_0_clk),
    .Q(net638),
    .Q_N(net637));
 sky130_fd_sc_hd__dlxtn_2 s871 (.D(net136),
    .GATE_N(clknet_4_8_0_clk),
    .Q(net639));
 sky130_fd_sc_hd__dlxtn_2 s872 (.D(net138),
    .GATE_N(clknet_4_8_0_clk),
    .Q(net640));
 sky130_fd_sc_hd__dlxtn_2 s873 (.D(net139),
    .GATE_N(clknet_4_2_0_clk),
    .Q(net641));
 sky130_fd_sc_hd__dlxtp_1 s874 (.D(net144),
    .GATE(clknet_4_8_0_clk),
    .Q(net642));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s875 (.D(net148),
    .SLEEP_B(clknet_4_3_0_clk),
    .Q(net643));
 sky130_fd_sc_hd__dfxbp_2 s876 (.CLK(clknet_4_8_0_clk),
    .D(net149),
    .Q(net645),
    .Q_N(net644));
 sky130_fd_sc_hd__dfxbp_2 s877 (.CLK(clknet_4_3_0_clk),
    .D(net151),
    .Q(net647),
    .Q_N(net646));
 sky130_fd_sc_hd__dfxtp_2 s878 (.CLK(clknet_4_3_0_clk),
    .D(net158),
    .Q(net648));
 sky130_fd_sc_hd__dfxtp_2 s879 (.CLK(clknet_4_3_0_clk),
    .D(net159),
    .Q(net649));
 sky130_fd_sc_hd__dfxtp_2 s880 (.CLK(clknet_4_1_0_clk),
    .D(net161),
    .Q(net650));
 sky130_fd_sc_hd__dlclkp_1 s881 (.CLK(clknet_4_3_0_clk),
    .GATE(net171),
    .GCLK(net651));
 sky130_fd_sc_hd__dlclkp_2 s882 (.CLK(clknet_4_4_0_clk),
    .GATE(net178),
    .GCLK(net652));
 sky130_fd_sc_hd__dlclkp_4 s883 (.CLK(clknet_4_1_0_clk),
    .GATE(net184),
    .GCLK(net653));
 sky130_fd_sc_hd__dlxbn_2 s884 (.D(net206),
    .GATE_N(clknet_4_11_0_clk),
    .Q(net655),
    .Q_N(net654));
 sky130_fd_sc_hd__dlxbn_2 s885 (.D(net207),
    .GATE_N(clknet_4_10_0_clk),
    .Q(net657),
    .Q_N(net656));
 sky130_fd_sc_hd__dlxbp_1 s886 (.D(net210),
    .GATE(clknet_4_10_0_clk),
    .Q(net659),
    .Q_N(net658));
 sky130_fd_sc_hd__dlxtn_2 s887 (.D(net224),
    .GATE_N(clknet_4_9_0_clk),
    .Q(net847));
 sky130_fd_sc_hd__dlxtn_4 s888 (.D(net226),
    .GATE_N(clknet_4_8_0_clk),
    .Q(net660));
 sky130_fd_sc_hd__dlxtn_4 s889 (.D(net228),
    .GATE_N(clknet_4_9_0_clk),
    .Q(net661));
 sky130_fd_sc_hd__dlxtp_1 s890 (.D(net232),
    .GATE(clknet_4_9_0_clk),
    .Q(net662));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s891 (.D(net234),
    .SLEEP_B(clknet_4_9_0_clk),
    .Q(net663));
 sky130_fd_sc_hd__dfxbp_2 s892 (.CLK(clknet_4_9_0_clk),
    .D(net237),
    .Q(net665),
    .Q_N(net664));
 sky130_fd_sc_hd__dfxbp_2 s893 (.CLK(clknet_4_3_0_clk),
    .D(net242),
    .Q(net667),
    .Q_N(net666));
 sky130_fd_sc_hd__dfxtp_1 s894 (.CLK(clknet_4_9_0_clk),
    .D(net245),
    .Q(net668));
 sky130_fd_sc_hd__dfxtp_1 s895 (.CLK(clknet_4_6_0_clk),
    .D(net254),
    .Q(net669));
 sky130_fd_sc_hd__dfxtp_1 s896 (.CLK(clknet_4_9_0_clk),
    .D(net255),
    .Q(net670));
 sky130_fd_sc_hd__dlclkp_1 s897 (.CLK(clknet_4_4_0_clk),
    .GATE(net267),
    .GCLK(net671));
 sky130_fd_sc_hd__dlclkp_2 s898 (.CLK(clknet_4_4_0_clk),
    .GATE(net286),
    .GCLK(net672));
 sky130_fd_sc_hd__dlclkp_4 s899 (.CLK(clknet_4_10_0_clk),
    .GATE(net305),
    .GCLK(net673));
 sky130_fd_sc_hd__dlxbn_2 s900 (.D(net306),
    .GATE_N(clknet_4_10_0_clk),
    .Q(net675),
    .Q_N(net674));
 sky130_fd_sc_hd__dlxbn_2 s901 (.D(net310),
    .GATE_N(clknet_4_11_0_clk),
    .Q(net677),
    .Q_N(net676));
 sky130_fd_sc_hd__dlxbp_1 s902 (.D(net312),
    .GATE(clknet_4_14_0_clk),
    .Q(net679),
    .Q_N(net678));
 sky130_fd_sc_hd__dlxtn_2 s903 (.D(net319),
    .GATE_N(clknet_4_14_0_clk),
    .Q(net680));
 sky130_fd_sc_hd__dlxtn_2 s904 (.D(net320),
    .GATE_N(clknet_4_14_0_clk),
    .Q(net681));
 sky130_fd_sc_hd__dlxtn_2 s905 (.D(net322),
    .GATE_N(clknet_4_11_0_clk),
    .Q(net682));
 sky130_fd_sc_hd__dlxtp_1 s906 (.D(net323),
    .GATE(clknet_4_11_0_clk),
    .Q(net683));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s907 (.D(net324),
    .SLEEP_B(clknet_4_14_0_clk),
    .Q(net684));
 sky130_fd_sc_hd__dfxbp_1 s908 (.CLK(clknet_4_9_0_clk),
    .D(net328),
    .Q(net686),
    .Q_N(net685));
 sky130_fd_sc_hd__dfxbp_1 s909 (.CLK(clknet_4_11_0_clk),
    .D(net329),
    .Q(net688),
    .Q_N(net687));
 sky130_fd_sc_hd__dfxtp_2 s910 (.CLK(clknet_4_14_0_clk),
    .D(net331),
    .Q(net689));
 sky130_fd_sc_hd__dfxtp_2 s911 (.CLK(clknet_4_9_0_clk),
    .D(net334),
    .Q(net690));
 sky130_fd_sc_hd__dfxtp_4 s912 (.CLK(clknet_4_14_0_clk),
    .D(net336),
    .Q(net831));
 sky130_fd_sc_hd__dlclkp_1 s913 (.CLK(clknet_4_12_0_clk),
    .GATE(net337),
    .GCLK(net691));
 sky130_fd_sc_hd__dlclkp_2 s914 (.CLK(clknet_4_14_0_clk),
    .GATE(net341),
    .GCLK(net692));
 sky130_fd_sc_hd__dlclkp_4 s915 (.CLK(clknet_4_14_0_clk),
    .GATE(net342),
    .GCLK(net693));
 sky130_fd_sc_hd__dlxbn_1 s916 (.D(net346),
    .GATE_N(clknet_4_12_0_clk),
    .Q(net695),
    .Q_N(net694));
 sky130_fd_sc_hd__dlxbn_1 s917 (.D(net356),
    .GATE_N(clknet_4_12_0_clk),
    .Q(net697),
    .Q_N(net696));
 sky130_fd_sc_hd__dlxbp_1 s918 (.D(net357),
    .GATE(clknet_4_12_0_clk),
    .Q(net699),
    .Q_N(net698));
 sky130_fd_sc_hd__dlxtn_1 s919 (.D(net365),
    .GATE_N(clknet_4_12_0_clk),
    .Q(net827));
 sky130_fd_sc_hd__dlxtn_1 s920 (.D(net366),
    .GATE_N(clknet_4_12_0_clk),
    .Q(net700));
 sky130_fd_sc_hd__dlxtn_1 s921 (.D(net370),
    .GATE_N(clknet_4_12_0_clk),
    .Q(net701));
 sky130_fd_sc_hd__dlxtp_1 s922 (.D(net372),
    .GATE(clknet_4_7_0_clk),
    .Q(net702));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s923 (.D(net377),
    .SLEEP_B(clknet_4_6_0_clk),
    .Q(net703));
 sky130_fd_sc_hd__dfxbp_1 s924 (.CLK(clknet_4_7_0_clk),
    .D(net390),
    .Q(net705),
    .Q_N(net704));
 sky130_fd_sc_hd__dfxbp_1 s925 (.CLK(clknet_4_14_0_clk),
    .D(net418),
    .Q(net707),
    .Q_N(net706));
 sky130_fd_sc_hd__dfxtp_4 s926 (.CLK(clknet_4_15_0_clk),
    .D(net427),
    .Q(net708));
 sky130_fd_sc_hd__dfxtp_4 s927 (.CLK(clknet_4_15_0_clk),
    .D(net430),
    .Q(net709));
 sky130_fd_sc_hd__dfxtp_2 s928 (.CLK(clknet_4_15_0_clk),
    .D(net431),
    .Q(net710));
 sky130_fd_sc_hd__dlclkp_1 s929 (.CLK(clknet_4_15_0_clk),
    .GATE(net432),
    .GCLK(net711));
 sky130_fd_sc_hd__dlclkp_2 s930 (.CLK(clknet_4_15_0_clk),
    .GATE(net433),
    .GCLK(net712));
 sky130_fd_sc_hd__dlclkp_4 s931 (.CLK(clknet_4_15_0_clk),
    .GATE(net434),
    .GCLK(net713));
 sky130_fd_sc_hd__dlxbn_1 s932 (.D(net436),
    .GATE_N(clknet_4_13_0_clk),
    .Q(net715),
    .Q_N(net714));
 sky130_fd_sc_hd__dlxbn_1 s933 (.D(net445),
    .GATE_N(clknet_4_15_0_clk),
    .Q(net717),
    .Q_N(net716));
 sky130_fd_sc_hd__dlxbp_1 s934 (.D(net446),
    .GATE(clknet_4_15_0_clk),
    .Q(net719),
    .Q_N(net718));
 sky130_fd_sc_hd__dlxtn_1 s935 (.D(net470),
    .GATE_N(clknet_4_13_0_clk),
    .Q(net720));
 sky130_fd_sc_hd__dlxtn_1 s936 (.D(net471),
    .GATE_N(clknet_4_13_0_clk),
    .Q(net721));
 sky130_fd_sc_hd__dlxtn_1 s937 (.D(net473),
    .GATE_N(clknet_4_12_0_clk),
    .Q(net722));
 sky130_fd_sc_hd__dlxtp_1 s938 (.D(net494),
    .GATE(clknet_4_13_0_clk),
    .Q(net723));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Right_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Right_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Right_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Right_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Right_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Right_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Right_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Right_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Right_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Right_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Right_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Right_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Right_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Right_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Right_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Right_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Right_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Right_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Right_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Right_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Right_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_161 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_162 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_163 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_164 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_165 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_166 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_167 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_168 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_169 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_170 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_171 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_172 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_173 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_174 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_175 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_176 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_177 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_178 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_179 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_180 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_181 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_182 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Left_183 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Left_184 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Left_185 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Left_186 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Left_187 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Left_188 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Left_189 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Left_190 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Left_191 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Left_192 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Left_193 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Left_194 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Left_195 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Left_196 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Left_197 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Left_198 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Left_199 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Left_200 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Left_201 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Left_202 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Left_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1347 ();
 sky130_fd_sc_hd__clkbuf_2 input1 (.A(in0),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_2 input2 (.A(in1),
    .X(net192));
 sky130_fd_sc_hd__buf_2 input3 (.A(in10),
    .X(net724));
 sky130_fd_sc_hd__buf_4 input4 (.A(in11),
    .X(net725));
 sky130_fd_sc_hd__buf_1 input5 (.A(in12),
    .X(net726));
 sky130_fd_sc_hd__clkbuf_4 input6 (.A(in13),
    .X(net727));
 sky130_fd_sc_hd__buf_12 input7 (.A(in14),
    .X(net728));
 sky130_fd_sc_hd__clkbuf_2 input8 (.A(in15),
    .X(net729));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(in16),
    .X(net730));
 sky130_fd_sc_hd__clkbuf_2 input10 (.A(in17),
    .X(net731));
 sky130_fd_sc_hd__buf_12 input11 (.A(in18),
    .X(net732));
 sky130_fd_sc_hd__buf_6 input12 (.A(in19),
    .X(net733));
 sky130_fd_sc_hd__clkbuf_2 input13 (.A(in2),
    .X(net734));
 sky130_fd_sc_hd__clkbuf_4 input14 (.A(in20),
    .X(net735));
 sky130_fd_sc_hd__buf_2 input15 (.A(in21),
    .X(net736));
 sky130_fd_sc_hd__clkbuf_8 input16 (.A(in22),
    .X(net737));
 sky130_fd_sc_hd__buf_4 input17 (.A(in23),
    .X(net738));
 sky130_fd_sc_hd__buf_2 input18 (.A(in24),
    .X(net739));
 sky130_fd_sc_hd__buf_4 input19 (.A(in25),
    .X(net740));
 sky130_fd_sc_hd__buf_4 input20 (.A(in26),
    .X(net741));
 sky130_fd_sc_hd__clkbuf_4 input21 (.A(in27),
    .X(net742));
 sky130_fd_sc_hd__clkbuf_4 input22 (.A(in28),
    .X(net743));
 sky130_fd_sc_hd__buf_4 input23 (.A(in29),
    .X(net744));
 sky130_fd_sc_hd__clkbuf_4 input24 (.A(in3),
    .X(net745));
 sky130_fd_sc_hd__clkbuf_4 input25 (.A(in30),
    .X(net746));
 sky130_fd_sc_hd__buf_2 input26 (.A(in31),
    .X(net747));
 sky130_fd_sc_hd__buf_4 input27 (.A(in32),
    .X(net748));
 sky130_fd_sc_hd__clkbuf_4 input28 (.A(in33),
    .X(net749));
 sky130_fd_sc_hd__clkbuf_4 input29 (.A(in34),
    .X(net750));
 sky130_fd_sc_hd__buf_2 input30 (.A(in35),
    .X(net751));
 sky130_fd_sc_hd__clkbuf_2 input31 (.A(in36),
    .X(net752));
 sky130_fd_sc_hd__buf_4 input32 (.A(in37),
    .X(net753));
 sky130_fd_sc_hd__buf_4 input33 (.A(in38),
    .X(net754));
 sky130_fd_sc_hd__buf_4 input34 (.A(in39),
    .X(net755));
 sky130_fd_sc_hd__clkbuf_4 input35 (.A(in4),
    .X(net756));
 sky130_fd_sc_hd__buf_4 input36 (.A(in40),
    .X(net757));
 sky130_fd_sc_hd__buf_2 input37 (.A(in41),
    .X(net758));
 sky130_fd_sc_hd__buf_2 input38 (.A(in42),
    .X(net759));
 sky130_fd_sc_hd__buf_4 input39 (.A(in43),
    .X(net760));
 sky130_fd_sc_hd__buf_4 input40 (.A(in44),
    .X(net761));
 sky130_fd_sc_hd__clkbuf_2 input41 (.A(in45),
    .X(net762));
 sky130_fd_sc_hd__dlymetal6s2s_1 input42 (.A(in46),
    .X(net763));
 sky130_fd_sc_hd__clkbuf_2 input43 (.A(in47),
    .X(net764));
 sky130_fd_sc_hd__buf_2 input44 (.A(in48),
    .X(net765));
 sky130_fd_sc_hd__clkbuf_1 input45 (.A(in49),
    .X(net766));
 sky130_fd_sc_hd__clkbuf_4 input46 (.A(in5),
    .X(net767));
 sky130_fd_sc_hd__buf_1 input47 (.A(in50),
    .X(net768));
 sky130_fd_sc_hd__buf_2 input48 (.A(in51),
    .X(net769));
 sky130_fd_sc_hd__buf_1 input49 (.A(in52),
    .X(net770));
 sky130_fd_sc_hd__clkbuf_4 input50 (.A(in53),
    .X(net771));
 sky130_fd_sc_hd__clkbuf_2 input51 (.A(in54),
    .X(net772));
 sky130_fd_sc_hd__clkbuf_2 input52 (.A(in55),
    .X(net773));
 sky130_fd_sc_hd__clkbuf_2 input53 (.A(in56),
    .X(net774));
 sky130_fd_sc_hd__clkbuf_2 input54 (.A(in57),
    .X(net775));
 sky130_fd_sc_hd__buf_4 input55 (.A(in58),
    .X(net776));
 sky130_fd_sc_hd__clkbuf_2 input56 (.A(in59),
    .X(net777));
 sky130_fd_sc_hd__clkbuf_2 input57 (.A(in6),
    .X(net778));
 sky130_fd_sc_hd__clkbuf_2 input58 (.A(in60),
    .X(net779));
 sky130_fd_sc_hd__buf_2 input59 (.A(in61),
    .X(net780));
 sky130_fd_sc_hd__buf_1 input60 (.A(in62),
    .X(net781));
 sky130_fd_sc_hd__buf_1 input61 (.A(in63),
    .X(net782));
 sky130_fd_sc_hd__clkbuf_1 input62 (.A(in64),
    .X(net783));
 sky130_fd_sc_hd__buf_1 input63 (.A(in65),
    .X(net784));
 sky130_fd_sc_hd__clkbuf_4 input64 (.A(in66),
    .X(net785));
 sky130_fd_sc_hd__buf_1 input65 (.A(in67),
    .X(net786));
 sky130_fd_sc_hd__buf_1 input66 (.A(in68),
    .X(net787));
 sky130_fd_sc_hd__buf_1 input67 (.A(in69),
    .X(net788));
 sky130_fd_sc_hd__clkbuf_2 input68 (.A(in7),
    .X(net789));
 sky130_fd_sc_hd__buf_1 input69 (.A(in70),
    .X(net790));
 sky130_fd_sc_hd__clkbuf_2 input70 (.A(in71),
    .X(net791));
 sky130_fd_sc_hd__clkbuf_1 input71 (.A(in72),
    .X(net792));
 sky130_fd_sc_hd__buf_1 input72 (.A(in73),
    .X(net793));
 sky130_fd_sc_hd__buf_1 input73 (.A(in74),
    .X(net794));
 sky130_fd_sc_hd__clkbuf_2 input74 (.A(in75),
    .X(net795));
 sky130_fd_sc_hd__buf_1 input75 (.A(in76),
    .X(net796));
 sky130_fd_sc_hd__clkbuf_1 input76 (.A(in77),
    .X(net797));
 sky130_fd_sc_hd__buf_1 input77 (.A(in78),
    .X(net798));
 sky130_fd_sc_hd__buf_1 input78 (.A(in79),
    .X(net799));
 sky130_fd_sc_hd__clkbuf_4 input79 (.A(in8),
    .X(net800));
 sky130_fd_sc_hd__clkbuf_4 input80 (.A(in80),
    .X(net801));
 sky130_fd_sc_hd__buf_2 input81 (.A(in81),
    .X(net802));
 sky130_fd_sc_hd__clkbuf_1 input82 (.A(in82),
    .X(net803));
 sky130_fd_sc_hd__buf_1 input83 (.A(in83),
    .X(net804));
 sky130_fd_sc_hd__dlymetal6s2s_1 input84 (.A(in84),
    .X(net805));
 sky130_fd_sc_hd__buf_1 input85 (.A(in85),
    .X(net806));
 sky130_fd_sc_hd__buf_1 input86 (.A(in86),
    .X(net807));
 sky130_fd_sc_hd__buf_1 input87 (.A(in87),
    .X(net808));
 sky130_fd_sc_hd__clkbuf_2 input88 (.A(in88),
    .X(net809));
 sky130_fd_sc_hd__buf_1 input89 (.A(in89),
    .X(net810));
 sky130_fd_sc_hd__buf_4 input90 (.A(in9),
    .X(net811));
 sky130_fd_sc_hd__buf_1 input91 (.A(in90),
    .X(net812));
 sky130_fd_sc_hd__buf_2 input92 (.A(in91),
    .X(net813));
 sky130_fd_sc_hd__buf_2 input93 (.A(in92),
    .X(net814));
 sky130_fd_sc_hd__dlymetal6s2s_1 input94 (.A(in93),
    .X(net815));
 sky130_fd_sc_hd__buf_1 input95 (.A(in94),
    .X(net816));
 sky130_fd_sc_hd__buf_2 input96 (.A(in95),
    .X(net817));
 sky130_fd_sc_hd__dlymetal6s2s_1 input97 (.A(in96),
    .X(net818));
 sky130_fd_sc_hd__buf_2 input98 (.A(in97),
    .X(net819));
 sky130_fd_sc_hd__clkbuf_2 input99 (.A(in98),
    .X(net820));
 sky130_fd_sc_hd__clkbuf_2 input100 (.A(in99),
    .X(net821));
 sky130_fd_sc_hd__clkbuf_4 output101 (.A(net933),
    .X(out0));
 sky130_fd_sc_hd__buf_2 output102 (.A(net823),
    .X(out10));
 sky130_fd_sc_hd__buf_2 output103 (.A(net824),
    .X(out11));
 sky130_fd_sc_hd__buf_2 output104 (.A(net825),
    .X(out12));
 sky130_fd_sc_hd__buf_2 output105 (.A(net826),
    .X(out13));
 sky130_fd_sc_hd__buf_2 output106 (.A(net827),
    .X(out14));
 sky130_fd_sc_hd__buf_2 output107 (.A(net828),
    .X(out15));
 sky130_fd_sc_hd__buf_2 output108 (.A(net829),
    .X(out18));
 sky130_fd_sc_hd__buf_2 output109 (.A(net830),
    .X(out19));
 sky130_fd_sc_hd__buf_2 output110 (.A(net831),
    .X(out2));
 sky130_fd_sc_hd__buf_2 output111 (.A(net832),
    .X(out21));
 sky130_fd_sc_hd__buf_2 output112 (.A(net833),
    .X(out23));
 sky130_fd_sc_hd__clkbuf_1 output113 (.A(clknet_1_1__leaf_net834),
    .X(out24));
 sky130_fd_sc_hd__buf_2 output114 (.A(net835),
    .X(out25));
 sky130_fd_sc_hd__clkbuf_1 output115 (.A(clknet_1_0__leaf_net836),
    .X(out27));
 sky130_fd_sc_hd__buf_2 output116 (.A(net837),
    .X(out3));
 sky130_fd_sc_hd__buf_2 output117 (.A(net838),
    .X(out30));
 sky130_fd_sc_hd__buf_2 output118 (.A(net928),
    .X(out31));
 sky130_fd_sc_hd__buf_2 output119 (.A(net840),
    .X(out32));
 sky130_fd_sc_hd__buf_2 output120 (.A(net841),
    .X(out33));
 sky130_fd_sc_hd__buf_2 output121 (.A(net842),
    .X(out34));
 sky130_fd_sc_hd__buf_2 output122 (.A(net903),
    .X(out35));
 sky130_fd_sc_hd__clkbuf_1 output123 (.A(clknet_1_0__leaf_net844),
    .X(out38));
 sky130_fd_sc_hd__buf_2 output124 (.A(net944),
    .X(out4));
 sky130_fd_sc_hd__buf_2 output125 (.A(net846),
    .X(out40));
 sky130_fd_sc_hd__clkbuf_4 output126 (.A(net847),
    .X(out41));
 sky130_fd_sc_hd__buf_2 output127 (.A(net848),
    .X(out42));
 sky130_fd_sc_hd__buf_2 output128 (.A(net849),
    .X(out43));
 sky130_fd_sc_hd__clkbuf_1 output129 (.A(net850),
    .X(out44));
 sky130_fd_sc_hd__clkbuf_1 output130 (.A(clknet_1_0__leaf_net851),
    .X(out47));
 sky130_fd_sc_hd__clkbuf_4 output131 (.A(net1055),
    .X(out5));
 sky130_fd_sc_hd__clkbuf_1 output132 (.A(clknet_1_0__leaf_net853),
    .X(out50));
 sky130_fd_sc_hd__buf_2 output133 (.A(net854),
    .X(out51));
 sky130_fd_sc_hd__clkbuf_1 output134 (.A(clknet_1_0__leaf_net855),
    .X(out52));
 sky130_fd_sc_hd__buf_2 output135 (.A(net856),
    .X(out53));
 sky130_fd_sc_hd__clkbuf_1 output136 (.A(net857),
    .X(out54));
 sky130_fd_sc_hd__buf_2 output137 (.A(net858),
    .X(out56));
 sky130_fd_sc_hd__buf_2 output138 (.A(net859),
    .X(out57));
 sky130_fd_sc_hd__clkbuf_1 output139 (.A(clknet_1_1__leaf_net860),
    .X(out58));
 sky130_fd_sc_hd__clkbuf_1 output140 (.A(net861),
    .X(out59));
 sky130_fd_sc_hd__clkbuf_4 output141 (.A(net918),
    .X(out6));
 sky130_fd_sc_hd__buf_2 output142 (.A(net863),
    .X(out60));
 sky130_fd_sc_hd__buf_2 output143 (.A(net864),
    .X(out61));
 sky130_fd_sc_hd__buf_2 output144 (.A(net865),
    .X(out64));
 sky130_fd_sc_hd__clkbuf_1 output145 (.A(clknet_1_0__leaf_net866),
    .X(out65));
 sky130_fd_sc_hd__buf_2 output146 (.A(net867),
    .X(out66));
 sky130_fd_sc_hd__clkbuf_1 output147 (.A(clknet_1_0__leaf_net868),
    .X(out68));
 sky130_fd_sc_hd__buf_2 output148 (.A(net869),
    .X(out7));
 sky130_fd_sc_hd__buf_2 output149 (.A(net870),
    .X(out70));
 sky130_fd_sc_hd__buf_2 output150 (.A(net871),
    .X(out72));
 sky130_fd_sc_hd__buf_2 output151 (.A(net872),
    .X(out74));
 sky130_fd_sc_hd__buf_2 output152 (.A(net873),
    .X(out76));
 sky130_fd_sc_hd__buf_2 output153 (.A(net1045),
    .X(out77));
 sky130_fd_sc_hd__clkbuf_1 output154 (.A(clknet_1_0__leaf_net875),
    .X(out78));
 sky130_fd_sc_hd__buf_2 output155 (.A(net876),
    .X(out79));
 sky130_fd_sc_hd__buf_2 output156 (.A(net877),
    .X(out81));
 sky130_fd_sc_hd__buf_2 output157 (.A(net878),
    .X(out82));
 sky130_fd_sc_hd__buf_2 output158 (.A(net879),
    .X(out83));
 sky130_fd_sc_hd__buf_2 output159 (.A(net880),
    .X(out86));
 sky130_fd_sc_hd__buf_2 output160 (.A(net881),
    .X(out87));
 sky130_fd_sc_hd__buf_2 output161 (.A(net882),
    .X(out88));
 sky130_fd_sc_hd__buf_2 output162 (.A(net883),
    .X(out89));
 sky130_fd_sc_hd__clkbuf_4 output163 (.A(net884),
    .X(out9));
 sky130_fd_sc_hd__buf_2 output164 (.A(net885),
    .X(out90));
 sky130_fd_sc_hd__buf_2 output165 (.A(net886),
    .X(out93));
 sky130_fd_sc_hd__buf_2 output166 (.A(net887),
    .X(out99));
 sky130_fd_sc_hd__buf_2 fanout167 (.A(net889),
    .X(net888));
 sky130_fd_sc_hd__buf_2 fanout168 (.A(net304),
    .X(net889));
 sky130_fd_sc_hd__clkbuf_4 fanout169 (.A(net891),
    .X(net890));
 sky130_fd_sc_hd__clkbuf_2 fanout170 (.A(net150),
    .X(net891));
 sky130_fd_sc_hd__clkbuf_4 fanout171 (.A(net893),
    .X(net892));
 sky130_fd_sc_hd__clkbuf_2 fanout172 (.A(net826),
    .X(net893));
 sky130_fd_sc_hd__clkbuf_4 fanout173 (.A(net205),
    .X(net894));
 sky130_fd_sc_hd__buf_4 fanout174 (.A(net114),
    .X(net895));
 sky130_fd_sc_hd__clkbuf_4 fanout175 (.A(net34),
    .X(net896));
 sky130_fd_sc_hd__clkbuf_4 fanout176 (.A(net126),
    .X(net897));
 sky130_fd_sc_hd__buf_4 fanout177 (.A(net30),
    .X(net898));
 sky130_fd_sc_hd__clkbuf_4 fanout178 (.A(net112),
    .X(net899));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout179 (.A(net112),
    .X(net900));
 sky130_fd_sc_hd__buf_8 fanout180 (.A(net31),
    .X(net901));
 sky130_fd_sc_hd__buf_4 fanout181 (.A(net843),
    .X(net902));
 sky130_fd_sc_hd__clkbuf_2 fanout182 (.A(net843),
    .X(net903));
 sky130_fd_sc_hd__clkbuf_4 fanout183 (.A(net47),
    .X(net904));
 sky130_fd_sc_hd__buf_12 fanout184 (.A(net22),
    .X(net905));
 sky130_fd_sc_hd__clkbuf_4 fanout185 (.A(net907),
    .X(net906));
 sky130_fd_sc_hd__buf_4 fanout186 (.A(net198),
    .X(net907));
 sky130_fd_sc_hd__buf_12 fanout187 (.A(net21),
    .X(net908));
 sky130_fd_sc_hd__buf_2 fanout188 (.A(net21),
    .X(net909));
 sky130_fd_sc_hd__buf_4 fanout189 (.A(net911),
    .X(net910));
 sky130_fd_sc_hd__buf_2 fanout190 (.A(net912),
    .X(net911));
 sky130_fd_sc_hd__buf_4 fanout191 (.A(net913),
    .X(net912));
 sky130_fd_sc_hd__buf_4 fanout192 (.A(net107),
    .X(net913));
 sky130_fd_sc_hd__clkbuf_4 fanout193 (.A(net105),
    .X(net914));
 sky130_fd_sc_hd__buf_12 fanout194 (.A(net20),
    .X(net915));
 sky130_fd_sc_hd__clkbuf_4 fanout195 (.A(net918),
    .X(net916));
 sky130_fd_sc_hd__buf_1 fanout196 (.A(net918),
    .X(net917));
 sky130_fd_sc_hd__buf_4 fanout197 (.A(net919),
    .X(net918));
 sky130_fd_sc_hd__buf_2 fanout198 (.A(net862),
    .X(net919));
 sky130_fd_sc_hd__buf_12 fanout199 (.A(net921),
    .X(net920));
 sky130_fd_sc_hd__buf_12 fanout200 (.A(net922),
    .X(net921));
 sky130_fd_sc_hd__buf_12 fanout201 (.A(net18),
    .X(net922));
 sky130_fd_sc_hd__clkbuf_4 fanout202 (.A(net16),
    .X(net923));
 sky130_fd_sc_hd__buf_8 fanout203 (.A(net14),
    .X(net924));
 sky130_fd_sc_hd__clkbuf_4 fanout204 (.A(net17),
    .X(net925));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout205 (.A(net17),
    .X(net926));
 sky130_fd_sc_hd__buf_12 fanout206 (.A(net13),
    .X(net927));
 sky130_fd_sc_hd__clkbuf_4 fanout207 (.A(net839),
    .X(net928));
 sky130_fd_sc_hd__buf_2 fanout208 (.A(net27),
    .X(net929));
 sky130_fd_sc_hd__buf_12 fanout209 (.A(net872),
    .X(net930));
 sky130_fd_sc_hd__buf_4 fanout210 (.A(net10),
    .X(net931));
 sky130_fd_sc_hd__buf_12 fanout211 (.A(net822),
    .X(net932));
 sky130_fd_sc_hd__buf_2 fanout212 (.A(net822),
    .X(net933));
 sky130_fd_sc_hd__clkbuf_4 fanout213 (.A(net935),
    .X(net934));
 sky130_fd_sc_hd__clkbuf_4 fanout214 (.A(net103),
    .X(net935));
 sky130_fd_sc_hd__buf_4 fanout215 (.A(net25),
    .X(net936));
 sky130_fd_sc_hd__buf_12 fanout216 (.A(net8),
    .X(net937));
 sky130_fd_sc_hd__buf_4 max_cap217 (.A(net662),
    .X(net938));
 sky130_fd_sc_hd__clkbuf_2 max_cap218 (.A(net642),
    .X(net939));
 sky130_fd_sc_hd__buf_4 fanout219 (.A(net639),
    .X(net940));
 sky130_fd_sc_hd__buf_2 max_cap220 (.A(net638),
    .X(net941));
 sky130_fd_sc_hd__buf_4 fanout221 (.A(net564),
    .X(net942));
 sky130_fd_sc_hd__clkbuf_4 fanout222 (.A(net559),
    .X(net943));
 sky130_fd_sc_hd__clkbuf_8 fanout223 (.A(net845),
    .X(net944));
 sky130_fd_sc_hd__buf_4 fanout224 (.A(net533),
    .X(net945));
 sky130_fd_sc_hd__buf_2 fanout225 (.A(net199),
    .X(net946));
 sky130_fd_sc_hd__buf_4 fanout226 (.A(net200),
    .X(net947));
 sky130_fd_sc_hd__buf_12 fanout227 (.A(net6),
    .X(net948));
 sky130_fd_sc_hd__clkbuf_4 fanout228 (.A(net950),
    .X(net949));
 sky130_fd_sc_hd__buf_12 fanout229 (.A(net811),
    .X(net950));
 sky130_fd_sc_hd__buf_4 fanout230 (.A(net811),
    .X(net951));
 sky130_fd_sc_hd__buf_4 fanout231 (.A(net954),
    .X(net952));
 sky130_fd_sc_hd__buf_4 fanout232 (.A(net954),
    .X(net953));
 sky130_fd_sc_hd__buf_4 fanout233 (.A(net730),
    .X(net954));
 sky130_fd_sc_hd__buf_4 fanout234 (.A(net729),
    .X(net955));
 sky130_fd_sc_hd__buf_4 fanout235 (.A(net800),
    .X(net956));
 sky130_fd_sc_hd__clkbuf_4 fanout236 (.A(net799),
    .X(net957));
 sky130_fd_sc_hd__clkbuf_4 fanout237 (.A(net791),
    .X(net958));
 sky130_fd_sc_hd__buf_12 fanout238 (.A(net728),
    .X(net959));
 sky130_fd_sc_hd__buf_4 fanout239 (.A(net789),
    .X(net960));
 sky130_fd_sc_hd__buf_4 fanout240 (.A(net778),
    .X(net961));
 sky130_fd_sc_hd__buf_4 fanout241 (.A(net777),
    .X(net962));
 sky130_fd_sc_hd__buf_4 fanout242 (.A(net774),
    .X(net963));
 sky130_fd_sc_hd__buf_4 fanout243 (.A(net726),
    .X(net964));
 sky130_fd_sc_hd__clkbuf_4 fanout244 (.A(net966),
    .X(net965));
 sky130_fd_sc_hd__clkbuf_4 fanout245 (.A(net967),
    .X(net966));
 sky130_fd_sc_hd__buf_12 fanout246 (.A(net767),
    .X(net967));
 sky130_fd_sc_hd__buf_4 fanout247 (.A(net724),
    .X(net968));
 sky130_fd_sc_hd__buf_4 fanout248 (.A(net192),
    .X(net969));
 sky130_fd_sc_hd__buf_4 fanout249 (.A(net739),
    .X(net970));
 sky130_fd_sc_hd__clkbuf_4 fanout250 (.A(net736),
    .X(net971));
 sky130_fd_sc_hd__clkbuf_8 fanout251 (.A(net734),
    .X(net972));
 sky130_fd_sc_hd__clkbuf_2 fanout252 (.A(net734),
    .X(net973));
 sky130_fd_sc_hd__buf_12 fanout253 (.A(net733),
    .X(net974));
 sky130_fd_sc_hd__buf_2 fanout254 (.A(net733),
    .X(net975));
 sky130_fd_sc_hd__clkbuf_4 fanout255 (.A(net977),
    .X(net976));
 sky130_fd_sc_hd__buf_12 fanout256 (.A(net978),
    .X(net977));
 sky130_fd_sc_hd__buf_12 fanout257 (.A(net732),
    .X(net978));
 sky130_fd_sc_hd__buf_4 fanout258 (.A(net731),
    .X(net979));
 sky130_fd_sc_hd__buf_4 fanout259 (.A(net101),
    .X(net980));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net713 (.A(net713),
    .X(clknet_0_net713));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net713 (.A(clknet_0_net713),
    .X(clknet_1_0__leaf_net713));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net713 (.A(clknet_0_net713),
    .X(clknet_1_1__leaf_net713));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net712 (.A(net712),
    .X(clknet_0_net712));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net712 (.A(clknet_0_net712),
    .X(clknet_1_0__leaf_net712));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net712 (.A(clknet_0_net712),
    .X(clknet_1_1__leaf_net712));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net711 (.A(net711),
    .X(clknet_0_net711));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net711 (.A(clknet_0_net711),
    .X(clknet_1_0__leaf_net711));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net711 (.A(clknet_0_net711),
    .X(clknet_1_1__leaf_net711));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net458 (.A(net458),
    .X(clknet_0_net458));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net458 (.A(clknet_0_net458),
    .X(clknet_1_0__leaf_net458));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net458 (.A(clknet_0_net458),
    .X(clknet_1_1__leaf_net458));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net482 (.A(net482),
    .X(clknet_0_net482));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net482 (.A(clknet_0_net482),
    .X(clknet_1_0__leaf_net482));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net482 (.A(clknet_0_net482),
    .X(clknet_1_1__leaf_net482));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net609 (.A(net609),
    .X(clknet_0_net609));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net609 (.A(clknet_0_net609),
    .X(clknet_1_0__leaf_net609));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net609 (.A(clknet_0_net609),
    .X(clknet_1_1__leaf_net609));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net483 (.A(net483),
    .X(clknet_0_net483));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net483 (.A(clknet_0_net483),
    .X(clknet_1_0__leaf_net483));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net483 (.A(clknet_0_net483),
    .X(clknet_1_1__leaf_net483));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net452 (.A(net452),
    .X(clknet_0_net452));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net452 (.A(clknet_0_net452),
    .X(clknet_1_0__leaf_net452));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net452 (.A(clknet_0_net452),
    .X(clknet_1_1__leaf_net452));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net457 (.A(net457),
    .X(clknet_0_net457));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net457 (.A(clknet_0_net457),
    .X(clknet_1_0__leaf_net457));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net457 (.A(clknet_0_net457),
    .X(clknet_1_1__leaf_net457));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net437 (.A(net437),
    .X(clknet_0_net437));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net437 (.A(clknet_0_net437),
    .X(clknet_1_0__leaf_net437));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net437 (.A(clknet_0_net437),
    .X(clknet_1_1__leaf_net437));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net454 (.A(net454),
    .X(clknet_0_net454));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net454 (.A(clknet_0_net454),
    .X(clknet_1_0__leaf_net454));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net454 (.A(clknet_0_net454),
    .X(clknet_1_1__leaf_net454));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net450 (.A(net450),
    .X(clknet_0_net450));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net450 (.A(clknet_0_net450),
    .X(clknet_1_0__leaf_net450));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net450 (.A(clknet_0_net450),
    .X(clknet_1_1__leaf_net450));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net444 (.A(net444),
    .X(clknet_0_net444));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net444 (.A(clknet_0_net444),
    .X(clknet_1_0__leaf_net444));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net444 (.A(clknet_0_net444),
    .X(clknet_1_1__leaf_net444));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net435 (.A(net435),
    .X(clknet_0_net435));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net435 (.A(clknet_0_net435),
    .X(clknet_1_0__leaf_net435));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net435 (.A(clknet_0_net435),
    .X(clknet_1_1__leaf_net435));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net451 (.A(net451),
    .X(clknet_0_net451));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net451 (.A(clknet_0_net451),
    .X(clknet_1_0__leaf_net451));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net451 (.A(clknet_0_net451),
    .X(clknet_1_1__leaf_net451));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net693 (.A(net693),
    .X(clknet_0_net693));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net693 (.A(clknet_0_net693),
    .X(clknet_1_0__leaf_net693));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net693 (.A(clknet_0_net693),
    .X(clknet_1_1__leaf_net693));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net345 (.A(net345),
    .X(clknet_0_net345));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net345 (.A(clknet_0_net345),
    .X(clknet_1_0__leaf_net345));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net345 (.A(clknet_0_net345),
    .X(clknet_1_1__leaf_net345));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net577 (.A(net577),
    .X(clknet_0_net577));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net577 (.A(clknet_0_net577),
    .X(clknet_1_0__leaf_net577));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net577 (.A(clknet_0_net577),
    .X(clknet_1_1__leaf_net577));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net466 (.A(net466),
    .X(clknet_0_net466));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net466 (.A(clknet_0_net466),
    .X(clknet_1_0__leaf_net466));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net466 (.A(clknet_0_net466),
    .X(clknet_1_1__leaf_net466));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net338 (.A(net338),
    .X(clknet_0_net338));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net338 (.A(clknet_0_net338),
    .X(clknet_1_0__leaf_net338));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net338 (.A(clknet_0_net338),
    .X(clknet_1_1__leaf_net338));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net343 (.A(net343),
    .X(clknet_0_net343));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net343 (.A(clknet_0_net343),
    .X(clknet_1_0__leaf_net343));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net343 (.A(clknet_0_net343),
    .X(clknet_1_1__leaf_net343));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net692 (.A(net692),
    .X(clknet_0_net692));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net692 (.A(clknet_0_net692),
    .X(clknet_1_0__leaf_net692));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net692 (.A(clknet_0_net692),
    .X(clknet_1_1__leaf_net692));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net691 (.A(net691),
    .X(clknet_0_net691));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net691 (.A(clknet_0_net691),
    .X(clknet_1_0__leaf_net691));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net691 (.A(clknet_0_net691),
    .X(clknet_1_1__leaf_net691));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net673 (.A(net673),
    .X(clknet_0_net673));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net673 (.A(clknet_0_net673),
    .X(clknet_1_0__leaf_net673));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net673 (.A(clknet_0_net673),
    .X(clknet_1_1__leaf_net673));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net463 (.A(net463),
    .X(clknet_0_net463));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net463 (.A(clknet_0_net463),
    .X(clknet_1_0__leaf_net463));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net463 (.A(clknet_0_net463),
    .X(clknet_1_1__leaf_net463));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net426 (.A(net426),
    .X(clknet_0_net426));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net426 (.A(clknet_0_net426),
    .X(clknet_1_0__leaf_net426));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net426 (.A(clknet_0_net426),
    .X(clknet_1_1__leaf_net426));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net428 (.A(net428),
    .X(clknet_0_net428));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net428 (.A(clknet_0_net428),
    .X(clknet_1_0__leaf_net428));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net428 (.A(clknet_0_net428),
    .X(clknet_1_1__leaf_net428));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net429 (.A(net429),
    .X(clknet_0_net429));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net429 (.A(clknet_0_net429),
    .X(clknet_1_0__leaf_net429));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net429 (.A(clknet_0_net429),
    .X(clknet_1_1__leaf_net429));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net316 (.A(net316),
    .X(clknet_0_net316));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net316 (.A(clknet_0_net316),
    .X(clknet_1_0__leaf_net316));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net316 (.A(clknet_0_net316),
    .X(clknet_1_1__leaf_net316));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net448 (.A(net448),
    .X(clknet_0_net448));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net448 (.A(clknet_0_net448),
    .X(clknet_1_0__leaf_net448));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net448 (.A(clknet_0_net448),
    .X(clknet_1_1__leaf_net448));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net610 (.A(net610),
    .X(clknet_0_net610));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net610 (.A(clknet_0_net610),
    .X(clknet_1_0__leaf_net610));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net610 (.A(clknet_0_net610),
    .X(clknet_1_1__leaf_net610));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net318 (.A(net318),
    .X(clknet_0_net318));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net318 (.A(clknet_0_net318),
    .X(clknet_1_0__leaf_net318));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net318 (.A(clknet_0_net318),
    .X(clknet_1_1__leaf_net318));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net440 (.A(net440),
    .X(clknet_0_net440));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net440 (.A(clknet_0_net440),
    .X(clknet_1_0__leaf_net440));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net440 (.A(clknet_0_net440),
    .X(clknet_1_1__leaf_net440));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net321 (.A(net321),
    .X(clknet_0_net321));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net321 (.A(clknet_0_net321),
    .X(clknet_1_0__leaf_net321));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net321 (.A(clknet_0_net321),
    .X(clknet_1_1__leaf_net321));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net315 (.A(net315),
    .X(clknet_0_net315));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net315 (.A(clknet_0_net315),
    .X(clknet_1_0__leaf_net315));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net315 (.A(clknet_0_net315),
    .X(clknet_1_1__leaf_net315));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net400 (.A(net400),
    .X(clknet_0_net400));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net400 (.A(clknet_0_net400),
    .X(clknet_1_0__leaf_net400));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net400 (.A(clknet_0_net400),
    .X(clknet_1_1__leaf_net400));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net349 (.A(net349),
    .X(clknet_0_net349));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net349 (.A(clknet_0_net349),
    .X(clknet_1_0__leaf_net349));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net349 (.A(clknet_0_net349),
    .X(clknet_1_1__leaf_net349));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net317 (.A(net317),
    .X(clknet_0_net317));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net317 (.A(clknet_0_net317),
    .X(clknet_1_0__leaf_net317));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net317 (.A(clknet_0_net317),
    .X(clknet_1_1__leaf_net317));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net367 (.A(net367),
    .X(clknet_0_net367));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net367 (.A(clknet_0_net367),
    .X(clknet_1_0__leaf_net367));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net367 (.A(clknet_0_net367),
    .X(clknet_1_1__leaf_net367));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net492 (.A(net492),
    .X(clknet_0_net492));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net492 (.A(clknet_0_net492),
    .X(clknet_1_0__leaf_net492));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net492 (.A(clknet_0_net492),
    .X(clknet_1_1__leaf_net492));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net672 (.A(net672),
    .X(clknet_0_net672));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net672 (.A(clknet_0_net672),
    .X(clknet_1_0__leaf_net672));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net672 (.A(clknet_0_net672),
    .X(clknet_1_1__leaf_net672));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net290 (.A(net290),
    .X(clknet_0_net290));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net290 (.A(clknet_0_net290),
    .X(clknet_1_0__leaf_net290));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net290 (.A(clknet_0_net290),
    .X(clknet_1_1__leaf_net290));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net671 (.A(net671),
    .X(clknet_0_net671));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net671 (.A(clknet_0_net671),
    .X(clknet_1_0__leaf_net671));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net671 (.A(clknet_0_net671),
    .X(clknet_1_1__leaf_net671));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net276 (.A(net276),
    .X(clknet_0_net276));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net276 (.A(clknet_0_net276),
    .X(clknet_1_0__leaf_net276));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net276 (.A(clknet_0_net276),
    .X(clknet_1_1__leaf_net276));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net653 (.A(net653),
    .X(clknet_0_net653));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net653 (.A(clknet_0_net653),
    .X(clknet_1_0__leaf_net653));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net653 (.A(clknet_0_net653),
    .X(clknet_1_1__leaf_net653));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net296 (.A(net296),
    .X(clknet_0_net296));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net296 (.A(clknet_0_net296),
    .X(clknet_1_0__leaf_net296));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net296 (.A(clknet_0_net296),
    .X(clknet_1_1__leaf_net296));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net292 (.A(net292),
    .X(clknet_0_net292));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net292 (.A(clknet_0_net292),
    .X(clknet_1_0__leaf_net292));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net292 (.A(clknet_0_net292),
    .X(clknet_1_1__leaf_net292));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net652 (.A(net652),
    .X(clknet_0_net652));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net652 (.A(clknet_0_net652),
    .X(clknet_1_0__leaf_net652));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net652 (.A(clknet_0_net652),
    .X(clknet_1_1__leaf_net652));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net866 (.A(net866),
    .X(clknet_0_net866));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net866 (.A(clknet_0_net866),
    .X(clknet_1_0__leaf_net866));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net866 (.A(clknet_0_net866),
    .X(clknet_1_1__leaf_net866));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net860 (.A(net860),
    .X(clknet_0_net860));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net860 (.A(clknet_0_net860),
    .X(clknet_1_0__leaf_net860));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net860 (.A(clknet_0_net860),
    .X(clknet_1_1__leaf_net860));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net853 (.A(net853),
    .X(clknet_0_net853));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net853 (.A(clknet_0_net853),
    .X(clknet_1_0__leaf_net853));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net853 (.A(clknet_0_net853),
    .X(clknet_1_1__leaf_net853));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net651 (.A(net651),
    .X(clknet_0_net651));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net651 (.A(clknet_0_net651),
    .X(clknet_1_0__leaf_net651));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net651 (.A(clknet_0_net651),
    .X(clknet_1_1__leaf_net651));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net177 (.A(net177),
    .X(clknet_0_net177));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net177 (.A(clknet_0_net177),
    .X(clknet_1_0__leaf_net177));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net177 (.A(clknet_0_net177),
    .X(clknet_1_1__leaf_net177));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net385 (.A(net385),
    .X(clknet_0_net385));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net385 (.A(clknet_0_net385),
    .X(clknet_1_0__leaf_net385));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net385 (.A(clknet_0_net385),
    .X(clknet_1_1__leaf_net385));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net176 (.A(net176),
    .X(clknet_0_net176));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net176 (.A(clknet_0_net176),
    .X(clknet_1_0__leaf_net176));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net176 (.A(clknet_0_net176),
    .X(clknet_1_1__leaf_net176));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net836 (.A(net836),
    .X(clknet_0_net836));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net836 (.A(clknet_0_net836),
    .X(clknet_1_0__leaf_net836));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net836 (.A(clknet_0_net836),
    .X(clknet_1_1__leaf_net836));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net281 (.A(net281),
    .X(clknet_0_net281));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net281 (.A(clknet_0_net281),
    .X(clknet_1_0__leaf_net281));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net281 (.A(clknet_0_net281),
    .X(clknet_1_1__leaf_net281));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net174 (.A(net174),
    .X(clknet_0_net174));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net174 (.A(clknet_0_net174),
    .X(clknet_1_0__leaf_net174));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net174 (.A(clknet_0_net174),
    .X(clknet_1_1__leaf_net174));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net371 (.A(net371),
    .X(clknet_0_net371));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net371 (.A(clknet_0_net371),
    .X(clknet_1_0__leaf_net371));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net371 (.A(clknet_0_net371),
    .X(clknet_1_1__leaf_net371));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net386 (.A(net386),
    .X(clknet_0_net386));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net386 (.A(clknet_0_net386),
    .X(clknet_1_0__leaf_net386));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net386 (.A(clknet_0_net386),
    .X(clknet_1_1__leaf_net386));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net173 (.A(net173),
    .X(clknet_0_net173));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net173 (.A(clknet_0_net173),
    .X(clknet_1_0__leaf_net173));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net173 (.A(clknet_0_net173),
    .X(clknet_1_1__leaf_net173));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net571 (.A(net571),
    .X(clknet_0_net571));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net571 (.A(clknet_0_net571),
    .X(clknet_1_0__leaf_net571));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net571 (.A(clknet_0_net571),
    .X(clknet_1_1__leaf_net571));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net189 (.A(net189),
    .X(clknet_0_net189));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net189 (.A(clknet_0_net189),
    .X(clknet_1_0__leaf_net189));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net189 (.A(clknet_0_net189),
    .X(clknet_1_1__leaf_net189));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net180 (.A(net180),
    .X(clknet_0_net180));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net180 (.A(clknet_0_net180),
    .X(clknet_1_0__leaf_net180));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net180 (.A(clknet_0_net180),
    .X(clknet_1_1__leaf_net180));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net155 (.A(net155),
    .X(clknet_0_net155));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net155 (.A(clknet_0_net155),
    .X(clknet_1_0__leaf_net155));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net155 (.A(clknet_0_net155),
    .X(clknet_1_1__leaf_net155));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net459 (.A(net459),
    .X(clknet_0_net459));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net459 (.A(clknet_0_net459),
    .X(clknet_1_0__leaf_net459));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net459 (.A(clknet_0_net459),
    .X(clknet_1_1__leaf_net459));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net250 (.A(net250),
    .X(clknet_0_net250));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net250 (.A(clknet_0_net250),
    .X(clknet_1_0__leaf_net250));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net250 (.A(clknet_0_net250),
    .X(clknet_1_1__leaf_net250));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net359 (.A(net359),
    .X(clknet_0_net359));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net359 (.A(clknet_0_net359),
    .X(clknet_1_0__leaf_net359));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net359 (.A(clknet_0_net359),
    .X(clknet_1_1__leaf_net359));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net355 (.A(net355),
    .X(clknet_0_net355));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net355 (.A(clknet_0_net355),
    .X(clknet_1_0__leaf_net355));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net355 (.A(clknet_0_net355),
    .X(clknet_1_1__leaf_net355));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net855 (.A(net855),
    .X(clknet_0_net855));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net855 (.A(clknet_0_net855),
    .X(clknet_1_0__leaf_net855));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net855 (.A(clknet_0_net855),
    .X(clknet_1_1__leaf_net855));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net632 (.A(net632),
    .X(clknet_0_net632));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net632 (.A(clknet_0_net632),
    .X(clknet_1_0__leaf_net632));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net632 (.A(clknet_0_net632),
    .X(clknet_1_1__leaf_net632));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net96 (.A(net96),
    .X(clknet_0_net96));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net96 (.A(clknet_0_net96),
    .X(clknet_1_0__leaf_net96));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net96 (.A(clknet_0_net96),
    .X(clknet_1_1__leaf_net96));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net868 (.A(net868),
    .X(clknet_0_net868));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net868 (.A(clknet_0_net868),
    .X(clknet_1_0__leaf_net868));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net868 (.A(clknet_0_net868),
    .X(clknet_1_1__leaf_net868));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net631 (.A(net631),
    .X(clknet_0_net631));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net631 (.A(clknet_0_net631),
    .X(clknet_1_0__leaf_net631));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net631 (.A(clknet_0_net631),
    .X(clknet_1_1__leaf_net631));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net875 (.A(net875),
    .X(clknet_0_net875));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net875 (.A(clknet_0_net875),
    .X(clknet_1_0__leaf_net875));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net875 (.A(clknet_0_net875),
    .X(clknet_1_1__leaf_net875));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net851 (.A(net851),
    .X(clknet_0_net851));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net851 (.A(clknet_0_net851),
    .X(clknet_1_0__leaf_net851));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net851 (.A(clknet_0_net851),
    .X(clknet_1_1__leaf_net851));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net84 (.A(net84),
    .X(clknet_0_net84));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net84 (.A(clknet_0_net84),
    .X(clknet_1_0__leaf_net84));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net84 (.A(clknet_0_net84),
    .X(clknet_1_1__leaf_net84));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net183 (.A(net183),
    .X(clknet_0_net183));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net183 (.A(clknet_0_net183),
    .X(clknet_1_0__leaf_net183));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net183 (.A(clknet_0_net183),
    .X(clknet_1_1__leaf_net183));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net834 (.A(net834),
    .X(clknet_0_net834));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net834 (.A(clknet_0_net834),
    .X(clknet_1_0__leaf_net834));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net834 (.A(clknet_0_net834),
    .X(clknet_1_1__leaf_net834));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net86 (.A(net86),
    .X(clknet_0_net86));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net86 (.A(clknet_0_net86),
    .X(clknet_1_0__leaf_net86));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net86 (.A(clknet_0_net86),
    .X(clknet_1_1__leaf_net86));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net78 (.A(net78),
    .X(clknet_0_net78));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net78 (.A(clknet_0_net78),
    .X(clknet_1_0__leaf_net78));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net78 (.A(clknet_0_net78),
    .X(clknet_1_1__leaf_net78));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net93 (.A(net93),
    .X(clknet_0_net93));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net93 (.A(clknet_0_net93),
    .X(clknet_1_0__leaf_net93));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net93 (.A(clknet_0_net93),
    .X(clknet_1_1__leaf_net93));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net630 (.A(net630),
    .X(clknet_0_net630));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net630 (.A(clknet_0_net630),
    .X(clknet_1_0__leaf_net630));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net630 (.A(clknet_0_net630),
    .X(clknet_1_1__leaf_net630));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net389 (.A(net389),
    .X(clknet_0_net389));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net389 (.A(clknet_0_net389),
    .X(clknet_1_0__leaf_net389));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net389 (.A(clknet_0_net389),
    .X(clknet_1_1__leaf_net389));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net844 (.A(net844),
    .X(clknet_0_net844));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net844 (.A(clknet_0_net844),
    .X(clknet_1_0__leaf_net844));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net844 (.A(clknet_0_net844),
    .X(clknet_1_1__leaf_net844));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer1 (.A(net22),
    .X(net981));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer2 (.A(net981),
    .X(net982));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer3 (.A(net260),
    .X(net983));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer4 (.A(net983),
    .X(net984));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer5 (.A(net984),
    .X(net985));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer6 (.A(net260),
    .X(net986));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer7 (.A(net24),
    .X(net987));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer8 (.A(net1065),
    .X(net988));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer9 (.A(net988),
    .X(net989));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer10 (.A(net23),
    .X(net990));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer11 (.A(net990),
    .X(net991));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer12 (.A(net991),
    .X(net992));
 sky130_fd_sc_hd__a41o_1 clone13 (.A1(net1018),
    .A2(net15),
    .A3(net1020),
    .A4(net1042),
    .B1(net12),
    .X(net993));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer14 (.A(net114),
    .X(net994));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer15 (.A(net994),
    .X(net995));
 sky130_fd_sc_hd__a41o_1 clone16 (.A1(net948),
    .A2(net960),
    .A3(net969),
    .A4(net949),
    .B1(net976),
    .X(net996));
 sky130_fd_sc_hd__clkbuf_1 clone17 (.A(net822),
    .X(net997));
 sky130_fd_sc_hd__clkbuf_4 clone18 (.A(net22),
    .X(net998));
 sky130_fd_sc_hd__clkbuf_1 clone19 (.A(net732),
    .X(net999));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer20 (.A(net1010),
    .X(net1000));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer21 (.A(net1008),
    .X(net1001));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer22 (.A(net927),
    .X(net1002));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer23 (.A(net1002),
    .X(net1003));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer24 (.A(net927),
    .X(net1004));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer25 (.A(net1004),
    .X(net1005));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer26 (.A(net260),
    .X(net1006));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer27 (.A(net1006),
    .X(net1007));
 sky130_fd_sc_hd__clkbuf_1 clone28 (.A(net6),
    .X(net1008));
 sky130_fd_sc_hd__clkbuf_1 clone29 (.A(net14),
    .X(net1009));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer30 (.A(net14),
    .X(net1010));
 sky130_fd_sc_hd__clkbuf_1 clone31 (.A(net1012),
    .X(net1011));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer32 (.A(net31),
    .X(net1012));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer33 (.A(net1015),
    .X(net1013));
 sky130_fd_sc_hd__clkbuf_1 clone34 (.A(net20),
    .X(net1014));
 sky130_fd_sc_hd__clkbuf_1 clone35 (.A(net21),
    .X(net1015));
 sky130_fd_sc_hd__clkbuf_1 clone36 (.A(net872),
    .X(net1016));
 sky130_fd_sc_hd__clkbuf_1 clone37 (.A(net8),
    .X(net1017));
 sky130_fd_sc_hd__clkbuf_1 clone38 (.A(net921),
    .X(net1018));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer39 (.A(net978),
    .X(net1019));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(net640),
    .X(net1024));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(net658),
    .X(net1025));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(net668),
    .X(net1026));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(net660),
    .X(net1027));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(net670),
    .X(net1028));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(net663),
    .X(net1029));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(net543),
    .X(net1030));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(net589),
    .X(net1031));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(net679),
    .X(net1032));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(net647),
    .X(net1033));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(net545),
    .X(net1034));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(net686),
    .X(net1035));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(net537),
    .X(net1036));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(net662),
    .X(net1037));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(net941),
    .X(net1038));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(net664),
    .X(net1039));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(net537),
    .X(net1040));
 sky130_fd_sc_hd__buf_6 fanout1 (.A(net925),
    .X(net1020));
 sky130_fd_sc_hd__clkbuf_2 fanout2 (.A(net976),
    .X(net1021));
 sky130_fd_sc_hd__buf_4 fanout3 (.A(net949),
    .X(net1022));
 sky130_fd_sc_hd__clkbuf_4 fanout4 (.A(net969),
    .X(net1023));
 sky130_fd_sc_hd__clkbuf_4 fanout5 (.A(net960),
    .X(net1041));
 sky130_fd_sc_hd__clkbuf_1 fanout6 (.A(net756),
    .X(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_A (.DIODE(clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(in0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(in1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(in10));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(in11));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(in12));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(in13));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(in14));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(in15));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(in16));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(in17));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(in18));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(in19));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(in2));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(in20));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(in21));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(in22));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(in23));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(in24));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(in25));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(in26));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(in27));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_A (.DIODE(in28));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_A (.DIODE(in29));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_A (.DIODE(in3));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_A (.DIODE(in30));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_A (.DIODE(in31));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_A (.DIODE(in32));
 sky130_fd_sc_hd__diode_2 ANTENNA_input28_A (.DIODE(in33));
 sky130_fd_sc_hd__diode_2 ANTENNA_input29_A (.DIODE(in34));
 sky130_fd_sc_hd__diode_2 ANTENNA_input30_A (.DIODE(in35));
 sky130_fd_sc_hd__diode_2 ANTENNA_input31_A (.DIODE(in36));
 sky130_fd_sc_hd__diode_2 ANTENNA_input32_A (.DIODE(in37));
 sky130_fd_sc_hd__diode_2 ANTENNA_input33_A (.DIODE(in38));
 sky130_fd_sc_hd__diode_2 ANTENNA_input34_A (.DIODE(in39));
 sky130_fd_sc_hd__diode_2 ANTENNA_input35_A (.DIODE(in4));
 sky130_fd_sc_hd__diode_2 ANTENNA_input36_A (.DIODE(in40));
 sky130_fd_sc_hd__diode_2 ANTENNA_input37_A (.DIODE(in41));
 sky130_fd_sc_hd__diode_2 ANTENNA_input38_A (.DIODE(in42));
 sky130_fd_sc_hd__diode_2 ANTENNA_input39_A (.DIODE(in43));
 sky130_fd_sc_hd__diode_2 ANTENNA_input40_A (.DIODE(in44));
 sky130_fd_sc_hd__diode_2 ANTENNA_input41_A (.DIODE(in45));
 sky130_fd_sc_hd__diode_2 ANTENNA_input42_A (.DIODE(in46));
 sky130_fd_sc_hd__diode_2 ANTENNA_input43_A (.DIODE(in47));
 sky130_fd_sc_hd__diode_2 ANTENNA_input44_A (.DIODE(in48));
 sky130_fd_sc_hd__diode_2 ANTENNA_input45_A (.DIODE(in49));
 sky130_fd_sc_hd__diode_2 ANTENNA_input46_A (.DIODE(in5));
 sky130_fd_sc_hd__diode_2 ANTENNA_input47_A (.DIODE(in50));
 sky130_fd_sc_hd__diode_2 ANTENNA_input48_A (.DIODE(in51));
 sky130_fd_sc_hd__diode_2 ANTENNA_input49_A (.DIODE(in52));
 sky130_fd_sc_hd__diode_2 ANTENNA_input50_A (.DIODE(in53));
 sky130_fd_sc_hd__diode_2 ANTENNA_input51_A (.DIODE(in54));
 sky130_fd_sc_hd__diode_2 ANTENNA_input52_A (.DIODE(in55));
 sky130_fd_sc_hd__diode_2 ANTENNA_input53_A (.DIODE(in56));
 sky130_fd_sc_hd__diode_2 ANTENNA_input54_A (.DIODE(in57));
 sky130_fd_sc_hd__diode_2 ANTENNA_input55_A (.DIODE(in58));
 sky130_fd_sc_hd__diode_2 ANTENNA_input56_A (.DIODE(in59));
 sky130_fd_sc_hd__diode_2 ANTENNA_input57_A (.DIODE(in6));
 sky130_fd_sc_hd__diode_2 ANTENNA_input58_A (.DIODE(in60));
 sky130_fd_sc_hd__diode_2 ANTENNA_input59_A (.DIODE(in61));
 sky130_fd_sc_hd__diode_2 ANTENNA_input60_A (.DIODE(in62));
 sky130_fd_sc_hd__diode_2 ANTENNA_input61_A (.DIODE(in63));
 sky130_fd_sc_hd__diode_2 ANTENNA_input62_A (.DIODE(in64));
 sky130_fd_sc_hd__diode_2 ANTENNA_input63_A (.DIODE(in65));
 sky130_fd_sc_hd__diode_2 ANTENNA_input64_A (.DIODE(in66));
 sky130_fd_sc_hd__diode_2 ANTENNA_input65_A (.DIODE(in67));
 sky130_fd_sc_hd__diode_2 ANTENNA_input66_A (.DIODE(in68));
 sky130_fd_sc_hd__diode_2 ANTENNA_input67_A (.DIODE(in69));
 sky130_fd_sc_hd__diode_2 ANTENNA_input68_A (.DIODE(in7));
 sky130_fd_sc_hd__diode_2 ANTENNA_input69_A (.DIODE(in70));
 sky130_fd_sc_hd__diode_2 ANTENNA_input70_A (.DIODE(in71));
 sky130_fd_sc_hd__diode_2 ANTENNA_input71_A (.DIODE(in72));
 sky130_fd_sc_hd__diode_2 ANTENNA_input72_A (.DIODE(in73));
 sky130_fd_sc_hd__diode_2 ANTENNA_input73_A (.DIODE(in74));
 sky130_fd_sc_hd__diode_2 ANTENNA_input74_A (.DIODE(in75));
 sky130_fd_sc_hd__diode_2 ANTENNA_input75_A (.DIODE(in76));
 sky130_fd_sc_hd__diode_2 ANTENNA_input76_A (.DIODE(in77));
 sky130_fd_sc_hd__diode_2 ANTENNA_input77_A (.DIODE(in78));
 sky130_fd_sc_hd__diode_2 ANTENNA_input78_A (.DIODE(in79));
 sky130_fd_sc_hd__diode_2 ANTENNA_input79_A (.DIODE(in8));
 sky130_fd_sc_hd__diode_2 ANTENNA_input80_A (.DIODE(in80));
 sky130_fd_sc_hd__diode_2 ANTENNA_input81_A (.DIODE(in81));
 sky130_fd_sc_hd__diode_2 ANTENNA_input82_A (.DIODE(in82));
 sky130_fd_sc_hd__diode_2 ANTENNA_input83_A (.DIODE(in83));
 sky130_fd_sc_hd__diode_2 ANTENNA_input84_A (.DIODE(in84));
 sky130_fd_sc_hd__diode_2 ANTENNA_input85_A (.DIODE(in85));
 sky130_fd_sc_hd__diode_2 ANTENNA_input86_A (.DIODE(in86));
 sky130_fd_sc_hd__diode_2 ANTENNA_input87_A (.DIODE(in87));
 sky130_fd_sc_hd__diode_2 ANTENNA_input88_A (.DIODE(in88));
 sky130_fd_sc_hd__diode_2 ANTENNA_input89_A (.DIODE(in89));
 sky130_fd_sc_hd__diode_2 ANTENNA_input90_A (.DIODE(in9));
 sky130_fd_sc_hd__diode_2 ANTENNA_input91_A (.DIODE(in90));
 sky130_fd_sc_hd__diode_2 ANTENNA_input92_A (.DIODE(in91));
 sky130_fd_sc_hd__diode_2 ANTENNA_input93_A (.DIODE(in92));
 sky130_fd_sc_hd__diode_2 ANTENNA_input94_A (.DIODE(in93));
 sky130_fd_sc_hd__diode_2 ANTENNA_input95_A (.DIODE(in94));
 sky130_fd_sc_hd__diode_2 ANTENNA_input96_A (.DIODE(in95));
 sky130_fd_sc_hd__diode_2 ANTENNA_input97_A (.DIODE(in96));
 sky130_fd_sc_hd__diode_2 ANTENNA_input98_A (.DIODE(in97));
 sky130_fd_sc_hd__diode_2 ANTENNA_input99_A (.DIODE(in98));
 sky130_fd_sc_hd__diode_2 ANTENNA_input100_A (.DIODE(in99));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_A2 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_A0 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_A3 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_S0 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_c369_A3 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_A2 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_S0 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_c106_S1 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_c105_A2 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_c104_S0 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_c102_X (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout210_A (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_A0 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_X (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA_c530_A1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_A0 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA_c311_S0 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_A2 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_A0 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA_c270_A1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA_c264_X (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_A0 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c560_A1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c542_A2 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c412_A0 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_S0 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c267_X (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout193_A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_S0 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_A2 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_X (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_A2 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_A0 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_A1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_A2 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_A2 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_A0 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c269_X (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c546_A3 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA_c541_S0 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA_c536_A0 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA_c533_D (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_A3 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA_c272_A1 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA_c271_X (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_A1 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_c544_A3 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_A0 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_A2 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_c295_A1 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_c273_A1 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_c272_X (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_A2 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_c313_A0 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_A0 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_A2 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_c279_A3 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_c278_S0 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_c277_A1 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_c276_A3 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_c274_X (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout179_A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout178_A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c276_X (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c562_A3 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c555_A0 (.DIODE(net1043));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_A2 (.DIODE(net1043));
 sky130_fd_sc_hd__diode_2 ANTENNA_c536_A1 (.DIODE(net1043));
 sky130_fd_sc_hd__diode_2 ANTENNA_c410_A3 (.DIODE(net1043));
 sky130_fd_sc_hd__diode_2 ANTENNA_c402_A2 (.DIODE(net1043));
 sky130_fd_sc_hd__diode_2 ANTENNA_c397_A3 (.DIODE(net1043));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_A4 (.DIODE(net1043));
 sky130_fd_sc_hd__diode_2 ANTENNA_c283_S0 (.DIODE(net1043));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_A1 (.DIODE(net1043));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_X (.DIODE(net1043));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_A0 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c534_A2 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c529_A2 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_S0 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_A0 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c283_A2 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_X (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_A0 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_A1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_A2 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c557_A1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c428_A2 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_A0 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c283_X (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_A0 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_A2 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A1 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_A2 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_c668_A1 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_c554_A1 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_c400_SCD (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_A1 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_X (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone13_B1 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_A0 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_A3 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_A4 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_A2 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_c148_A1 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_B1 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_A2 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_c143_B1 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_X (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_A2 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_S0 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_A1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_A3 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c344_A2 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_A1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_A0 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c286_X (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_A0 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_A3 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_A4 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_A2 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_A1 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_X (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_A1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_A3 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_A0 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c558_A0 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c365_A2 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_A1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_A3 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_A1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_A4 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_A3 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_X (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_A2 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_A3 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_A1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_A3 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_A1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_A2 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_A0 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_X (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_A0 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_A2 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_A2 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c587_A2 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_A2 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c297_A2 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c295_A0 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_X (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_A0 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_A1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_S0 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c297_A1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c295_A2 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_X (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout176_A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_A2 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_X (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_A1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_A2 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_A2 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_S0 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_A1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_A0 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_A2 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_A1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_X (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_A0 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_A3 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_A2 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_c371_A1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_A1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_A2 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_A3 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_B1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_c295_X (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_A0 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_A3 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_A1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_A3 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_A2 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_S1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_X (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout206_A (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_S0 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_X (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_A0 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_c321_A3 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_S1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_A2 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_A2 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_X (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_A0 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA_c559_A1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_A2 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_A1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_A0 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_A4 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_X (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_A1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_A0 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_A1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_c323_A1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_A0 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_X (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_c757_A2 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_S0 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_A0 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_A1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_A0 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_X (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone13_A2 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_c283_A0 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_c270_A0 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_A1 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_c148_A4 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_A2 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_c143_X (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_A3 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_A1 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_A0 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_A3 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_A0 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_S0 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_X (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout202_A (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c677_A0 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_X (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_A1 (.DIODE(net1051));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_A0 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_A2 (.DIODE(net1051));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_S1 (.DIODE(net1051));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_S0 (.DIODE(net1051));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_X (.DIODE(net1051));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge797_B (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA_c372_X (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_A3 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_A0 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_c610_A1 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_S0 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_c402_A4 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_c400_D (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_c397_B1 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_X (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_A1 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_A0 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_A0 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_A2 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA_c542_A3 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA_c428_S0 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA_c406_A3 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA_c397_X (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_A1 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_c564_A3 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_c416_A2 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_c409_A0 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_c406_A0 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_c398_X (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout186_A (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_c533_RESET_B (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_A1 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_c400_SET_B (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_c399_X (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone34_A (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout194_A (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA_c586_A2 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_X (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout226_A (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_A3 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_c400_Q (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_c685_A0 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_A1 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_A1 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_c403_B1 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_c402_A1 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_c401_X (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_A0 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_c669_A2 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_A3 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_A0 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_A2 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_A3 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_c415_S1 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_c410_A0 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_c409_X (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone35_A (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout188_A (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout187_A (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_X (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_A0 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_A1 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_S0 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_A0 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA_c416_A0 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA_c414_A2 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA_c412_X (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_A2 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_S0 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA_c686_A0 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA_c555_A1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA_c427_A0 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_A1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_A2 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_X (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA_c577_A0 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA_c565_A1 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_A1 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_A2 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_X (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone18_A (.DIODE(net1050));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer1_A (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout184_A (.DIODE(net1050));
 sky130_fd_sc_hd__diode_2 ANTENNA_c671_A2 (.DIODE(net1050));
 sky130_fd_sc_hd__diode_2 ANTENNA_c661_A2 (.DIODE(net1050));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_X (.DIODE(net1050));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_A0 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_A1 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_S0 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA_c430_A1 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_A1 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_A2 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_S0 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_X (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_A0 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_A3 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_S0 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA_c430_A4 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_X (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA_c763_A2 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_c695_A3 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_A2 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_A1 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_A3 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_A0 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_A1 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_c427_X (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_c571_A0 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_A2 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA_c560_A0 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_A2 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA_c437_A1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA_c434_A3 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_X (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_A0 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_A0 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_A3 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_A1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA_c434_A1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_A0 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA_c431_D (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA_c430_X (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_A2 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_A3 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_A2 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_c434_A2 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_c431_Q_N (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_c687_A0 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_A1 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_A2 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_A3 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_X (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA_c482_A0 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_A2 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_X (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA_c739_A2 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A0 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_A3 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_A2 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_A1 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_X (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_A1 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_A1 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA_c577_A1 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_A3 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_A2 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA_c458_A1 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_A1 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_A3 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_A0 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_A2 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_X (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout215_A (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_A3 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_X (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_A0 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_A3 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_A1 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_X (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA_c323_A0 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c313_A1 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_S0 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_A2 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_A1 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_A3 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_A4 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_A1 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_A0 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_A4 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_X (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c743_A2 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_A1 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_c610_A3 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_A1 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_X (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_A0 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_A1 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_A0 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c437_A2 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_A4 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c286_A4 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_A1 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_A1 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_X (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net290_A (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_X (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_A0 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_S0 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_A2 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_A1 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c237_A3 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c235_A2 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c104_X (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout177_A (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_A0 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_c757_A1 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_X (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_A0 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_A1 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA_c546_A2 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA_c545_A3 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA_c532_X (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_A0 (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA_c571_A1 (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA_c558_A3 (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA_c533_Q (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net315_A (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_c538_X (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_A0 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_A2 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_A2 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_A1 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA_c677_A3 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA_c660_A2 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA_c571_A2 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA_c563_A1 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA_c549_X (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_A0 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_S0 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_A2 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_A2 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_c557_A2 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_c556_A3 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_c554_A0 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_X (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_c562_A0 (.DIODE(net1075));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_A3 (.DIODE(net1075));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_A0 (.DIODE(net1075));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_S0 (.DIODE(net1075));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_A0 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_A3 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_X (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout175_A (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_A0 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_X (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net345_A (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_X (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_A0 (.DIODE(net1068));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_A2 (.DIODE(net1069));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_A1 (.DIODE(net1067));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_A0 (.DIODE(net1066));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_A0 (.DIODE(net1066));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_A2 (.DIODE(net1066));
 sky130_fd_sc_hd__diode_2 ANTENNA_c198_S0 (.DIODE(net1070));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_A3 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_X (.DIODE(net1066));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_A0 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_A2 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_A0 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_A2 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_A1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_A0 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_X (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge805_D (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_X (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_S0 (.DIODE(net1072));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_A3 (.DIODE(net1072));
 sky130_fd_sc_hd__diode_2 ANTENNA_c691_A0 (.DIODE(net1071));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_A3 (.DIODE(net1072));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_A3 (.DIODE(net1071));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_S1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_A0 (.DIODE(net1074));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_A0 (.DIODE(net1071));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_S0 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_X (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_A0 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_A3 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_A2 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_A2 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_A1 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_A1 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_X (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_c764_A2 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_A2 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_A3 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_X (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A2 (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_A1 (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_A3 (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_X (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_A0 (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA_c745_A1 (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_A1 (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA_c681_A1 (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA_c677_A2 (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA_c669_X (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA_c241_A1 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_c240_A2 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_c237_A0 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_c222_S0 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_A4 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_c184_A2 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_X (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge835_B (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA_c686_X (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_A2 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_A0 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_A1 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_A1 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_A0 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_c311_A2 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_A2 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_c184_A0 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_S0 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_X (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_A0 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_S0 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_S1 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_S0 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_c180_A0 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_X (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout183_A (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_A1 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA_c446_A0 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA_c180_X (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_A0 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_A0 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_A3 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_B1 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_c182_X (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge773_Q (.DIODE(net529));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_S1 (.DIODE(net529));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_S0 (.DIODE(net529));
 sky130_fd_sc_hd__diode_2 ANTENNA_c566_A3 (.DIODE(net529));
 sky130_fd_sc_hd__diode_2 ANTENNA_c549_A2 (.DIODE(net529));
 sky130_fd_sc_hd__diode_2 ANTENNA_c545_S0 (.DIODE(net529));
 sky130_fd_sc_hd__diode_2 ANTENNA_c539_S0 (.DIODE(net529));
 sky130_fd_sc_hd__diode_2 ANTENNA_c538_A2 (.DIODE(net529));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_A3 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_S0 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_A0 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_A2 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA_c577_A3 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_S0 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_A1 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_A2 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_A2 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_X (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout224_A (.DIODE(net533));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_S0 (.DIODE(net533));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge777_Q (.DIODE(net533));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge779_Q (.DIODE(net536));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_S0 (.DIODE(net536));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_A3 (.DIODE(net536));
 sky130_fd_sc_hd__diode_2 ANTENNA_c437_A3 (.DIODE(net536));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge780_Q (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_S0 (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_A3 (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_S0 (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA_c191_S1 (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_A3 (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge784_Q (.DIODE(net542));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_S0 (.DIODE(net542));
 sky130_fd_sc_hd__diode_2 ANTENNA_c723_A3 (.DIODE(net542));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_A3 (.DIODE(net542));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_A3 (.DIODE(net542));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold50_A (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge785_Q (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_S0 (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA_c372_S1 (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_A3 (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_A1 (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA_c234_S0 (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA_c203_S1 (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge792_Q (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA_c371_S0 (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA_c368_S0 (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_A3 (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_A3 (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_A4 (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_S0 (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_A3 (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_S0 (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_S1 (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_B1 (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_B1 (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA_c286_B1 (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA_c221_A3 (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_B1 (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_A0 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_A1 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_S0 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_A2 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_A1 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_c194_A3 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_c191_S0 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_c190_X (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge809_Q (.DIODE(net567));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_A2 (.DIODE(net567));
 sky130_fd_sc_hd__diode_2 ANTENNA_c696_A3 (.DIODE(net567));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_S1 (.DIODE(net567));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_A2 (.DIODE(net567));
 sky130_fd_sc_hd__diode_2 ANTENNA_c666_A3 (.DIODE(net567));
 sky130_fd_sc_hd__diode_2 ANTENNA_c661_S1 (.DIODE(net567));
 sky130_fd_sc_hd__diode_2 ANTENNA_c565_A3 (.DIODE(net567));
 sky130_fd_sc_hd__diode_2 ANTENNA_c563_A2 (.DIODE(net567));
 sky130_fd_sc_hd__diode_2 ANTENNA_c542_S1 (.DIODE(net567));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_A0 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_A3 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_A1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_c587_A1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_A2 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_A3 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_A3 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_c191_X (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge822_Q_N (.DIODE(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_A1 (.DIODE(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA_c373_S0 (.DIODE(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge828_Q (.DIODE(net584));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_A2 (.DIODE(net584));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_A2 (.DIODE(net584));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_S0 (.DIODE(net584));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_S0 (.DIODE(net584));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge830_Q (.DIODE(net586));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_S0 (.DIODE(net586));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_S0 (.DIODE(net586));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_A3 (.DIODE(net586));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_A1 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_A0 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_A2 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_A2 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_A2 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_B1 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA_c194_A1 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_X (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge833_Q (.DIODE(net590));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_S0 (.DIODE(net590));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_S0 (.DIODE(net590));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_A2 (.DIODE(net590));
 sky130_fd_sc_hd__diode_2 ANTENNA_c371_S1 (.DIODE(net590));
 sky130_fd_sc_hd__diode_2 ANTENNA_c366_S1 (.DIODE(net590));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_S0 (.DIODE(net590));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_S0 (.DIODE(net590));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_S0 (.DIODE(net590));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone28_A (.DIODE(net1048));
 sky130_fd_sc_hd__diode_2 ANTENNA_c134_A3 (.DIODE(net1048));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout227_A (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_S0 (.DIODE(net1048));
 sky130_fd_sc_hd__diode_2 ANTENNA_c191_A3 (.DIODE(net1048));
 sky130_fd_sc_hd__diode_2 ANTENNA_c143_A4 (.DIODE(net1048));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_X (.DIODE(net1048));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_A1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_A1 (.DIODE(net1049));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_A1 (.DIODE(net1049));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_A1 (.DIODE(net1049));
 sky130_fd_sc_hd__diode_2 ANTENNA_c228_A1 (.DIODE(net1049));
 sky130_fd_sc_hd__diode_2 ANTENNA_c220_A1 (.DIODE(net1049));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_S0 (.DIODE(net1049));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_A2 (.DIODE(net1049));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_A0 (.DIODE(net1049));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_A1 (.DIODE(net1049));
 sky130_fd_sc_hd__diode_2 ANTENNA_c194_X (.DIODE(net1049));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge841_Q (.DIODE(net601));
 sky130_fd_sc_hd__diode_2 ANTENNA_c764_S0 (.DIODE(net601));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_A3 (.DIODE(net601));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_S1 (.DIODE(net601));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_S0 (.DIODE(net601));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge842_Q (.DIODE(net602));
 sky130_fd_sc_hd__diode_2 ANTENNA_c742_S0 (.DIODE(net602));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_A1 (.DIODE(net602));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_S0 (.DIODE(net602));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_A2 (.DIODE(net602));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge847_Q_N (.DIODE(net605));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_A3 (.DIODE(net605));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_S1 (.DIODE(net605));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_S1 (.DIODE(net605));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_S0 (.DIODE(net605));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge852_Q (.DIODE(net612));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_A3 (.DIODE(net612));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_A3 (.DIODE(net612));
 sky130_fd_sc_hd__diode_2 ANTENNA_c723_S1 (.DIODE(net612));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge853_Q_N (.DIODE(net613));
 sky130_fd_sc_hd__diode_2 ANTENNA_c745_S0 (.DIODE(net613));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_S0 (.DIODE(net613));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_A3 (.DIODE(net613));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge854_Q (.DIODE(net615));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_S0 (.DIODE(net615));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_S1 (.DIODE(net615));
 sky130_fd_sc_hd__diode_2 ANTENNA_c615_S0 (.DIODE(net615));
 sky130_fd_sc_hd__diode_2 ANTENNA_c502_S1 (.DIODE(net615));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_S0 (.DIODE(net615));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_S1 (.DIODE(net615));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge855_Q (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_S0 (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_A3 (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA_c747_A3 (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA_c742_S1 (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA_c698_A2 (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_A1 (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge856_Q (.DIODE(net617));
 sky130_fd_sc_hd__diode_2 ANTENNA_c745_S1 (.DIODE(net617));
 sky130_fd_sc_hd__diode_2 ANTENNA_c744_A3 (.DIODE(net617));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_A2 (.DIODE(net617));
 sky130_fd_sc_hd__diode_2 ANTENNA_c482_S1 (.DIODE(net617));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_S1 (.DIODE(net617));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_S0 (.DIODE(net617));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_A3 (.DIODE(net617));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge857_Q (.DIODE(net618));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_S0 (.DIODE(net618));
 sky130_fd_sc_hd__diode_2 ANTENNA_c724_A2 (.DIODE(net618));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_A2 (.DIODE(net618));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_A3 (.DIODE(net618));
 sky130_fd_sc_hd__diode_2 ANTENNA_c703_A1 (.DIODE(net618));
 sky130_fd_sc_hd__diode_2 ANTENNA_c702_A4 (.DIODE(net618));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge858_Q_N (.DIODE(net619));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_S0 (.DIODE(net619));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_A3 (.DIODE(net619));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_S1 (.DIODE(net619));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge859_Q (.DIODE(net622));
 sky130_fd_sc_hd__diode_2 ANTENNA_c701_S0 (.DIODE(net622));
 sky130_fd_sc_hd__diode_2 ANTENNA_c685_A3 (.DIODE(net622));
 sky130_fd_sc_hd__diode_2 ANTENNA_c672_S0 (.DIODE(net622));
 sky130_fd_sc_hd__diode_2 ANTENNA_s860_Q_N (.DIODE(net623));
 sky130_fd_sc_hd__diode_2 ANTENNA_c695_S0 (.DIODE(net623));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_A3 (.DIODE(net623));
 sky130_fd_sc_hd__diode_2 ANTENNA_c685_S0 (.DIODE(net623));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_S0 (.DIODE(net623));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_S1 (.DIODE(net623));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_S0 (.DIODE(net623));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_S1 (.DIODE(net623));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_S1 (.DIODE(net623));
 sky130_fd_sc_hd__diode_2 ANTENNA_s860_Q (.DIODE(net624));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_S1 (.DIODE(net624));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_S1 (.DIODE(net624));
 sky130_fd_sc_hd__diode_2 ANTENNA_c724_A3 (.DIODE(net624));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_A3 (.DIODE(net624));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_S1 (.DIODE(net624));
 sky130_fd_sc_hd__diode_2 ANTENNA_c236_A2 (.DIODE(net624));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_S1 (.DIODE(net624));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_S1 (.DIODE(net624));
 sky130_fd_sc_hd__diode_2 ANTENNA_s861_Q_N (.DIODE(net625));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_A3 (.DIODE(net625));
 sky130_fd_sc_hd__diode_2 ANTENNA_c226_S0 (.DIODE(net625));
 sky130_fd_sc_hd__diode_2 ANTENNA_c220_S1 (.DIODE(net625));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_S1 (.DIODE(net625));
 sky130_fd_sc_hd__diode_2 ANTENNA_c190_S1 (.DIODE(net625));
 sky130_fd_sc_hd__diode_2 ANTENNA_s861_Q (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA_c762_S0 (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_S0 (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA_c747_S0 (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_A3 (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_S0 (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_S1 (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA_s862_Q (.DIODE(net627));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_S1 (.DIODE(net627));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_S0 (.DIODE(net627));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_S1 (.DIODE(net627));
 sky130_fd_sc_hd__diode_2 ANTENNA_c231_S1 (.DIODE(net627));
 sky130_fd_sc_hd__diode_2 ANTENNA_c226_S1 (.DIODE(net627));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_S1 (.DIODE(net627));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_B1 (.DIODE(net627));
 sky130_fd_sc_hd__diode_2 ANTENNA_s863_Q (.DIODE(net628));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_A3 (.DIODE(net628));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_A3 (.DIODE(net628));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_S1 (.DIODE(net628));
 sky130_fd_sc_hd__diode_2 ANTENNA_c370_S0 (.DIODE(net628));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_S0 (.DIODE(net628));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_A3 (.DIODE(net628));
 sky130_fd_sc_hd__diode_2 ANTENNA_c311_S1 (.DIODE(net628));
 sky130_fd_sc_hd__diode_2 ANTENNA_c240_S1 (.DIODE(net628));
 sky130_fd_sc_hd__diode_2 ANTENNA_c206_S1 (.DIODE(net628));
 sky130_fd_sc_hd__diode_2 ANTENNA_s864_Q (.DIODE(net629));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_A3 (.DIODE(net629));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_S1 (.DIODE(net629));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_S1 (.DIODE(net629));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_S0 (.DIODE(net629));
 sky130_fd_sc_hd__diode_2 ANTENNA_c241_S0 (.DIODE(net629));
 sky130_fd_sc_hd__diode_2 ANTENNA_c216_S1 (.DIODE(net629));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_S0 (.DIODE(net629));
 sky130_fd_sc_hd__diode_2 ANTENNA_s870_Q_N (.DIODE(net637));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_S1 (.DIODE(net637));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_S0 (.DIODE(net637));
 sky130_fd_sc_hd__diode_2 ANTENNA_c672_S1 (.DIODE(net637));
 sky130_fd_sc_hd__diode_2 ANTENNA_c528_B1 (.DIODE(net637));
 sky130_fd_sc_hd__diode_2 ANTENNA_c404_S1 (.DIODE(net637));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_B1 (.DIODE(net637));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap220_A (.DIODE(net638));
 sky130_fd_sc_hd__diode_2 ANTENNA_s870_Q (.DIODE(net638));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_S0 (.DIODE(net638));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout219_A (.DIODE(net639));
 sky130_fd_sc_hd__diode_2 ANTENNA_c698_A3 (.DIODE(net639));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_A2 (.DIODE(net639));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_S1 (.DIODE(net639));
 sky130_fd_sc_hd__diode_2 ANTENNA_c764_S1 (.DIODE(net639));
 sky130_fd_sc_hd__diode_2 ANTENNA_s871_Q (.DIODE(net639));
 sky130_fd_sc_hd__diode_2 ANTENNA_s873_Q (.DIODE(net641));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_S1 (.DIODE(net641));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_S1 (.DIODE(net641));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_S0 (.DIODE(net641));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_S1 (.DIODE(net641));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_S1 (.DIODE(net641));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_S1 (.DIODE(net641));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap218_A (.DIODE(net642));
 sky130_fd_sc_hd__diode_2 ANTENNA_s874_Q (.DIODE(net642));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_S0 (.DIODE(net642));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_S0 (.DIODE(net642));
 sky130_fd_sc_hd__diode_2 ANTENNA_s875_Q (.DIODE(net643));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_S1 (.DIODE(net643));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_S1 (.DIODE(net643));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_S0 (.DIODE(net643));
 sky130_fd_sc_hd__diode_2 ANTENNA_c321_S1 (.DIODE(net643));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_S1 (.DIODE(net643));
 sky130_fd_sc_hd__diode_2 ANTENNA_s876_Q_N (.DIODE(net644));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_A3 (.DIODE(net644));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_A3 (.DIODE(net644));
 sky130_fd_sc_hd__diode_2 ANTENNA_c323_S0 (.DIODE(net644));
 sky130_fd_sc_hd__diode_2 ANTENNA_s876_Q (.DIODE(net645));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_S0 (.DIODE(net645));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_S0 (.DIODE(net645));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_S1 (.DIODE(net645));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold53_A (.DIODE(net647));
 sky130_fd_sc_hd__diode_2 ANTENNA_s877_Q (.DIODE(net647));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_S0 (.DIODE(net647));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_S1 (.DIODE(net647));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_S0 (.DIODE(net647));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_S1 (.DIODE(net647));
 sky130_fd_sc_hd__diode_2 ANTENNA_s878_Q (.DIODE(net648));
 sky130_fd_sc_hd__diode_2 ANTENNA_c496_S1 (.DIODE(net648));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_S1 (.DIODE(net648));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_S1 (.DIODE(net648));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_S0 (.DIODE(net648));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_S1 (.DIODE(net648));
 sky130_fd_sc_hd__diode_2 ANTENNA_s879_Q (.DIODE(net649));
 sky130_fd_sc_hd__diode_2 ANTENNA_c610_S1 (.DIODE(net649));
 sky130_fd_sc_hd__diode_2 ANTENNA_c587_S1 (.DIODE(net649));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_S0 (.DIODE(net649));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_S1 (.DIODE(net649));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_A2 (.DIODE(net649));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_S1 (.DIODE(net649));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net653_A (.DIODE(net653));
 sky130_fd_sc_hd__diode_2 ANTENNA_s883_GCLK (.DIODE(net653));
 sky130_fd_sc_hd__diode_2 ANTENNA_s884_Q_N (.DIODE(net654));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_A3 (.DIODE(net654));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_S0 (.DIODE(net654));
 sky130_fd_sc_hd__diode_2 ANTENNA_c531_S1 (.DIODE(net654));
 sky130_fd_sc_hd__diode_2 ANTENNA_c413_S0 (.DIODE(net654));
 sky130_fd_sc_hd__diode_2 ANTENNA_c412_A3 (.DIODE(net654));
 sky130_fd_sc_hd__diode_2 ANTENNA_c411_S1 (.DIODE(net654));
 sky130_fd_sc_hd__diode_2 ANTENNA_c409_S0 (.DIODE(net654));
 sky130_fd_sc_hd__diode_2 ANTENNA_s884_Q (.DIODE(net655));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_A3 (.DIODE(net655));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_S1 (.DIODE(net655));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_S1 (.DIODE(net655));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_A3 (.DIODE(net655));
 sky130_fd_sc_hd__diode_2 ANTENNA_c586_S0 (.DIODE(net655));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_S1 (.DIODE(net655));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_A2 (.DIODE(net655));
 sky130_fd_sc_hd__diode_2 ANTENNA_c414_S0 (.DIODE(net655));
 sky130_fd_sc_hd__diode_2 ANTENNA_s885_Q_N (.DIODE(net656));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_S0 (.DIODE(net656));
 sky130_fd_sc_hd__diode_2 ANTENNA_c529_B1 (.DIODE(net656));
 sky130_fd_sc_hd__diode_2 ANTENNA_c412_S0 (.DIODE(net656));
 sky130_fd_sc_hd__diode_2 ANTENNA_c409_S1 (.DIODE(net656));
 sky130_fd_sc_hd__diode_2 ANTENNA_s885_Q (.DIODE(net657));
 sky130_fd_sc_hd__diode_2 ANTENNA_c665_S0 (.DIODE(net657));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_S1 (.DIODE(net657));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_S1 (.DIODE(net657));
 sky130_fd_sc_hd__diode_2 ANTENNA_c408_S1 (.DIODE(net657));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_A1 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_A0 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_A0 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_A0 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_X (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold47_A (.DIODE(net660));
 sky130_fd_sc_hd__diode_2 ANTENNA_s888_Q (.DIODE(net660));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_S0 (.DIODE(net660));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_S1 (.DIODE(net660));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_S1 (.DIODE(net660));
 sky130_fd_sc_hd__diode_2 ANTENNA_c430_B1 (.DIODE(net660));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_B1 (.DIODE(net660));
 sky130_fd_sc_hd__diode_2 ANTENNA_c427_S1 (.DIODE(net660));
 sky130_fd_sc_hd__diode_2 ANTENNA_s889_Q (.DIODE(net661));
 sky130_fd_sc_hd__diode_2 ANTENNA_c633_S1 (.DIODE(net661));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_S0 (.DIODE(net661));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_S1 (.DIODE(net661));
 sky130_fd_sc_hd__diode_2 ANTENNA_c615_S1 (.DIODE(net661));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_A3 (.DIODE(net661));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_S0 (.DIODE(net661));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_S1 (.DIODE(net661));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_S1 (.DIODE(net661));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_S1 (.DIODE(net661));
 sky130_fd_sc_hd__diode_2 ANTENNA_s892_Q (.DIODE(net665));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_A3 (.DIODE(net665));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_A3 (.DIODE(net665));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_S1 (.DIODE(net665));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_S1 (.DIODE(net665));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_S1 (.DIODE(net665));
 sky130_fd_sc_hd__diode_2 ANTENNA_s893_Q_N (.DIODE(net666));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_A3 (.DIODE(net666));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_S1 (.DIODE(net666));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_S0 (.DIODE(net666));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_S1 (.DIODE(net666));
 sky130_fd_sc_hd__diode_2 ANTENNA_s893_Q (.DIODE(net667));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_A3 (.DIODE(net667));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_S1 (.DIODE(net667));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_S1 (.DIODE(net667));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_S1 (.DIODE(net667));
 sky130_fd_sc_hd__diode_2 ANTENNA_c446_S1 (.DIODE(net667));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_A0 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_S1 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_A3 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_A1 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_X (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net673_A (.DIODE(net673));
 sky130_fd_sc_hd__diode_2 ANTENNA_s899_GCLK (.DIODE(net673));
 sky130_fd_sc_hd__diode_2 ANTENNA_s900_Q_N (.DIODE(net674));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_S0 (.DIODE(net674));
 sky130_fd_sc_hd__diode_2 ANTENNA_c541_S1 (.DIODE(net674));
 sky130_fd_sc_hd__diode_2 ANTENNA_c536_S0 (.DIODE(net674));
 sky130_fd_sc_hd__diode_2 ANTENNA_c532_S1 (.DIODE(net674));
 sky130_fd_sc_hd__diode_2 ANTENNA_s900_Q (.DIODE(net675));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_S1 (.DIODE(net675));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_S1 (.DIODE(net675));
 sky130_fd_sc_hd__diode_2 ANTENNA_c549_A3 (.DIODE(net675));
 sky130_fd_sc_hd__diode_2 ANTENNA_c538_S1 (.DIODE(net675));
 sky130_fd_sc_hd__diode_2 ANTENNA_s901_Q_N (.DIODE(net676));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_S1 (.DIODE(net676));
 sky130_fd_sc_hd__diode_2 ANTENNA_c548_A3 (.DIODE(net676));
 sky130_fd_sc_hd__diode_2 ANTENNA_c547_A3 (.DIODE(net676));
 sky130_fd_sc_hd__diode_2 ANTENNA_s901_Q (.DIODE(net677));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_S1 (.DIODE(net677));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_S1 (.DIODE(net677));
 sky130_fd_sc_hd__diode_2 ANTENNA_c544_S0 (.DIODE(net677));
 sky130_fd_sc_hd__diode_2 ANTENNA_c536_S1 (.DIODE(net677));
 sky130_fd_sc_hd__diode_2 ANTENNA_c494_A0 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_S0 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_A3 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_A3 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_A1 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c216_A0 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_A2 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c203_X (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_s904_Q (.DIODE(net681));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_S1 (.DIODE(net681));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_S0 (.DIODE(net681));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_S1 (.DIODE(net681));
 sky130_fd_sc_hd__diode_2 ANTENNA_c549_S0 (.DIODE(net681));
 sky130_fd_sc_hd__diode_2 ANTENNA_c547_S1 (.DIODE(net681));
 sky130_fd_sc_hd__diode_2 ANTENNA_c546_S0 (.DIODE(net681));
 sky130_fd_sc_hd__diode_2 ANTENNA_s906_Q (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_S0 (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_S1 (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA_c556_S1 (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA_c548_S1 (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA_s907_Q (.DIODE(net684));
 sky130_fd_sc_hd__diode_2 ANTENNA_c702_B1 (.DIODE(net684));
 sky130_fd_sc_hd__diode_2 ANTENNA_c695_S1 (.DIODE(net684));
 sky130_fd_sc_hd__diode_2 ANTENNA_c676_A3 (.DIODE(net684));
 sky130_fd_sc_hd__diode_2 ANTENNA_c665_S1 (.DIODE(net684));
 sky130_fd_sc_hd__diode_2 ANTENNA_c549_S1 (.DIODE(net684));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_A0 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_A1 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_S0 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_c208_A0 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_X (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_s911_Q (.DIODE(net690));
 sky130_fd_sc_hd__diode_2 ANTENNA_c582_S0 (.DIODE(net690));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_S1 (.DIODE(net690));
 sky130_fd_sc_hd__diode_2 ANTENNA_c565_S0 (.DIODE(net690));
 sky130_fd_sc_hd__diode_2 ANTENNA_c563_S0 (.DIODE(net690));
 sky130_fd_sc_hd__diode_2 ANTENNA_c561_S1 (.DIODE(net690));
 sky130_fd_sc_hd__diode_2 ANTENNA_c560_S0 (.DIODE(net690));
 sky130_fd_sc_hd__diode_2 ANTENNA_c559_S1 (.DIODE(net690));
 sky130_fd_sc_hd__diode_2 ANTENNA_s918_Q_N (.DIODE(net698));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_S0 (.DIODE(net698));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_S0 (.DIODE(net698));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_S1 (.DIODE(net698));
 sky130_fd_sc_hd__diode_2 ANTENNA_c582_S1 (.DIODE(net698));
 sky130_fd_sc_hd__diode_2 ANTENNA_s918_Q (.DIODE(net699));
 sky130_fd_sc_hd__diode_2 ANTENNA_c757_S1 (.DIODE(net699));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_S0 (.DIODE(net699));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_S1 (.DIODE(net699));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_S1 (.DIODE(net699));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_S1 (.DIODE(net699));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_A1 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_A1 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_A1 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA_c228_S0 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA_c218_A2 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_A1 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_A3 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA_c205_X (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA_s920_Q (.DIODE(net700));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_S1 (.DIODE(net700));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_S1 (.DIODE(net700));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_S1 (.DIODE(net700));
 sky130_fd_sc_hd__diode_2 ANTENNA_s922_Q (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_S0 (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_S0 (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_S1 (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA_c743_S1 (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA_c614_S0 (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_S1 (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA_s923_Q (.DIODE(net703));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_S1 (.DIODE(net703));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_S1 (.DIODE(net703));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_S1 (.DIODE(net703));
 sky130_fd_sc_hd__diode_2 ANTENNA_c611_S1 (.DIODE(net703));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_S1 (.DIODE(net703));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_S1 (.DIODE(net703));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_S1 (.DIODE(net703));
 sky130_fd_sc_hd__diode_2 ANTENNA_s925_Q (.DIODE(net707));
 sky130_fd_sc_hd__diode_2 ANTENNA_c703_A3 (.DIODE(net707));
 sky130_fd_sc_hd__diode_2 ANTENNA_c671_S1 (.DIODE(net707));
 sky130_fd_sc_hd__diode_2 ANTENNA_c667_S1 (.DIODE(net707));
 sky130_fd_sc_hd__diode_2 ANTENNA_s926_Q (.DIODE(net708));
 sky130_fd_sc_hd__diode_2 ANTENNA_c746_S1 (.DIODE(net708));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_S1 (.DIODE(net708));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_S1 (.DIODE(net708));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_S0 (.DIODE(net708));
 sky130_fd_sc_hd__diode_2 ANTENNA_c686_S1 (.DIODE(net708));
 sky130_fd_sc_hd__diode_2 ANTENNA_c680_S0 (.DIODE(net708));
 sky130_fd_sc_hd__diode_2 ANTENNA_c678_A2 (.DIODE(net708));
 sky130_fd_sc_hd__diode_2 ANTENNA_c676_S0 (.DIODE(net708));
 sky130_fd_sc_hd__diode_2 ANTENNA_c674_S1 (.DIODE(net708));
 sky130_fd_sc_hd__diode_2 ANTENNA_s927_Q (.DIODE(net709));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_S1 (.DIODE(net709));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_S0 (.DIODE(net709));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_S1 (.DIODE(net709));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_A2 (.DIODE(net709));
 sky130_fd_sc_hd__diode_2 ANTENNA_c693_S0 (.DIODE(net709));
 sky130_fd_sc_hd__diode_2 ANTENNA_c681_S0 (.DIODE(net709));
 sky130_fd_sc_hd__diode_2 ANTENNA_c679_S1 (.DIODE(net709));
 sky130_fd_sc_hd__diode_2 ANTENNA_c678_A3 (.DIODE(net709));
 sky130_fd_sc_hd__diode_2 ANTENNA_c676_S1 (.DIODE(net709));
 sky130_fd_sc_hd__diode_2 ANTENNA_s928_Q (.DIODE(net710));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_S1 (.DIODE(net710));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_S0 (.DIODE(net710));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_S1 (.DIODE(net710));
 sky130_fd_sc_hd__diode_2 ANTENNA_c685_S1 (.DIODE(net710));
 sky130_fd_sc_hd__diode_2 ANTENNA_c678_S0 (.DIODE(net710));
 sky130_fd_sc_hd__diode_2 ANTENNA_s934_Q (.DIODE(net719));
 sky130_fd_sc_hd__diode_2 ANTENNA_c759_S1 (.DIODE(net719));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_S1 (.DIODE(net719));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_S1 (.DIODE(net719));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_A0 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_A3 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_A1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_A2 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_A2 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_c238_A2 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_B1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_X (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_A0 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_A2 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_S0 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_A0 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_c215_X (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone37_A (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout216_A (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_A1 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c134_X (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_A3 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_S1 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_A2 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_A0 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_c370_A1 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_A1 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_X (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_A1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_A3 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_c240_A1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_c238_A1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_S1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_c229_A0 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_c226_X (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_A2 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_c496_A1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_c239_A1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_c234_A0 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_A2 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_c229_A1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_c228_S1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_X (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_c427_A2 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_A1 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c278_A3 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_A1 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c266_A4 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_A2 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_A2 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_A1 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_A1 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c136_X (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c760_A0 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_c633_A1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_A3 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_A3 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_c232_A1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_c230_X (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout259_A (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_X (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_A2 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_S1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout248_A (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_X (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_A2 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout247_A (.DIODE(net724));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_X (.DIODE(net724));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_S0 (.DIODE(net724));
 sky130_fd_sc_hd__diode_2 ANTENNA_c271_A3 (.DIODE(net724));
 sky130_fd_sc_hd__diode_2 ANTENNA_c267_A4 (.DIODE(net724));
 sky130_fd_sc_hd__diode_2 ANTENNA_c266_A1 (.DIODE(net724));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_X (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA_c428_A0 (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_B1 (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA_c413_A0 (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA_c401_A1 (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_A4 (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_B1 (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA_c265_A2 (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_S1 (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_A2 (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_A2 (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout243_A (.DIODE(net726));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_X (.DIODE(net726));
 sky130_fd_sc_hd__diode_2 ANTENNA_c685_A2 (.DIODE(net726));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_X (.DIODE(net727));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_A0 (.DIODE(net727));
 sky130_fd_sc_hd__diode_2 ANTENNA_c212_A3 (.DIODE(net727));
 sky130_fd_sc_hd__diode_2 ANTENNA_c208_A1 (.DIODE(net727));
 sky130_fd_sc_hd__diode_2 ANTENNA_c180_S0 (.DIODE(net727));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_A1 (.DIODE(net727));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_B1 (.DIODE(net727));
 sky130_fd_sc_hd__diode_2 ANTENNA_c130_A1 (.DIODE(net727));
 sky130_fd_sc_hd__diode_2 ANTENNA_c123_A0 (.DIODE(net727));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout238_A (.DIODE(net728));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_X (.DIODE(net728));
 sky130_fd_sc_hd__diode_2 ANTENNA_c759_A0 (.DIODE(net728));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_A2 (.DIODE(net728));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_S0 (.DIODE(net728));
 sky130_fd_sc_hd__diode_2 ANTENNA_c660_A1 (.DIODE(net728));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout234_A (.DIODE(net729));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_X (.DIODE(net729));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_A1 (.DIODE(net729));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_A3 (.DIODE(net729));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout258_A (.DIODE(net731));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_X (.DIODE(net731));
 sky130_fd_sc_hd__diode_2 ANTENNA_c674_A1 (.DIODE(net731));
 sky130_fd_sc_hd__diode_2 ANTENNA_c662_A3 (.DIODE(net731));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone19_A (.DIODE(net732));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout257_A (.DIODE(net732));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_X (.DIODE(net732));
 sky130_fd_sc_hd__diode_2 ANTENNA_c744_A1 (.DIODE(net732));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout254_A (.DIODE(net733));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout253_A (.DIODE(net733));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_X (.DIODE(net733));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout252_A (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout251_A (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_X (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_X (.DIODE(net735));
 sky130_fd_sc_hd__diode_2 ANTENNA_c529_A1 (.DIODE(net735));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_A2 (.DIODE(net735));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_A0 (.DIODE(net735));
 sky130_fd_sc_hd__diode_2 ANTENNA_c405_A1 (.DIODE(net735));
 sky130_fd_sc_hd__diode_2 ANTENNA_c398_A1 (.DIODE(net735));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_A1 (.DIODE(net735));
 sky130_fd_sc_hd__diode_2 ANTENNA_c286_A3 (.DIODE(net735));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_A3 (.DIODE(net735));
 sky130_fd_sc_hd__diode_2 ANTENNA_c134_B1 (.DIODE(net735));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout250_A (.DIODE(net736));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_X (.DIODE(net736));
 sky130_fd_sc_hd__diode_2 ANTENNA_c744_A2 (.DIODE(net736));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_S1 (.DIODE(net736));
 sky130_fd_sc_hd__diode_2 ANTENNA_c680_A2 (.DIODE(net736));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_X (.DIODE(net737));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_A0 (.DIODE(net737));
 sky130_fd_sc_hd__diode_2 ANTENNA_c558_S0 (.DIODE(net737));
 sky130_fd_sc_hd__diode_2 ANTENNA_c557_A3 (.DIODE(net737));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_A3 (.DIODE(net737));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_S1 (.DIODE(net737));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_A1 (.DIODE(net737));
 sky130_fd_sc_hd__diode_2 ANTENNA_c235_A3 (.DIODE(net737));
 sky130_fd_sc_hd__diode_2 ANTENNA_c198_A3 (.DIODE(net737));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_A2 (.DIODE(net737));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_X (.DIODE(net738));
 sky130_fd_sc_hd__diode_2 ANTENNA_c502_A0 (.DIODE(net738));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_A1 (.DIODE(net738));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_A0 (.DIODE(net738));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_A2 (.DIODE(net738));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_A0 (.DIODE(net738));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_A1 (.DIODE(net738));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_A2 (.DIODE(net738));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_A3 (.DIODE(net738));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_A3 (.DIODE(net738));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout249_A (.DIODE(net739));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_X (.DIODE(net739));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_A2 (.DIODE(net739));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_A2 (.DIODE(net739));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_A0 (.DIODE(net739));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_A1 (.DIODE(net739));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_X (.DIODE(net740));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_A3 (.DIODE(net740));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_A3 (.DIODE(net740));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_A1 (.DIODE(net740));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_A1 (.DIODE(net740));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_S0 (.DIODE(net740));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_A4 (.DIODE(net740));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_A3 (.DIODE(net740));
 sky130_fd_sc_hd__diode_2 ANTENNA_c100_A0 (.DIODE(net740));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_X (.DIODE(net741));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_A0 (.DIODE(net741));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_A3 (.DIODE(net741));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_A2 (.DIODE(net741));
 sky130_fd_sc_hd__diode_2 ANTENNA_c701_A2 (.DIODE(net741));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_A3 (.DIODE(net741));
 sky130_fd_sc_hd__diode_2 ANTENNA_c587_A3 (.DIODE(net741));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_A3 (.DIODE(net741));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_S1 (.DIODE(net741));
 sky130_fd_sc_hd__diode_2 ANTENNA_c295_S0 (.DIODE(net741));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_A1 (.DIODE(net741));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_X (.DIODE(net742));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_A0 (.DIODE(net742));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_A0 (.DIODE(net742));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_A0 (.DIODE(net742));
 sky130_fd_sc_hd__diode_2 ANTENNA_c430_A2 (.DIODE(net742));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_A1 (.DIODE(net742));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_A3 (.DIODE(net742));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_A3 (.DIODE(net742));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_A3 (.DIODE(net742));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_X (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_S0 (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_A0 (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA_c183_A3 (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_S1 (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_A2 (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_A4 (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_B1 (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_X (.DIODE(net744));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_A0 (.DIODE(net744));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_A2 (.DIODE(net744));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_A2 (.DIODE(net744));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_A0 (.DIODE(net744));
 sky130_fd_sc_hd__diode_2 ANTENNA_c431_SCD (.DIODE(net744));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_A1 (.DIODE(net744));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_A3 (.DIODE(net744));
 sky130_fd_sc_hd__diode_2 ANTENNA_c311_A1 (.DIODE(net744));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_B1 (.DIODE(net744));
 sky130_fd_sc_hd__diode_2 ANTENNA_c159_A4 (.DIODE(net744));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_A4 (.DIODE(net745));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_X (.DIODE(net745));
 sky130_fd_sc_hd__diode_2 ANTENNA_c668_A0 (.DIODE(net745));
 sky130_fd_sc_hd__diode_2 ANTENNA_c663_S1 (.DIODE(net745));
 sky130_fd_sc_hd__diode_2 ANTENNA_c662_A2 (.DIODE(net745));
 sky130_fd_sc_hd__diode_2 ANTENNA_c543_A2 (.DIODE(net745));
 sky130_fd_sc_hd__diode_2 ANTENNA_c403_A2 (.DIODE(net745));
 sky130_fd_sc_hd__diode_2 ANTENNA_c400_RESET_B (.DIODE(net745));
 sky130_fd_sc_hd__diode_2 ANTENNA_c267_A1 (.DIODE(net745));
 sky130_fd_sc_hd__diode_2 ANTENNA_c136_A1 (.DIODE(net745));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_X (.DIODE(net746));
 sky130_fd_sc_hd__diode_2 ANTENNA_c366_A1 (.DIODE(net746));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_A1 (.DIODE(net746));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_A1 (.DIODE(net746));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_A4 (.DIODE(net746));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_B1 (.DIODE(net746));
 sky130_fd_sc_hd__diode_2 ANTENNA_c102_A1 (.DIODE(net746));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_X (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA_c191_A0 (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_A3 (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_A2 (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_A1 (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_A2 (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_X (.DIODE(net748));
 sky130_fd_sc_hd__diode_2 ANTENNA_c742_A3 (.DIODE(net748));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_A1 (.DIODE(net748));
 sky130_fd_sc_hd__diode_2 ANTENNA_c615_A3 (.DIODE(net748));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_A1 (.DIODE(net748));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_A0 (.DIODE(net748));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_A3 (.DIODE(net748));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_A1 (.DIODE(net748));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_S0 (.DIODE(net748));
 sky130_fd_sc_hd__diode_2 ANTENNA_c215_A2 (.DIODE(net748));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_A4 (.DIODE(net748));
 sky130_fd_sc_hd__diode_2 ANTENNA_input28_X (.DIODE(net749));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_A0 (.DIODE(net749));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_B1 (.DIODE(net749));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_B1 (.DIODE(net749));
 sky130_fd_sc_hd__diode_2 ANTENNA_c234_A3 (.DIODE(net749));
 sky130_fd_sc_hd__diode_2 ANTENNA_c205_A3 (.DIODE(net749));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_A1 (.DIODE(net749));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_A0 (.DIODE(net749));
 sky130_fd_sc_hd__diode_2 ANTENNA_c129_A1 (.DIODE(net749));
 sky130_fd_sc_hd__diode_2 ANTENNA_input29_X (.DIODE(net750));
 sky130_fd_sc_hd__diode_2 ANTENNA_c458_A0 (.DIODE(net750));
 sky130_fd_sc_hd__diode_2 ANTENNA_c424_A1 (.DIODE(net750));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_A2 (.DIODE(net750));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_A2 (.DIODE(net750));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_S0 (.DIODE(net750));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_A3 (.DIODE(net750));
 sky130_fd_sc_hd__diode_2 ANTENNA_c180_A1 (.DIODE(net750));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_A2 (.DIODE(net750));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_A3 (.DIODE(net750));
 sky130_fd_sc_hd__diode_2 ANTENNA_input30_X (.DIODE(net751));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_A0 (.DIODE(net751));
 sky130_fd_sc_hd__diode_2 ANTENNA_c286_A1 (.DIODE(net751));
 sky130_fd_sc_hd__diode_2 ANTENNA_c205_A2 (.DIODE(net751));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_A2 (.DIODE(net751));
 sky130_fd_sc_hd__diode_2 ANTENNA_c129_A0 (.DIODE(net751));
 sky130_fd_sc_hd__diode_2 ANTENNA_input31_X (.DIODE(net752));
 sky130_fd_sc_hd__diode_2 ANTENNA_c230_A1 (.DIODE(net752));
 sky130_fd_sc_hd__diode_2 ANTENNA_c205_A1 (.DIODE(net752));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_A1 (.DIODE(net752));
 sky130_fd_sc_hd__diode_2 ANTENNA_c158_A3 (.DIODE(net752));
 sky130_fd_sc_hd__diode_2 ANTENNA_input32_X (.DIODE(net753));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_A1 (.DIODE(net753));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A3 (.DIODE(net753));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_A2 (.DIODE(net753));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_A2 (.DIODE(net753));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_A3 (.DIODE(net753));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_A2 (.DIODE(net753));
 sky130_fd_sc_hd__diode_2 ANTENNA_c313_A3 (.DIODE(net753));
 sky130_fd_sc_hd__diode_2 ANTENNA_c182_A1 (.DIODE(net753));
 sky130_fd_sc_hd__diode_2 ANTENNA_input33_X (.DIODE(net754));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_A1 (.DIODE(net754));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_A1 (.DIODE(net754));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_A2 (.DIODE(net754));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_A1 (.DIODE(net754));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_S0 (.DIODE(net754));
 sky130_fd_sc_hd__diode_2 ANTENNA_c340_S0 (.DIODE(net754));
 sky130_fd_sc_hd__diode_2 ANTENNA_c231_A0 (.DIODE(net754));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_S0 (.DIODE(net754));
 sky130_fd_sc_hd__diode_2 ANTENNA_input34_X (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA_c739_S0 (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_A2 (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_A1 (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_A0 (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_A3 (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_A2 (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_A2 (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA_input36_X (.DIODE(net757));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_A2 (.DIODE(net757));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_A0 (.DIODE(net757));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_A2 (.DIODE(net757));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_A3 (.DIODE(net757));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_A0 (.DIODE(net757));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_S0 (.DIODE(net757));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_S1 (.DIODE(net757));
 sky130_fd_sc_hd__diode_2 ANTENNA_c180_A2 (.DIODE(net757));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_S0 (.DIODE(net757));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_S0 (.DIODE(net757));
 sky130_fd_sc_hd__diode_2 ANTENNA_input37_X (.DIODE(net758));
 sky130_fd_sc_hd__diode_2 ANTENNA_c371_A3 (.DIODE(net758));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_A1 (.DIODE(net758));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_A2 (.DIODE(net758));
 sky130_fd_sc_hd__diode_2 ANTENNA_c124_A0 (.DIODE(net758));
 sky130_fd_sc_hd__diode_2 ANTENNA_input38_X (.DIODE(net759));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_A0 (.DIODE(net759));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_A0 (.DIODE(net759));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_A2 (.DIODE(net759));
 sky130_fd_sc_hd__diode_2 ANTENNA_c191_A1 (.DIODE(net759));
 sky130_fd_sc_hd__diode_2 ANTENNA_c158_A2 (.DIODE(net759));
 sky130_fd_sc_hd__diode_2 ANTENNA_input39_X (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA_c760_A1 (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA_c759_A3 (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_A2 (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_A2 (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_A2 (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA_c566_A1 (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_A3 (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA_c228_A3 (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA_c203_A0 (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA_input40_X (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_A3 (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_A1 (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_A0 (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_A1 (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_A2 (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_S0 (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_c222_A3 (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_c194_A2 (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_S0 (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_input41_X (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_A0 (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_A1 (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_A2 (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_A1 (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA_input43_X (.DIODE(net764));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_A2 (.DIODE(net764));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_A0 (.DIODE(net764));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_B1 (.DIODE(net764));
 sky130_fd_sc_hd__diode_2 ANTENNA_c183_S1 (.DIODE(net764));
 sky130_fd_sc_hd__diode_2 ANTENNA_input44_X (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_A4 (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_A3 (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_c124_A1 (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_c122_A3 (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_input48_X (.DIODE(net769));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_A2 (.DIODE(net769));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_A1 (.DIODE(net769));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_A1 (.DIODE(net769));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_A0 (.DIODE(net769));
 sky130_fd_sc_hd__diode_2 ANTENNA_c203_A2 (.DIODE(net769));
 sky130_fd_sc_hd__diode_2 ANTENNA_input50_X (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_c368_A2 (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_c346_A2 (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_A0 (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_A1 (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_c206_A2 (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_A3 (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_c184_A1 (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_c183_S0 (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_c127_A0 (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_c122_A2 (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_input51_X (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_A0 (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_A3 (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_c191_A2 (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_c182_A2 (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_input52_X (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_A0 (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_A2 (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_S1 (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout242_A (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_input53_X (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_A2 (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_S0 (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_A0 (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_input54_X (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_c228_A0 (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_c206_A1 (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_A3 (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_B1 (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_c102_S1 (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_input55_X (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_A1 (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_A0 (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_A2 (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_A1 (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_A2 (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_S0 (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c190_A1 (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_A2 (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c131_S1 (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c124_S0 (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout241_A (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_input56_X (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_c757_A0 (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_A2 (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout240_A (.DIODE(net778));
 sky130_fd_sc_hd__diode_2 ANTENNA_input57_X (.DIODE(net778));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_S0 (.DIODE(net778));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_A1 (.DIODE(net778));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_S0 (.DIODE(net778));
 sky130_fd_sc_hd__diode_2 ANTENNA_input58_X (.DIODE(net779));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_A3 (.DIODE(net779));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_A2 (.DIODE(net779));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_A0 (.DIODE(net779));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_A4 (.DIODE(net779));
 sky130_fd_sc_hd__diode_2 ANTENNA_input59_X (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_A2 (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_A1 (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_A4 (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA_c129_S0 (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA_c124_A3 (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA_input64_X (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_A0 (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_S0 (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_c236_A0 (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_A3 (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_c130_A3 (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_c128_A2 (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_c122_A1 (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_c109_S1 (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_input67_X (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_A0 (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_A1 (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_A1 (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout239_A (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_input68_X (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_c723_A2 (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_c720_A0 (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_A0 (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout237_A (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_input70_X (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_A1 (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_S0 (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_A2 (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_input74_X (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_c239_A0 (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_c215_S1 (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_c106_A2 (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout235_A (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_input79_X (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c759_A1 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A2 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_A2 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_input80_X (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_A0 (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_A2 (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_A3 (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_A2 (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_A3 (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_S1 (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_c344_S0 (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_A1 (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_A2 (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_c216_A2 (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_input81_X (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_A0 (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_A0 (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_A2 (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_B1 (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_c123_A2 (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_c107_A1 (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_c106_A3 (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_c103_A1 (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_input83_X (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c231_A2 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_A3 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_input84_X (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_A1 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_A0 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_c340_A1 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_input88_X (.DIODE(net809));
 sky130_fd_sc_hd__diode_2 ANTENNA_c494_A1 (.DIODE(net809));
 sky130_fd_sc_hd__diode_2 ANTENNA_c128_S0 (.DIODE(net809));
 sky130_fd_sc_hd__diode_2 ANTENNA_c106_A1 (.DIODE(net809));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout230_A (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout229_A (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_input90_X (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_A2 (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_A1 (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_input92_X (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c373_A0 (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c368_A3 (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_A2 (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_A1 (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c105_S0 (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c100_S1 (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_input93_X (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_c633_A2 (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_A0 (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_A0 (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_c373_A2 (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_c109_S0 (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_c101_A3 (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_input94_X (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_c365_A1 (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_c107_A3 (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_c104_A1 (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_c102_A0 (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_input96_X (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_A3 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_S1 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_A0 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_A3 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c103_S1 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_input97_X (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_A0 (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c107_A2 (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c105_A3 (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c104_A3 (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c100_A2 (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_input100_X (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_c372_A2 (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_c123_S0 (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_c104_A2 (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_c100_S0 (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone17_A (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout212_A (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout211_A (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_X (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_output104_A (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge793_Q_N (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_S0 (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout172_A (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_output105_A (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_A2 (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_S0 (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_c297_X (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_output106_A (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_s919_Q (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_S1 (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_S1 (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_output107_A (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_A2 (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_A0 (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_A3 (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_c372_S0 (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_c350_A2 (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_A0 (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_c340_A2 (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_X (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_output108_A (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_A2 (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_S0 (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_A0 (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_A2 (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_A2 (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_A2 (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_X (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_output109_A (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_A3 (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_S1 (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_A1 (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_A2 (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_A1 (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA_c446_A2 (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_X (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA_output110_A (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_s912_Q (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_S1 (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_S1 (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c571_S0 (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_S0 (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c566_S0 (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c564_S1 (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c563_S1 (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c560_S1 (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_output111_A (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_A2 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_A2 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_A3 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_S0 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_A0 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_A1 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_X (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_output112_A (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_c411_A2 (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_A2 (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_c369_A1 (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_A1 (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_c278_X (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_output114_A (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge845_Q (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_A3 (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_S0 (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_S1 (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c350_S0 (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_A3 (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_A2 (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_A3 (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout207_A (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_A3 (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_A1 (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_X (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_output120_A (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_A1 (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_A1 (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_A0 (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_A2 (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_c275_X (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_output121_A (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_A0 (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_A1 (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_c369_A2 (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_A2 (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_A1 (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_S1 (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_X (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout223_A (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge795_Q (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_S0 (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_c557_S1 (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_output125_A (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_S0 (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_S0 (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_S0 (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_c364_A2 (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_A1 (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_X (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_output126_A (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_s887_Q (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_S1 (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_S0 (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_c437_S0 (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_c434_S0 (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_c428_S1 (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_output127_A (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_A2 (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_A1 (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_X (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_output128_A (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_A2 (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c370_A2 (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c237_S0 (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c221_A1 (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c216_A1 (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c215_A1 (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_X (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_output131_A (.DIODE(net1055));
 sky130_fd_sc_hd__diode_2 ANTENNA_c536_A2 (.DIODE(net1054));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_A3 (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_A1 (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_A2 (.DIODE(net1053));
 sky130_fd_sc_hd__diode_2 ANTENNA_c283_A1 (.DIODE(net1053));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_A0 (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_S1 (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_X (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_output137_A (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_c364_A1 (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_A2 (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_A3 (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_X (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_output138_A (.DIODE(net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_A0 (.DIODE(net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_A1 (.DIODE(net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_A0 (.DIODE(net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_c365_A3 (.DIODE(net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_c236_A1 (.DIODE(net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_A1 (.DIODE(net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_c222_X (.DIODE(net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_output142_A (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_A1 (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_c125_A2 (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_c103_S0 (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_c101_X (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_output143_A (.DIODE(net864));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_A2 (.DIODE(net864));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_A3 (.DIODE(net864));
 sky130_fd_sc_hd__diode_2 ANTENNA_c350_A3 (.DIODE(net864));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_A0 (.DIODE(net864));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_A0 (.DIODE(net864));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_X (.DIODE(net864));
 sky130_fd_sc_hd__diode_2 ANTENNA_output144_A (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge824_Q (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c458_S0 (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c446_S0 (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_A3 (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_S0 (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_S1 (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_S1 (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_A4 (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_output148_A (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge834_Q (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_A3 (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_S1 (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_A3 (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_output150_A (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA_c237_A2 (.DIODE(net1052));
 sky130_fd_sc_hd__diode_2 ANTENNA_c230_A3 (.DIODE(net1052));
 sky130_fd_sc_hd__diode_2 ANTENNA_c203_S0 (.DIODE(net1052));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_A1 (.DIODE(net1052));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_A0 (.DIODE(net1052));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_A4 (.DIODE(net1052));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_A4 (.DIODE(net1052));
 sky130_fd_sc_hd__diode_2 ANTENNA_c148_X (.DIODE(net1052));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone36_A (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout209_A (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_output151_A (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_c140_X (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_output153_A (.DIODE(net1045));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_A4 (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_c198_A1 (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_A2 (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_c183_A1 (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_S0 (.DIODE(net1044));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_A0 (.DIODE(net1045));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_S0 (.DIODE(net1046));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_X (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_output159_A (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge801_Q (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_S0 (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c482_S0 (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_S1 (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_A3 (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c218_S0 (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c212_S1 (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_S1 (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_output160_A (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_A3 (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_A2 (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c194_S1 (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_S0 (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_A1 (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_A0 (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_X (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_output163_A (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_c577_A2 (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_A1 (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_A2 (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_c431_Q (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout168_X (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c663_A2 (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c543_A3 (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c536_A3 (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c537_RESET_B (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout167_A (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c545_A0 (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c535_S1 (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c533_SCD (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c531_A3 (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c530_A3 (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout169_X (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_A0 (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_A1 (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_A1 (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c321_A2 (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_S0 (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_A2 (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c344_A3 (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c340_S1 (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_S0 (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_S1 (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout170_X (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_A0 (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_A2 (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_A1 (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_A1 (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout169_A (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout171_X (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_A2 (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_S0 (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_A3 (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_A3 (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_A1 (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_A1 (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_S0 (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_A3 (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_A2 (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_A3 (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout172_X (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_A3 (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_A2 (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c424_S1 (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_A3 (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout171_A (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout173_X (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c406_S0 (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c541_A3 (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c564_A0 (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c409_A1 (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c535_A1 (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_A2 (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_A4 (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c414_A3 (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c413_A2 (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c410_S1 (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout174_X (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_c662_A0 (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_c661_A3 (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_c739_A0 (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_S0 (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_A3 (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_A3 (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_S1 (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_c546_A1 (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_A2 (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_A2 (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout175_X (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_A3 (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_A4 (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_A2 (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_A3 (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_A1 (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_A1 (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_A3 (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_S1 (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_S1 (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_S1 (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout176_X (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_A1 (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_A1 (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c561_A1 (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_A1 (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_A3 (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c321_S0 (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_A1 (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_A2 (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_A4 (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_A2 (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout177_X (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_A1 (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_A0 (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_A1 (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_A1 (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_S0 (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_A3 (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c297_A4 (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c295_A3 (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_A3 (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_A2 (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout180_X (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_c427_A1 (.DIODE(net1064));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_A0 (.DIODE(net1064));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_A3 (.DIODE(net1064));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_S1 (.DIODE(net1064));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_A2 (.DIODE(net1064));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout181_X (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_A1 (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_B1 (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_A1 (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_A2 (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_c372_A3 (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_A3 (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_A3 (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_A2 (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_c222_A1 (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_c205_S0 (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout182_X (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_output122_A (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_A2 (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_S0 (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_A3 (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_A4 (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout183_X (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_A3 (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c232_A0 (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_A1 (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_A3 (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c194_A0 (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_A3 (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_S0 (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c184_S0 (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c182_A3 (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c183_A2 (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout184_X (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c275_A2 (.DIODE(net1063));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_A3 (.DIODE(net1063));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_A2 (.DIODE(net1063));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_A1 (.DIODE(net1063));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_A0 (.DIODE(net1063));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout185_X (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_c693_A0 (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_c406_S1 (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_c413_A3 (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_c412_A1 (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_c405_S1 (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_c404_A1 (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_c403_A4 (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_c402_B1 (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_c401_A2 (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_S0 (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout186_X (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_c558_A1 (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout185_A (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_c761_S0 (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_A0 (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_A3 (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_A3 (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_A3 (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_A3 (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_A3 (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_S0 (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout187_X (.DIODE(net1058));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_S1 (.DIODE(net1058));
 sky130_fd_sc_hd__diode_2 ANTENNA_c203_A3 (.DIODE(net1058));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_B1 (.DIODE(net1058));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_A2 (.DIODE(net1058));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_S1 (.DIODE(net1058));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout188_X (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_c742_A0 (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_c723_A1 (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_A3 (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_c664_A2 (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_A3 (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_A1 (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout190_X (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_c404_S0 (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout189_A (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_c277_A0 (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_A4 (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_c275_B1 (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout191_X (.DIODE(net912));
 sky130_fd_sc_hd__diode_2 ANTENNA_c673_A1 (.DIODE(net912));
 sky130_fd_sc_hd__diode_2 ANTENNA_c678_A1 (.DIODE(net912));
 sky130_fd_sc_hd__diode_2 ANTENNA_c675_S0 (.DIODE(net912));
 sky130_fd_sc_hd__diode_2 ANTENNA_c670_A3 (.DIODE(net912));
 sky130_fd_sc_hd__diode_2 ANTENNA_c667_S0 (.DIODE(net912));
 sky130_fd_sc_hd__diode_2 ANTENNA_c665_A3 (.DIODE(net912));
 sky130_fd_sc_hd__diode_2 ANTENNA_c555_S1 (.DIODE(net912));
 sky130_fd_sc_hd__diode_2 ANTENNA_c528_A4 (.DIODE(net912));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout190_A (.DIODE(net912));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout192_X (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout191_A (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_S0 (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A0 (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_A2 (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_A1 (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout193_X (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_A1 (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA_c274_A2 (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA_c273_A2 (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA_c271_A4 (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA_c269_B1 (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_A0 (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA_c368_A0 (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_S0 (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_A3 (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_A1 (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout194_X (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_c399_A2 (.DIODE(net1060));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_A3 (.DIODE(net1060));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_A1 (.DIODE(net1060));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_A1 (.DIODE(net1060));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_A2 (.DIODE(net1060));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout197_X (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_output141_A (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_A1 (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_c411_A1 (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_c410_A1 (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_c398_A3 (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_c267_A2 (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout195_A (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout196_A (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout198_X (.DIODE(net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout197_A (.DIODE(net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_A2 (.DIODE(net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_A2 (.DIODE(net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_A3 (.DIODE(net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_S1 (.DIODE(net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_c275_A3 (.DIODE(net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone38_A (.DIODE(net1086));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout200_X (.DIODE(net1086));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_S1 (.DIODE(net1086));
 sky130_fd_sc_hd__diode_2 ANTENNA_c408_A3 (.DIODE(net1086));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout199_A (.DIODE(net1086));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_S1 (.DIODE(net1086));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_S0 (.DIODE(net1086));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_A2 (.DIODE(net1086));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout201_X (.DIODE(net1077));
 sky130_fd_sc_hd__diode_2 ANTENNA_c669_A1 (.DIODE(net1056));
 sky130_fd_sc_hd__diode_2 ANTENNA_c664_S0 (.DIODE(net1056));
 sky130_fd_sc_hd__diode_2 ANTENNA_c424_A3 (.DIODE(net1056));
 sky130_fd_sc_hd__diode_2 ANTENNA_c746_A0 (.DIODE(net1056));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_A1 (.DIODE(net1056));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_A1 (.DIODE(net1056));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_A0 (.DIODE(net1056));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout200_A (.DIODE(net1056));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout202_X (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c663_A1 (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_A2 (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_A1 (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_A2 (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_A1 (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_A3 (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c283_A3 (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c275_A4 (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c267_A3 (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c159_A1 (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer24_A (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer22_A (.DIODE(net1061));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout206_X (.DIODE(net1061));
 sky130_fd_sc_hd__diode_2 ANTENNA_c680_A3 (.DIODE(net1061));
 sky130_fd_sc_hd__diode_2 ANTENNA_c405_A2 (.DIODE(net1061));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_A2 (.DIODE(net1061));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_A1 (.DIODE(net1061));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout207_X (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_A1 (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c194_S0 (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_A0 (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_output118_A (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_A1 (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_A2 (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_A2 (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_A1 (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_S1 (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c226_A3 (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout210_X (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_c693_A1 (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_c668_A3 (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_c667_A2 (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_c663_S0 (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_c661_A1 (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_c586_A1 (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_c555_S0 (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_c397_A1 (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_c321_A1 (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_A1 (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_A2 (.DIODE(net1059));
 sky130_fd_sc_hd__diode_2 ANTENNA_c140_A1 (.DIODE(net1059));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout211_X (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_A2 (.DIODE(net1059));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_A1 (.DIODE(net1059));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_A2 (.DIODE(net1059));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout212_X (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_output101_A (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c540_A3 (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c528_A1 (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_A3 (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_A3 (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c400_SCE (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout213_X (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c397_A2 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c537_SCD (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c313_S0 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c276_A1 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c274_A1 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c272_A3 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c269_A3 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_A2 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c535_A2 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c399_B1 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout214_X (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_A1 (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c687_A3 (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout213_A (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c760_S1 (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A0 (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_A3 (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout215_X (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c577_S0 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_A1 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_A1 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c430_A3 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_A3 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_A1 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_A2 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_A3 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_A0 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_S0 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_A1 (.DIODE(net1062));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout216_X (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_A3 (.DIODE(net1062));
 sky130_fd_sc_hd__diode_2 ANTENNA_c138_A2 (.DIODE(net1062));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_A1 (.DIODE(net1062));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_A0 (.DIODE(net1062));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap217_X (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_c743_A3 (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_S0 (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_A2 (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_S0 (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_S1 (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_S1 (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap218_X (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c744_S0 (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_S0 (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_A3 (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout219_X (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_c564_S0 (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_S0 (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_A3 (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_c687_S1 (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_S0 (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_B1 (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_S1 (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_S1 (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_S1 (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_S1 (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold58_A (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap220_X (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c703_A2 (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_A3 (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_S1 (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c538_A3 (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout221_X (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_S0 (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_S1 (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_A4 (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_S0 (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_S1 (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_S1 (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_S0 (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_A2 (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_S0 (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_S0 (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout222_X (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c205_S1 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c230_S1 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c235_S1 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c232_S0 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c229_S1 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_S1 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c221_S0 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c220_S0 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c218_A3 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_S0 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout223_X (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_S0 (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_S0 (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_B1 (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_S1 (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_output124_A (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_S0 (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_A3 (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_S0 (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_c206_S0 (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_S1 (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout224_X (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_c561_A2 (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_c557_S0 (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_c556_S0 (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_S0 (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_S0 (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_B1 (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_S0 (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_S0 (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_S1 (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_S0 (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout225_X (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c674_A3 (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c672_A3 (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c663_A3 (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c554_A2 (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_A2 (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c412_A2 (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c411_A3 (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c406_A2 (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c404_A2 (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c401_A4 (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout226_X (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c415_S0 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c410_A2 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c405_A0 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c403_A3 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c402_A3 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_A2 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c763_A1 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c494_A2 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_A1 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_A1 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone16_A1 (.DIODE(net1084));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_A1 (.DIODE(net1084));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout227_X (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c264_A2 (.DIODE(net1084));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_S0 (.DIODE(net1084));
 sky130_fd_sc_hd__diode_2 ANTENNA_c180_S1 (.DIODE(net1084));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout229_X (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_S1 (.DIODE(net1083));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_A3 (.DIODE(net1083));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout228_A (.DIODE(net1083));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_A4 (.DIODE(net1083));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_A1 (.DIODE(net1083));
 sky130_fd_sc_hd__diode_2 ANTENNA_c126_S1 (.DIODE(net1083));
 sky130_fd_sc_hd__diode_2 ANTENNA_c124_S1 (.DIODE(net1083));
 sky130_fd_sc_hd__diode_2 ANTENNA_c122_S0 (.DIODE(net1083));
 sky130_fd_sc_hd__diode_2 ANTENNA_c107_S1 (.DIODE(net1083));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout230_X (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_c679_A1 (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_c676_A2 (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_c668_S0 (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_c664_A3 (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_c547_A1 (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_c530_A2 (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_c529_A4 (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_c401_B1 (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_A2 (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_A1 (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_A2 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout231_X (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_A4 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_A0 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_B1 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c138_B1 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_A3 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c311_A3 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_A3 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_S1 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_B1 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout232_X (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c666_A1 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c662_A1 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c660_S0 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c537_D (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c534_A1 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c531_S0 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_A3 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A3 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c614_A1 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_S0 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout233_X (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c668_S1 (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c673_A4 (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c686_A2 (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout232_A (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c159_B1 (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c265_B1 (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_S0 (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c270_S1 (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout231_A (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout234_X (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_c667_A0 (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_c562_A2 (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_S0 (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_c403_A1 (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_c407_A2 (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_c398_A2 (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_A3 (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_A2 (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_A1 (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_S0 (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout235_X (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_S0 (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_A1 (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_S1 (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_A3 (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_A2 (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_A3 (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_A2 (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_A0 (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_c180_A3 (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_c107_S0 (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout236_X (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_A0 (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_S0 (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_A1 (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_S0 (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_A2 (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_S1 (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_A2 (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_A3 (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c368_A1 (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c232_A2 (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout237_X (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_A1 (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_S1 (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_A3 (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_A0 (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_S0 (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c230_A2 (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_A1 (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c212_A1 (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_A2 (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c108_A3 (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_A3 (.DIODE(net1081));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout238_X (.DIODE(net1081));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_S0 (.DIODE(net1081));
 sky130_fd_sc_hd__diode_2 ANTENNA_c611_A3 (.DIODE(net1081));
 sky130_fd_sc_hd__diode_2 ANTENNA_c610_A2 (.DIODE(net1081));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_A3 (.DIODE(net1081));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_A0 (.DIODE(net1081));
 sky130_fd_sc_hd__diode_2 ANTENNA_c279_A2 (.DIODE(net1081));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_A3 (.DIODE(net1081));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_A3 (.DIODE(net1081));
 sky130_fd_sc_hd__diode_2 ANTENNA_c134_A2 (.DIODE(net1081));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout5_A (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone16_A2 (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout239_X (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout240_X (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A2 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_A3 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_A3 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_A2 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_A3 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_A0 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_A4 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_A3 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_A0 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_A3 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout241_X (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_A1 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_A1 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_A2 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_A2 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c587_A0 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_A3 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_A3 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_A2 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_S1 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_A3 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout242_X (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_A3 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_S0 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_A2 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_A3 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_A2 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_A1 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_S1 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_A3 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_S0 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_A2 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout243_X (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_A0 (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c667_A1 (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c663_A0 (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c556_A1 (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c532_A3 (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_S1 (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_A1 (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_S0 (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c270_A3 (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c138_A1 (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c140_A4 (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout244_X (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c264_A3 (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c143_A3 (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_A4 (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_A4 (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c134_A4 (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_A3 (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_A3 (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c297_B1 (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_A3 (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout245_X (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c679_A3 (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c665_A1 (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c556_A2 (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c528_A3 (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c265_A1 (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c267_B1 (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c270_S0 (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c535_S0 (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout244_A (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout246_X (.DIODE(net1080));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout245_A (.DIODE(net1080));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_A0 (.DIODE(net1080));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_A3 (.DIODE(net1080));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_A3 (.DIODE(net1080));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_A3 (.DIODE(net1080));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_A2 (.DIODE(net1080));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_A0 (.DIODE(net1080));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_A3 (.DIODE(net1080));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_A4 (.DIODE(net1080));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout247_X (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_S0 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_B1 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_A2 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_A0 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_A2 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c496_A3 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_A1 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_A3 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_A0 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c125_S1 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout4_A (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone16_A3 (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout248_X (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout249_X (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_A2 (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_A2 (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_A1 (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_A3 (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_c286_A2 (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_c212_S0 (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_S0 (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_A2 (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_B1 (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_A2 (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout250_X (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_c529_A3 (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_S1 (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_S0 (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_c408_A0 (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_c405_A3 (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_c278_A0 (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_A0 (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_A2 (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_A3 (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_A2 (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout251_X (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_A1 (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_S0 (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_A1 (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c537_SCE (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c397_A4 (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c535_A3 (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_A3 (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_A4 (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c140_A2 (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c102_S0 (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout252_X (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_c762_A1 (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_A3 (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_A1 (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_A3 (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_A3 (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_A2 (.DIODE(net1079));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_S0 (.DIODE(net1079));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_A1 (.DIODE(net1079));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_A1 (.DIODE(net1079));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_A1 (.DIODE(net1079));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout253_X (.DIODE(net1079));
 sky130_fd_sc_hd__diode_2 ANTENNA_c140_B1 (.DIODE(net1079));
 sky130_fd_sc_hd__diode_2 ANTENNA_c230_A0 (.DIODE(net1079));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_A2 (.DIODE(net1079));
 sky130_fd_sc_hd__diode_2 ANTENNA_c215_S0 (.DIODE(net1079));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_A2 (.DIODE(net1079));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout254_X (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c547_A2 (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c540_A1 (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c530_A0 (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_A3 (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c266_A3 (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_A2 (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_A1 (.DIODE(net1078));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout256_X (.DIODE(net1078));
 sky130_fd_sc_hd__diode_2 ANTENNA_c274_B1 (.DIODE(net1078));
 sky130_fd_sc_hd__diode_2 ANTENNA_c313_S1 (.DIODE(net1078));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout255_A (.DIODE(net1078));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_A1 (.DIODE(net1078));
 sky130_fd_sc_hd__diode_2 ANTENNA_c446_A3 (.DIODE(net1078));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_S0 (.DIODE(net1078));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_A2 (.DIODE(net1078));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer39_A (.DIODE(net1082));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout257_X (.DIODE(net1082));
 sky130_fd_sc_hd__diode_2 ANTENNA_c661_A0 (.DIODE(net1082));
 sky130_fd_sc_hd__diode_2 ANTENNA_c660_A3 (.DIODE(net1082));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_A2 (.DIODE(net1082));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout256_A (.DIODE(net1082));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout258_X (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_B1 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_A1 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c136_A3 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c760_A2 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_A1 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_S1 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_A1 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_S0 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_A2 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c235_A1 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout259_X (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_A2 (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_A2 (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_A0 (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c555_A3 (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c548_A1 (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_A2 (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_A1 (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c398_A0 (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_A3 (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c108_A1 (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_15_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_14_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_13_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_12_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_11_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_10_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_9_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_8_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_7_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_6_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_5_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_4_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_3_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_2_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_1_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_0_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_X (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge772_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge785_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge801_GATE_N (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge803_GATE_N (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge812_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s864_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s867_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s868_GATE_N (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s869_GATE_N (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_0_0_clk_X (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge820_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge833_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge845_GATE (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge847_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s866_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s880_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s883_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_1_0_clk_X (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge780_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge799_GATE_N (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge830_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s861_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s862_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s863_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s865_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s873_GATE_N (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_2_0_clk_X (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge770_CLK_N (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge792_GATE_N (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge813_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge824_CLK_N (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge856_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s875_SLEEP_B (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s877_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s878_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s879_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s881_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s893_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_3_0_clk_X (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge793_GATE (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge825_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge829_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge834_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge843_GATE_N (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge848_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge853_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s882_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s897_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s898_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_4_0_clk_X (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge781_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge838_GATE_N (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge840_GATE (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge849_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge854_CLK_N (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s895_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s923_SLEEP_B (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_6_0_clk_X (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge836_GATE_N (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge841_GATE_N (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge842_GATE_N (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge850_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s922_GATE (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s924_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_7_0_clk_X (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge777_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge795_GATE (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge806_GATE (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s860_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s871_GATE_N (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s872_GATE_N (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s874_GATE (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s876_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s888_GATE_N (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_8_0_clk_X (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge819_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge831_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge844_GATE (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge859_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s913_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s916_GATE_N (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s917_GATE_N (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s918_GATE (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s919_GATE_N (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s920_GATE_N (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s921_GATE_N (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s937_GATE_N (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_12_0_clk_X (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge805_GATE (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge823_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge839_GATE (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge851_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge855_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge857_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s932_GATE_N (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s935_GATE_N (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s936_GATE_N (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s938_GATE (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_13_0_clk_X (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c400_CLK_N (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge765_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s902_GATE (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s903_GATE_N (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s904_GATE_N (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s907_SLEEP_B (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s910_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s912_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s914_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s915_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s925_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_14_0_clk_X (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge766_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge784_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge811_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s926_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s927_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s928_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s929_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s930_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s931_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s933_GATE_N (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s934_GATE (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_15_0_clk_X (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_S1 (.DIODE(clknet_1_0__leaf_net692));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_S1 (.DIODE(clknet_1_0__leaf_net692));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_S0 (.DIODE(clknet_1_0__leaf_net692));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_S1 (.DIODE(clknet_1_0__leaf_net692));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net692_X (.DIODE(clknet_1_0__leaf_net692));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net673_A (.DIODE(clknet_0_net673));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net673_A (.DIODE(clknet_0_net673));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net673_X (.DIODE(clknet_0_net673));
 sky130_fd_sc_hd__diode_2 ANTENNA_c679_S0 (.DIODE(clknet_1_0__leaf_net673));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_S0 (.DIODE(clknet_1_0__leaf_net673));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_A3 (.DIODE(clknet_1_0__leaf_net673));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_S1 (.DIODE(clknet_1_0__leaf_net673));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_S1 (.DIODE(clknet_1_0__leaf_net673));
 sky130_fd_sc_hd__diode_2 ANTENNA_c762_S1 (.DIODE(clknet_1_0__leaf_net673));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net673_X (.DIODE(clknet_1_0__leaf_net673));
 sky130_fd_sc_hd__diode_2 ANTENNA_c537_SET_B (.DIODE(clknet_1_1__leaf_net673));
 sky130_fd_sc_hd__diode_2 ANTENNA_c538_S0 (.DIODE(clknet_1_1__leaf_net673));
 sky130_fd_sc_hd__diode_2 ANTENNA_c539_S1 (.DIODE(clknet_1_1__leaf_net673));
 sky130_fd_sc_hd__diode_2 ANTENNA_c543_S0 (.DIODE(clknet_1_1__leaf_net673));
 sky130_fd_sc_hd__diode_2 ANTENNA_c545_S1 (.DIODE(clknet_1_1__leaf_net673));
 sky130_fd_sc_hd__diode_2 ANTENNA_c670_S0 (.DIODE(clknet_1_1__leaf_net673));
 sky130_fd_sc_hd__diode_2 ANTENNA_c671_A3 (.DIODE(clknet_1_1__leaf_net673));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net673_X (.DIODE(clknet_1_1__leaf_net673));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_A1 (.DIODE(clknet_1_0__leaf_net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_A1 (.DIODE(clknet_1_0__leaf_net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_A0 (.DIODE(clknet_1_0__leaf_net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net315_X (.DIODE(clknet_1_0__leaf_net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_S1 (.DIODE(clknet_1_0__leaf_net652));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_S1 (.DIODE(clknet_1_0__leaf_net652));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_S1 (.DIODE(clknet_1_0__leaf_net652));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_S1 (.DIODE(clknet_1_0__leaf_net652));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_S0 (.DIODE(clknet_1_0__leaf_net652));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net652_X (.DIODE(clknet_1_0__leaf_net652));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_S1 (.DIODE(clknet_1_0__leaf_net651));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_S1 (.DIODE(clknet_1_0__leaf_net651));
 sky130_fd_sc_hd__diode_2 ANTENNA_c350_S1 (.DIODE(clknet_1_0__leaf_net651));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_S1 (.DIODE(clknet_1_0__leaf_net651));
 sky130_fd_sc_hd__diode_2 ANTENNA_c370_S1 (.DIODE(clknet_1_0__leaf_net651));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_S0 (.DIODE(clknet_1_0__leaf_net651));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net651_X (.DIODE(clknet_1_0__leaf_net651));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_S1 (.DIODE(clknet_1_1__leaf_net651));
 sky130_fd_sc_hd__diode_2 ANTENNA_c344_S1 (.DIODE(clknet_1_1__leaf_net651));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_S1 (.DIODE(clknet_1_1__leaf_net651));
 sky130_fd_sc_hd__diode_2 ANTENNA_c346_S1 (.DIODE(clknet_1_1__leaf_net651));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_S1 (.DIODE(clknet_1_1__leaf_net651));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_S1 (.DIODE(clknet_1_1__leaf_net651));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_S0 (.DIODE(clknet_1_1__leaf_net651));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net651_X (.DIODE(clknet_1_1__leaf_net651));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_A1 (.DIODE(clknet_1_1__leaf_net177));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_A2 (.DIODE(clknet_1_1__leaf_net177));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_A2 (.DIODE(clknet_1_1__leaf_net177));
 sky130_fd_sc_hd__diode_2 ANTENNA_c615_A2 (.DIODE(clknet_1_1__leaf_net177));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_A0 (.DIODE(clknet_1_1__leaf_net177));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net177_X (.DIODE(clknet_1_1__leaf_net177));
 sky130_fd_sc_hd__diode_2 ANTENNA_c350_A0 (.DIODE(clknet_1_1__leaf_net173));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_S0 (.DIODE(clknet_1_1__leaf_net173));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_A3 (.DIODE(clknet_1_1__leaf_net173));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_A2 (.DIODE(clknet_1_1__leaf_net173));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net173_X (.DIODE(clknet_1_1__leaf_net173));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_S0 (.DIODE(clknet_1_0__leaf_net155));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_A2 (.DIODE(clknet_1_0__leaf_net155));
 sky130_fd_sc_hd__diode_2 ANTENNA_c446_A1 (.DIODE(clknet_1_0__leaf_net155));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_A1 (.DIODE(clknet_1_0__leaf_net155));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_A2 (.DIODE(clknet_1_0__leaf_net155));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_A0 (.DIODE(clknet_1_0__leaf_net155));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net155_X (.DIODE(clknet_1_0__leaf_net155));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_A3 (.DIODE(clknet_1_1__leaf_net155));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_A3 (.DIODE(clknet_1_1__leaf_net155));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_A2 (.DIODE(clknet_1_1__leaf_net155));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_A0 (.DIODE(clknet_1_1__leaf_net155));
 sky130_fd_sc_hd__diode_2 ANTENNA_c742_A2 (.DIODE(clknet_1_1__leaf_net155));
 sky130_fd_sc_hd__diode_2 ANTENNA_c747_A2 (.DIODE(clknet_1_1__leaf_net155));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net155_X (.DIODE(clknet_1_1__leaf_net155));
 sky130_fd_sc_hd__diode_2 ANTENNA_c205_A0 (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer7_X (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA_c613_A1 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer9_A (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer8_X (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c190_A2 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_A1 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_A2 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_A1 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_B1 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone13_X (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer15_A (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c673_A3 (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer14_X (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_A2 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c234_A1 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_A2 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_S1 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_A3 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone17_X (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c660_A0 (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c757_A3 (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c761_A0 (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c531_A2 (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_S0 (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone18_X (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c669_A3 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c428_A3 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c613_A0 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c672_A2 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_A2 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone19_X (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_A3 (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_A1 (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer21_X (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer23_A (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_A3 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_A3 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer22_X (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c747_A0 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A2 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer25_A (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer24_X (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_A2 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer21_A (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_A0 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_A0 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_A1 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone28_X (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c582_A0 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c414_A1 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c183_A0 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_S1 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_A3 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone29_X (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_A3 (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_A2 (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_c366_A2 (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_A2 (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_A2 (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone31_X (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone31_A (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer32_X (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_A1 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_A3 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c611_A1 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c761_A1 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_S0 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone34_X (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer33_A (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_A1 (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c208_A2 (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_A3 (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone35_X (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_S0 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_A3 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c218_A0 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c228_A2 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_A3 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone36_X (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_A2 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_A3 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_A1 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_A2 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c229_A3 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone37_X (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_S1 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_S1 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone13_A1 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_A3 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_A3 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone38_X (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c720_A3 (.DIODE(net1038));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold58_X (.DIODE(net1038));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1_X (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_A1 (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_A3 (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_A3 (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_c148_A3 (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_A3 (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_B1 (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone13_A3 (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_A4 (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_A3 (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_S0 (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout2_X (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c136_A2 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_B1 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_S1 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_S1 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_A4 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_B1 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c138_A3 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_B1 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_A1 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_B1 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout4_X (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c431_RESET_B (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c399_A1 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_S0 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_A0 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c136_S1 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_A3 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_A0 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_S0 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_A1 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c103_A2 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout5_X (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_c549_A1 (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_c398_S0 (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_A0 (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_A2 (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_A1 (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_c264_A4 (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_c158_B1 (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_A3 (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_A3 (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_c124_A2 (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout6_X (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_c528_A2 (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone13_A4 (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_A4 (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_c530_S0 (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_c273_B1 (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_c269_A2 (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_c266_A2 (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_A3 (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_A3 (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_c136_A0 (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(net282));
 sky130_fd_sc_hd__mux4_1 clone1 (.A0(net106),
    .A1(net914),
    .A2(net111),
    .A3(net917),
    .S0(net964),
    .S1(net1054),
    .X(net1043));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer13 (.A(net874),
    .X(net1044));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer16 (.A(net1044),
    .X(net1045));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer17 (.A(net874),
    .X(net1046));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer18 (.A(net874),
    .X(net1047));
 sky130_fd_sc_hd__a41o_1 clone20 (.A1(net977),
    .A2(net974),
    .A3(net959),
    .A4(net967),
    .B1(net727),
    .X(net1048));
 sky130_fd_sc_hd__mux4_1 clone21 (.A0(net904),
    .A1(net59),
    .A2(net761),
    .A3(net56),
    .S0(net928),
    .S1(net881),
    .X(net1049));
 sky130_fd_sc_hd__mux4_1 clone22 (.A0(net1085),
    .A1(net15),
    .A2(net924),
    .A3(net1020),
    .S0(net1016),
    .S1(net908),
    .X(net1050));
 sky130_fd_sc_hd__a41o_1 clone23 (.A1(net1085),
    .A2(net15),
    .A3(net1020),
    .A4(net1042),
    .B1(net12),
    .X(net1051));
 sky130_fd_sc_hd__a41o_1 clone24 (.A1(net12),
    .A2(net924),
    .A3(net1020),
    .A4(net15),
    .B1(net1085),
    .X(net1052));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer28 (.A(net852),
    .X(net1053));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer29 (.A(net1053),
    .X(net1054));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer31 (.A(net1054),
    .X(net1055));
 sky130_fd_sc_hd__clkbuf_1 clone32 (.A(net18),
    .X(net1056));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer34 (.A(net416),
    .X(net1057));
 sky130_fd_sc_hd__clkbuf_1 clone39 (.A(net21),
    .X(net1058));
 sky130_fd_sc_hd__clkbuf_1 clone40 (.A(net822),
    .X(net1059));
 sky130_fd_sc_hd__clkbuf_1 clone41 (.A(net20),
    .X(net1060));
 sky130_fd_sc_hd__clkbuf_1 clone42 (.A(net13),
    .X(net1061));
 sky130_fd_sc_hd__clkbuf_1 clone43 (.A(net8),
    .X(net1062));
 sky130_fd_sc_hd__clkbuf_1 clone44 (.A(net22),
    .X(net1063));
 sky130_fd_sc_hd__clkbuf_1 clone45 (.A(net1065),
    .X(net1064));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer46 (.A(net31),
    .X(net1065));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer47 (.A(net35),
    .X(net1066));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer48 (.A(net1066),
    .X(net1067));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer49 (.A(net1067),
    .X(net1068));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer50 (.A(net1068),
    .X(net1069));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer51 (.A(net35),
    .X(net1070));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer52 (.A(net37),
    .X(net1071));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer53 (.A(net1071),
    .X(net1072));
 sky130_fd_sc_hd__clkbuf_1 rebuffer54 (.A(net1072),
    .X(net1073));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer55 (.A(net37),
    .X(net1074));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer56 (.A(net33),
    .X(net1075));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer57 (.A(net1075),
    .X(net1076));
 sky130_fd_sc_hd__clkbuf_1 clone58 (.A(net18),
    .X(net1077));
 sky130_fd_sc_hd__clkbuf_1 clone59 (.A(net978),
    .X(net1078));
 sky130_fd_sc_hd__clkbuf_1 clone60 (.A(net733),
    .X(net1079));
 sky130_fd_sc_hd__clkbuf_1 clone61 (.A(net767),
    .X(net1080));
 sky130_fd_sc_hd__clkbuf_1 clone62 (.A(net728),
    .X(net1081));
 sky130_fd_sc_hd__clkbuf_1 clone63 (.A(net732),
    .X(net1082));
 sky130_fd_sc_hd__clkbuf_1 clone64 (.A(net811),
    .X(net1083));
 sky130_fd_sc_hd__clkbuf_1 clone65 (.A(net6),
    .X(net1084));
 sky130_fd_sc_hd__clkbuf_1 clone66 (.A(net921),
    .X(net1085));
 sky130_fd_sc_hd__clkbuf_1 clone67 (.A(net922),
    .X(net1086));
 sky130_fd_sc_hd__decap_6 FILLER_0_0_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_79 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_303 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_115 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_20 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_267 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_198 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_104 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_280 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_115 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_64 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_508 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_140 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_423 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_435 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_31 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_227 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_507 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_511 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_128 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_368 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_86 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_245 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_367 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_387 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_438 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_351 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_435 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_527 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_560 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_198 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_525 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_471 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_455 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_452 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_74 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_104 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_339 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_88 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_471 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_525 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_506 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_115 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_415 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_497 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_543 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_308 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_525 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_431 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_442 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_384 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_103 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_448 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_479 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_487 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_507 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_5 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_131 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_219 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_135 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_242 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_462 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_395 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_219 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_275 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_5 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_523 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_5 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_490 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_617 ();
endmodule
