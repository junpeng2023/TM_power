module netlist_2 (clk,
    in0,
    in1,
    in10,
    in11,
    in12,
    in13,
    in14,
    in15,
    in16,
    in17,
    in18,
    in19,
    in2,
    in20,
    in21,
    in22,
    in23,
    in24,
    in25,
    in26,
    in27,
    in28,
    in29,
    in3,
    in30,
    in31,
    in32,
    in33,
    in34,
    in35,
    in36,
    in37,
    in38,
    in39,
    in4,
    in40,
    in41,
    in42,
    in43,
    in44,
    in45,
    in46,
    in47,
    in48,
    in49,
    in5,
    in50,
    in51,
    in52,
    in53,
    in54,
    in55,
    in56,
    in57,
    in58,
    in59,
    in6,
    in60,
    in61,
    in62,
    in63,
    in64,
    in65,
    in66,
    in67,
    in68,
    in69,
    in7,
    in70,
    in71,
    in72,
    in73,
    in74,
    in75,
    in76,
    in77,
    in78,
    in79,
    in8,
    in80,
    in81,
    in82,
    in83,
    in84,
    in85,
    in86,
    in87,
    in88,
    in89,
    in9,
    in90,
    in91,
    in92,
    in93,
    in94,
    in95,
    in96,
    in97,
    in98,
    in99,
    out0,
    out1,
    out10,
    out11,
    out12,
    out13,
    out14,
    out15,
    out16,
    out17,
    out18,
    out19,
    out2,
    out20,
    out21,
    out22,
    out23,
    out24,
    out25,
    out26,
    out27,
    out28,
    out29,
    out3,
    out30,
    out31,
    out32,
    out33,
    out34,
    out35,
    out36,
    out37,
    out38,
    out39,
    out4,
    out40,
    out41,
    out42,
    out43,
    out44,
    out45,
    out46,
    out47,
    out48,
    out49,
    out5,
    out50,
    out51,
    out52,
    out53,
    out54,
    out55,
    out56,
    out57,
    out58,
    out59,
    out6,
    out60,
    out61,
    out62,
    out63,
    out64,
    out65,
    out66,
    out67,
    out68,
    out69,
    out7,
    out70,
    out71,
    out72,
    out73,
    out74,
    out75,
    out76,
    out77,
    out78,
    out79,
    out8,
    out80,
    out81,
    out82,
    out83,
    out84,
    out85,
    out86,
    out87,
    out88,
    out89,
    out9,
    out90,
    out91,
    out92,
    out93,
    out94,
    out95,
    out96,
    out97,
    out98,
    out99,
    rst);
 input clk;
 input in0;
 input in1;
 input in10;
 input in11;
 input in12;
 input in13;
 input in14;
 input in15;
 input in16;
 input in17;
 input in18;
 input in19;
 input in2;
 input in20;
 input in21;
 input in22;
 input in23;
 input in24;
 input in25;
 input in26;
 input in27;
 input in28;
 input in29;
 input in3;
 input in30;
 input in31;
 input in32;
 input in33;
 input in34;
 input in35;
 input in36;
 input in37;
 input in38;
 input in39;
 input in4;
 input in40;
 input in41;
 input in42;
 input in43;
 input in44;
 input in45;
 input in46;
 input in47;
 input in48;
 input in49;
 input in5;
 input in50;
 input in51;
 input in52;
 input in53;
 input in54;
 input in55;
 input in56;
 input in57;
 input in58;
 input in59;
 input in6;
 input in60;
 input in61;
 input in62;
 input in63;
 input in64;
 input in65;
 input in66;
 input in67;
 input in68;
 input in69;
 input in7;
 input in70;
 input in71;
 input in72;
 input in73;
 input in74;
 input in75;
 input in76;
 input in77;
 input in78;
 input in79;
 input in8;
 input in80;
 input in81;
 input in82;
 input in83;
 input in84;
 input in85;
 input in86;
 input in87;
 input in88;
 input in89;
 input in9;
 input in90;
 input in91;
 input in92;
 input in93;
 input in94;
 input in95;
 input in96;
 input in97;
 input in98;
 input in99;
 output out0;
 output out1;
 output out10;
 output out11;
 output out12;
 output out13;
 output out14;
 output out15;
 output out16;
 output out17;
 output out18;
 output out19;
 output out2;
 output out20;
 output out21;
 output out22;
 output out23;
 output out24;
 output out25;
 output out26;
 output out27;
 output out28;
 output out29;
 output out3;
 output out30;
 output out31;
 output out32;
 output out33;
 output out34;
 output out35;
 output out36;
 output out37;
 output out38;
 output out39;
 output out4;
 output out40;
 output out41;
 output out42;
 output out43;
 output out44;
 output out45;
 output out46;
 output out47;
 output out48;
 output out49;
 output out5;
 output out50;
 output out51;
 output out52;
 output out53;
 output out54;
 output out55;
 output out56;
 output out57;
 output out58;
 output out59;
 output out6;
 output out60;
 output out61;
 output out62;
 output out63;
 output out64;
 output out65;
 output out66;
 output out67;
 output out68;
 output out69;
 output out7;
 output out70;
 output out71;
 output out72;
 output out73;
 output out74;
 output out75;
 output out76;
 output out77;
 output out78;
 output out79;
 output out8;
 output out80;
 output out81;
 output out82;
 output out83;
 output out84;
 output out85;
 output out86;
 output out87;
 output out88;
 output out89;
 output out9;
 output out90;
 output out91;
 output out92;
 output out93;
 output out94;
 output out95;
 output out96;
 output out97;
 output out98;
 output out99;
 input rst;

 wire net0;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net63;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net64;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net65;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net66;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net67;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net68;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net69;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net7;
 wire net70;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net144;
 wire net557;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_0_net698;
 wire clknet_1_0__leaf_net698;
 wire clknet_1_1__leaf_net698;
 wire clknet_0_net697;
 wire clknet_1_0__leaf_net697;
 wire clknet_1_1__leaf_net697;
 wire clknet_0_net696;
 wire clknet_1_0__leaf_net696;
 wire clknet_1_1__leaf_net696;
 wire clknet_0_net521;
 wire clknet_1_0__leaf_net521;
 wire clknet_1_1__leaf_net521;
 wire clknet_0_net522;
 wire clknet_1_0__leaf_net522;
 wire clknet_1_1__leaf_net522;
 wire clknet_0_net526;
 wire clknet_1_0__leaf_net526;
 wire clknet_1_1__leaf_net526;
 wire clknet_0_net502;
 wire clknet_1_0__leaf_net502;
 wire clknet_1_1__leaf_net502;
 wire clknet_0_net677;
 wire clknet_1_0__leaf_net677;
 wire clknet_1_1__leaf_net677;
 wire clknet_0_net463;
 wire clknet_1_0__leaf_net463;
 wire clknet_1_1__leaf_net463;
 wire clknet_0_net482;
 wire clknet_1_0__leaf_net482;
 wire clknet_1_1__leaf_net482;
 wire clknet_0_net488;
 wire clknet_1_0__leaf_net488;
 wire clknet_1_1__leaf_net488;
 wire clknet_0_net676;
 wire clknet_1_0__leaf_net676;
 wire clknet_1_1__leaf_net676;
 wire clknet_0_net459;
 wire clknet_1_0__leaf_net459;
 wire clknet_1_1__leaf_net459;
 wire clknet_0_net466;
 wire clknet_1_0__leaf_net466;
 wire clknet_1_1__leaf_net466;
 wire clknet_0_net473;
 wire clknet_1_0__leaf_net473;
 wire clknet_1_1__leaf_net473;
 wire clknet_0_net675;
 wire clknet_1_0__leaf_net675;
 wire clknet_1_1__leaf_net675;
 wire clknet_0_net656;
 wire clknet_1_0__leaf_net656;
 wire clknet_1_1__leaf_net656;
 wire clknet_0_net314;
 wire clknet_1_0__leaf_net314;
 wire clknet_1_1__leaf_net314;
 wire clknet_0_net655;
 wire clknet_1_0__leaf_net655;
 wire clknet_1_1__leaf_net655;
 wire clknet_0_net420;
 wire clknet_1_0__leaf_net420;
 wire clknet_1_1__leaf_net420;
 wire clknet_0_net412;
 wire clknet_1_0__leaf_net412;
 wire clknet_1_1__leaf_net412;
 wire clknet_0_net809;
 wire clknet_1_0__leaf_net809;
 wire clknet_1_1__leaf_net809;
 wire clknet_0_net855;
 wire clknet_1_0__leaf_net855;
 wire clknet_1_1__leaf_net855;
 wire clknet_0_net317;
 wire clknet_1_0__leaf_net317;
 wire clknet_1_1__leaf_net317;
 wire clknet_0_net318;
 wire clknet_1_0__leaf_net318;
 wire clknet_1_1__leaf_net318;
 wire clknet_0_net654;
 wire clknet_1_0__leaf_net654;
 wire clknet_1_1__leaf_net654;
 wire clknet_0_net821;
 wire clknet_1_0__leaf_net821;
 wire clknet_1_1__leaf_net821;
 wire clknet_0_net638;
 wire clknet_1_0__leaf_net638;
 wire clknet_1_1__leaf_net638;
 wire clknet_0_net207;
 wire clknet_1_0__leaf_net207;
 wire clknet_1_1__leaf_net207;
 wire clknet_0_net824;
 wire clknet_1_0__leaf_net824;
 wire clknet_1_1__leaf_net824;
 wire clknet_0_net204;
 wire clknet_1_0__leaf_net204;
 wire clknet_1_1__leaf_net204;
 wire clknet_0_net816;
 wire clknet_1_0__leaf_net816;
 wire clknet_1_1__leaf_net816;
 wire clknet_0_net812;
 wire clknet_1_0__leaf_net812;
 wire clknet_1_1__leaf_net812;
 wire clknet_0_net637;
 wire clknet_1_0__leaf_net637;
 wire clknet_1_1__leaf_net637;
 wire clknet_0_net289;
 wire clknet_1_0__leaf_net289;
 wire clknet_1_1__leaf_net289;
 wire clknet_0_net285;
 wire clknet_1_0__leaf_net285;
 wire clknet_1_1__leaf_net285;
 wire clknet_0_net401;
 wire clknet_1_0__leaf_net401;
 wire clknet_1_1__leaf_net401;
 wire clknet_0_net504;
 wire clknet_1_0__leaf_net504;
 wire clknet_1_1__leaf_net504;
 wire clknet_0_net511;
 wire clknet_1_0__leaf_net511;
 wire clknet_1_1__leaf_net511;
 wire clknet_0_net396;
 wire clknet_1_0__leaf_net396;
 wire clknet_1_1__leaf_net396;
 wire clknet_0_net605;
 wire clknet_1_0__leaf_net605;
 wire clknet_1_1__leaf_net605;
 wire clknet_0_net398;
 wire clknet_1_0__leaf_net398;
 wire clknet_1_1__leaf_net398;
 wire clknet_0_net380;
 wire clknet_1_0__leaf_net380;
 wire clknet_1_1__leaf_net380;
 wire clknet_0_net392;
 wire clknet_1_0__leaf_net392;
 wire clknet_1_1__leaf_net392;
 wire clknet_0_net282;
 wire clknet_1_0__leaf_net282;
 wire clknet_1_1__leaf_net282;
 wire clknet_0_net286;
 wire clknet_1_0__leaf_net286;
 wire clknet_1_1__leaf_net286;
 wire clknet_0_net290;
 wire clknet_1_0__leaf_net290;
 wire clknet_1_1__leaf_net290;
 wire clknet_0_net291;
 wire clknet_1_0__leaf_net291;
 wire clknet_1_1__leaf_net291;
 wire clknet_0_net852;
 wire clknet_1_0__leaf_net852;
 wire clknet_1_1__leaf_net852;
 wire clknet_0_net841;
 wire clknet_1_0__leaf_net841;
 wire clknet_1_1__leaf_net841;
 wire clknet_0_net191;
 wire clknet_1_0__leaf_net191;
 wire clknet_1_1__leaf_net191;
 wire clknet_0_net604;
 wire clknet_1_0__leaf_net604;
 wire clknet_1_1__leaf_net604;
 wire clknet_0_net838;
 wire clknet_1_0__leaf_net838;
 wire clknet_1_1__leaf_net838;
 wire clknet_0_net862;
 wire clknet_1_0__leaf_net862;
 wire clknet_1_1__leaf_net862;
 wire clknet_0_net94;
 wire clknet_1_0__leaf_net94;
 wire clknet_1_1__leaf_net94;
 wire clknet_0_net836;
 wire clknet_1_0__leaf_net836;
 wire clknet_1_1__leaf_net836;
 wire clknet_0_net75;
 wire clknet_1_0__leaf_net75;
 wire clknet_1_1__leaf_net75;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net942;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;

 sky130_fd_sc_hd__a41o_1 c100 (.A1(net793),
    .A2(net796),
    .A3(net751),
    .A4(net740),
    .B1(net794),
    .X(net0));
 sky130_fd_sc_hd__a41o_1 c101 (.A1(net775),
    .A2(net767),
    .A3(net793),
    .A4(net0),
    .B1(net782),
    .X(net1));
 sky130_fd_sc_hd__a31o_1 c102 (.A1(net794),
    .A2(net1),
    .A3(net721),
    .B1(net801),
    .X(net873));
 sky130_fd_sc_hd__mux4_2 c103 (.A0(net799),
    .A1(net782),
    .A2(net1),
    .A3(net719),
    .S0(net797),
    .S1(net776),
    .X(net869));
 sky130_fd_sc_hd__a31o_1 c104 (.A1(net756),
    .A2(net797),
    .A3(net744),
    .B1(net773),
    .X(net2));
 sky130_fd_sc_hd__a41o_1 c105 (.A1(net802),
    .A2(net797),
    .A3(net2),
    .A4(net869),
    .B1(net791),
    .X(net3));
 sky130_fd_sc_hd__a41o_1 c106 (.A1(net2),
    .A2(net3),
    .A3(net795),
    .A4(net797),
    .B1(net796),
    .X(net864));
 sky130_fd_sc_hd__mux4_1 c107 (.A0(net1),
    .A1(net796),
    .A2(net3),
    .A3(net786),
    .S0(net744),
    .S1(net873),
    .X(net4));
 sky130_fd_sc_hd__mux4_2 c108 (.A0(net4),
    .A1(net723),
    .A2(net790),
    .A3(net740),
    .S0(net751),
    .S1(net3),
    .X(net5));
 sky130_fd_sc_hd__mux4_1 c109 (.A0(net799),
    .A1(net2),
    .A2(net801),
    .A3(net864),
    .S0(net4),
    .S1(net1),
    .X(net857));
 sky130_fd_sc_hd__a31o_4 c122 (.A1(net3),
    .A2(net789),
    .A3(net796),
    .B1(net791),
    .X(net860));
 sky130_fd_sc_hd__mux4_2 c123 (.A0(net751),
    .A1(net780),
    .A2(net796),
    .A3(net860),
    .S0(net765),
    .S1(net791),
    .X(net6));
 sky130_fd_sc_hd__a41o_1 c124 (.A1(net766),
    .A2(net6),
    .A3(net860),
    .A4(net797),
    .B1(net801),
    .X(net7));
 sky130_fd_sc_hd__a41o_1 c125 (.A1(net791),
    .A2(net860),
    .A3(net6),
    .A4(net765),
    .B1(net908),
    .X(net858));
 sky130_fd_sc_hd__a41o_1 c126 (.A1(net0),
    .A2(net860),
    .A3(net858),
    .A4(net7),
    .B1(net6),
    .X(net875));
 sky130_fd_sc_hd__mux4_2 c127 (.A0(net740),
    .A1(net751),
    .A2(net776),
    .A3(net797),
    .S0(net860),
    .S1(net858),
    .X(net865));
 sky130_fd_sc_hd__mux4_2 c128 (.A0(net6),
    .A1(net875),
    .A2(net865),
    .A3(net858),
    .S0(net908),
    .S1(net860),
    .X(net872));
 sky130_fd_sc_hd__mux4_1 c129 (.A0(net7),
    .A1(net858),
    .A2(net865),
    .A3(net875),
    .S0(net860),
    .S1(net872),
    .X(net874));
 sky130_fd_sc_hd__mux4_1 c130 (.A0(net765),
    .A1(net6),
    .A2(net872),
    .A3(net865),
    .S0(net779),
    .S1(net874),
    .X(net842));
 sky130_fd_sc_hd__mux4_1 c131 (.A0(net753),
    .A1(net875),
    .A2(net842),
    .A3(net860),
    .S0(net872),
    .S1(net858),
    .X(net870));
 sky130_fd_sc_hd__xnor2_4 c132 (.A(net760),
    .B(net708),
    .Y(net8));
 sky130_fd_sc_hd__a21bo_1 c133 (.A1(net770),
    .A2(net739),
    .B1_N(net905),
    .X(net9));
 sky130_fd_sc_hd__a21bo_4 c134 (.A1(net144),
    .A2(net707),
    .B1_N(net750),
    .X(net10));
 sky130_fd_sc_hd__xnor2_4 c135 (.A(net712),
    .B(net10),
    .Y(net11));
 sky130_fd_sc_hd__a21bo_2 c136 (.A1(net781),
    .A2(net11),
    .B1_N(net760),
    .X(net12));
 sky130_fd_sc_hd__mux4_2 c137 (.A0(net12),
    .A1(net781),
    .A2(net10),
    .A3(net714),
    .S0(net715),
    .S1(net905),
    .X(net13));
 sky130_fd_sc_hd__xnor2_1 c138 (.A(net11),
    .B(net792),
    .Y(net14));
 sky130_fd_sc_hd__xnor2_4 c139 (.A(net8),
    .B(net750),
    .Y(net15));
 sky130_fd_sc_hd__xnor2_2 c140 (.A(net718),
    .B(net719),
    .Y(net16));
 sky130_fd_sc_hd__a41o_4 c141 (.A1(net9),
    .A2(net8),
    .A3(net14),
    .A4(net717),
    .B1(net12),
    .X(net17));
 sky130_fd_sc_hd__xnor2_1 c142 (.A(net10),
    .B(net709),
    .Y(net18));
 sky130_fd_sc_hd__xnor2_4 c143 (.A(net717),
    .B(net15),
    .Y(net19));
 sky130_fd_sc_hd__a41o_2 c144 (.A1(net714),
    .A2(net19),
    .A3(net9),
    .A4(net715),
    .B1(net716),
    .X(net20));
 sky130_fd_sc_hd__a21bo_4 c145 (.A1(net14),
    .A2(net13),
    .B1_N(net11),
    .X(net21));
 sky130_fd_sc_hd__a41o_2 c146 (.A1(net17),
    .A2(net11),
    .A3(net770),
    .A4(net715),
    .B1(net905),
    .X(net22));
 sky130_fd_sc_hd__xnor2_2 c147 (.A(net16),
    .B(net19),
    .Y(net23));
 sky130_fd_sc_hd__a21bo_4 c148 (.A1(net11),
    .A2(net16),
    .B1_N(net718),
    .X(net24));
 sky130_fd_sc_hd__a21bo_4 c149 (.A1(net24),
    .A2(net710),
    .B1_N(net11),
    .X(net871));
 sky130_fd_sc_hd__a21bo_1 c150 (.A1(net12),
    .A2(net21),
    .B1_N(net905),
    .X(net25));
 sky130_fd_sc_hd__a41o_1 c151 (.A1(net24),
    .A2(net770),
    .A3(net557),
    .A4(net17),
    .B1(net18),
    .X(net26));
 sky130_fd_sc_hd__mux4_2 c152 (.A0(net15),
    .A1(net750),
    .A2(net18),
    .A3(net19),
    .S0(net892),
    .S1(net24),
    .X(net27));
 sky130_fd_sc_hd__a21bo_4 c153 (.A1(net26),
    .A2(net27),
    .B1_N(net916),
    .X(net28));
 sky130_fd_sc_hd__a21bo_1 c154 (.A1(net707),
    .A2(net731),
    .B1_N(net715),
    .X(net29));
 sky130_fd_sc_hd__a31o_1 c155 (.A1(net712),
    .A2(net709),
    .A3(net750),
    .B1(net905),
    .X(net30));
 sky130_fd_sc_hd__a21bo_4 c156 (.A1(net743),
    .A2(net731),
    .B1_N(net725),
    .X(net863));
 sky130_fd_sc_hd__a21bo_4 c157 (.A1(net30),
    .A2(net707),
    .B1_N(net901),
    .X(net31));
 sky130_fd_sc_hd__a31o_4 c158 (.A1(net750),
    .A2(net792),
    .A3(net31),
    .B1(net901),
    .X(net32));
 sky130_fd_sc_hd__a21bo_1 c159 (.A1(net734),
    .A2(net30),
    .B1_N(net732),
    .X(net33));
 sky130_fd_sc_hd__a41o_4 c160 (.A1(net31),
    .A2(net742),
    .A3(net735),
    .A4(net32),
    .B1(net901),
    .X(net34));
 sky130_fd_sc_hd__a31o_4 c161 (.A1(net732),
    .A2(net27),
    .A3(net34),
    .B1(net901),
    .X(net35));
 sky130_fd_sc_hd__a41o_4 c162 (.A1(net737),
    .A2(net34),
    .A3(net724),
    .A4(net35),
    .B1(net901),
    .X(net808));
 sky130_fd_sc_hd__mux4_1 c163 (.A0(net31),
    .A1(net729),
    .A2(net35),
    .A3(net723),
    .S0(net34),
    .S1(net901),
    .X(net36));
 sky130_fd_sc_hd__a31o_4 c164 (.A1(net719),
    .A2(net35),
    .A3(net32),
    .B1(net901),
    .X(net37));
 sky130_fd_sc_hd__mux4_1 c165 (.A0(net731),
    .A1(net32),
    .A2(net33),
    .A3(net36),
    .S0(net908),
    .S1(net939),
    .X(net38));
 sky130_fd_sc_hd__a21bo_4 c166 (.A1(net33),
    .A2(net725),
    .B1_N(net34),
    .X(net39));
 sky130_fd_sc_hd__a41o_1 c167 (.A1(net808),
    .A2(net722),
    .A3(net727),
    .A4(net901),
    .B1(net39),
    .X(net40));
 sky130_fd_sc_hd__mux4_2 c168 (.A0(net18),
    .A1(net37),
    .A2(net735),
    .A3(net738),
    .S0(net720),
    .S1(net901),
    .X(net41));
 sky130_fd_sc_hd__a21bo_1 c169 (.A1(net715),
    .A2(net740),
    .B1_N(net926),
    .X(net42));
 sky130_fd_sc_hd__mux4_2 c170 (.A0(net735),
    .A1(net738),
    .A2(net36),
    .A3(net41),
    .S0(net35),
    .S1(net10),
    .X(net43));
 sky130_fd_sc_hd__mux4_2 c171 (.A0(net36),
    .A1(net908),
    .A2(net39),
    .A3(net43),
    .S0(net41),
    .S1(net40),
    .X(net44));
 sky130_fd_sc_hd__mux4_2 c172 (.A0(net43),
    .A1(net927),
    .A2(net40),
    .A3(net42),
    .S0(net887),
    .S1(net743),
    .X(net45));
 sky130_fd_sc_hd__mux4_2 c173 (.A0(net35),
    .A1(net42),
    .A2(net45),
    .A3(net33),
    .S0(net808),
    .S1(net887),
    .X(net46));
 sky130_fd_sc_hd__mux4_2 c174 (.A0(net42),
    .A1(net46),
    .A2(net27),
    .A3(net713),
    .S0(net34),
    .S1(net887),
    .X(net47));
 sky130_fd_sc_hd__mux4_2 c175 (.A0(net40),
    .A1(net887),
    .A2(net735),
    .A3(net45),
    .S0(net723),
    .S1(net46),
    .X(net48));
 sky130_fd_sc_hd__a21bo_1 c176 (.A1(net30),
    .A2(net738),
    .B1_N(net759),
    .X(net49));
 sky130_fd_sc_hd__a31o_2 c177 (.A1(net720),
    .A2(net726),
    .A3(net749),
    .B1(net756),
    .X(net50));
 sky130_fd_sc_hd__a41o_1 c178 (.A1(net727),
    .A2(net762),
    .A3(net755),
    .A4(net941),
    .B1(net898),
    .X(net51));
 sky130_fd_sc_hd__a41o_1 c179 (.A1(net755),
    .A2(net725),
    .A3(net38),
    .A4(net898),
    .B1(net39),
    .X(net52));
 sky130_fd_sc_hd__a21bo_1 c180 (.A1(net709),
    .A2(net744),
    .B1_N(net898),
    .X(net53));
 sky130_fd_sc_hd__a21bo_1 c181 (.A1(net754),
    .A2(net888),
    .B1_N(net745),
    .X(net847));
 sky130_fd_sc_hd__a21bo_1 c182 (.A1(net708),
    .A2(net29),
    .B1_N(net892),
    .X(net54));
 sky130_fd_sc_hd__a21bo_1 c183 (.A1(net729),
    .A2(net748),
    .B1_N(net885),
    .X(net55));
 sky130_fd_sc_hd__mux4_2 c184 (.A0(net723),
    .A1(net733),
    .A2(net908),
    .A3(net885),
    .S0(net888),
    .S1(net898),
    .X(net56));
 sky130_fd_sc_hd__a31o_1 c185 (.A1(net733),
    .A2(net885),
    .A3(net888),
    .B1(net898),
    .X(net57));
 sky130_fd_sc_hd__a31o_1 c186 (.A1(net757),
    .A2(net723),
    .A3(net57),
    .B1(net898),
    .X(net861));
 sky130_fd_sc_hd__a21bo_1 c187 (.A1(net29),
    .A2(net708),
    .B1_N(net55),
    .X(net58));
 sky130_fd_sc_hd__a21bo_1 c188 (.A1(net49),
    .A2(net902),
    .B1_N(net57),
    .X(net59));
 sky130_fd_sc_hd__mux4_2 c189 (.A0(net45),
    .A1(net761),
    .A2(net54),
    .A3(net861),
    .S0(net941),
    .S1(net898),
    .X(net60));
 sky130_fd_sc_hd__a31o_1 c190 (.A1(net10),
    .A2(net888),
    .A3(net754),
    .B1(net898),
    .X(net61));
 sky130_fd_sc_hd__a21bo_1 c191 (.A1(net53),
    .A2(net861),
    .B1_N(net888),
    .X(net62));
 sky130_fd_sc_hd__mux4_2 c192 (.A0(net61),
    .A1(net56),
    .A2(net51),
    .A3(net60),
    .S0(net758),
    .S1(net54),
    .X(net63));
 sky130_fd_sc_hd__mux4_1 c193 (.A0(net38),
    .A1(net59),
    .A2(net53),
    .A3(net10),
    .S0(net941),
    .S1(net898),
    .X(net64));
 sky130_fd_sc_hd__mux4_1 c194 (.A0(net54),
    .A1(net62),
    .A2(net63),
    .A3(net29),
    .S0(net756),
    .S1(net61),
    .X(net65));
 sky130_fd_sc_hd__mux4_1 c195 (.A0(net62),
    .A1(net64),
    .A2(net63),
    .A3(net60),
    .S0(net898),
    .S1(net896),
    .X(net66));
 sky130_fd_sc_hd__a41o_2 c196 (.A1(net759),
    .A2(net60),
    .A3(net885),
    .A4(net29),
    .B1(net896),
    .X(net67));
 sky130_fd_sc_hd__mux4_1 c197 (.A0(net748),
    .A1(net64),
    .A2(net746),
    .A3(net38),
    .S0(net62),
    .S1(net67),
    .X(net68));
 sky130_fd_sc_hd__a21bo_2 c198 (.A1(net774),
    .A2(net782),
    .B1_N(net19),
    .X(net837));
 sky130_fd_sc_hd__a21bo_1 c199 (.A1(net39),
    .A2(net19),
    .B1_N(net761),
    .X(net69));
 sky130_fd_sc_hd__a21bo_1 c200 (.A1(net761),
    .A2(net786),
    .B1_N(net740),
    .X(net70));
 sky130_fd_sc_hd__a21bo_4 c201 (.A1(net59),
    .A2(net70),
    .B1_N(net773),
    .X(net849));
 sky130_fd_sc_hd__a21bo_1 c202 (.A1(net57),
    .A2(net849),
    .B1_N(net896),
    .X(net71));
 sky130_fd_sc_hd__a31o_1 c203 (.A1(net725),
    .A2(net837),
    .A3(net773),
    .B1(net849),
    .X(net72));
 sky130_fd_sc_hd__a41o_1 c204 (.A1(net70),
    .A2(net69),
    .A3(net769),
    .A4(net13),
    .B1(net774),
    .X(net73));
 sky130_fd_sc_hd__a31o_1 c205 (.A1(net72),
    .A2(net63),
    .A3(net849),
    .B1(net787),
    .X(net74));
 sky130_fd_sc_hd__a41o_1 c206 (.A1(net69),
    .A2(net784),
    .A3(net849),
    .A4(net763),
    .B1(clknet_1_0__leaf_net604),
    .X(net75));
 sky130_fd_sc_hd__buf_1 c207 (.A(net859),
    .X(net853));
 sky130_fd_sc_hd__clkbuf_4 c208 (.A(net859),
    .X(net868));
 sky130_fd_sc_hd__a21bo_1 c209 (.A1(net769),
    .A2(net885),
    .B1_N(net787),
    .X(net76));
 sky130_fd_sc_hd__a21bo_1 c210 (.A1(net749),
    .A2(net853),
    .B1_N(net849),
    .X(net77));
 sky130_fd_sc_hd__a21bo_1 c211 (.A1(net19),
    .A2(net76),
    .B1_N(net725),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_1 c212 (.A(net630),
    .X(net79));
 sky130_fd_sc_hd__a21bo_1 c213 (.A1(net777),
    .A2(net78),
    .B1_N(net896),
    .X(net80));
 sky130_fd_sc_hd__buf_1 c214 (.A(net851),
    .X(net81));
 sky130_fd_sc_hd__mux4_1 c215 (.A0(net48),
    .A1(net849),
    .A2(net79),
    .A3(net784),
    .S0(net78),
    .S1(net77),
    .X(net82));
 sky130_fd_sc_hd__mux4_1 c216 (.A0(net81),
    .A1(net767),
    .A2(net80),
    .A3(net70),
    .S0(net71),
    .S1(net948),
    .X(net83));
 sky130_fd_sc_hd__mux4_1 c217 (.A0(net78),
    .A1(net853),
    .A2(net868),
    .A3(net81),
    .S0(net606),
    .S1(net632),
    .X(net84));
 sky130_fd_sc_hd__mux4_1 c218 (.A0(net79),
    .A1(clknet_1_0__leaf_net75),
    .A2(net81),
    .A3(net78),
    .S0(net606),
    .S1(net856),
    .X(net85));
 sky130_fd_sc_hd__a31o_1 c219 (.A1(net84),
    .A2(net81),
    .A3(net606),
    .B1(net632),
    .X(net86));
 sky130_fd_sc_hd__clkbuf_2 c220 (.A(net851),
    .X(net87));
 sky130_fd_sc_hd__a21bo_1 c221 (.A1(net800),
    .A2(net87),
    .B1_N(net778),
    .X(net88));
 sky130_fd_sc_hd__a41o_1 c222 (.A1(clknet_1_1__leaf_net75),
    .A2(net87),
    .A3(net853),
    .A4(net837),
    .B1(net896),
    .X(net89));
 sky130_fd_sc_hd__a31o_2 c223 (.A1(net87),
    .A2(net885),
    .A3(net598),
    .B1(net606),
    .X(net867));
 sky130_fd_sc_hd__a41o_1 c224 (.A1(net88),
    .A2(net789),
    .A3(net867),
    .A4(net756),
    .B1(net51),
    .X(net90));
 sky130_fd_sc_hd__a21bo_1 c225 (.A1(net798),
    .A2(net726),
    .B1_N(net849),
    .X(net91));
 sky130_fd_sc_hd__a41o_2 c226 (.A1(net90),
    .A2(net802),
    .A3(net785),
    .A4(net758),
    .B1(net897),
    .X(net92));
 sky130_fd_sc_hd__a21bo_1 c227 (.A1(net73),
    .A2(net763),
    .B1_N(net859),
    .X(net866));
 sky130_fd_sc_hd__a31o_1 c228 (.A1(net91),
    .A2(net867),
    .A3(net808),
    .B1(net632),
    .X(net93));
 sky130_fd_sc_hd__a41o_1 c229 (.A1(net787),
    .A2(net802),
    .A3(net87),
    .A4(net798),
    .B1(clknet_1_1__leaf_net604),
    .X(net862));
 sky130_fd_sc_hd__a21bo_1 c230 (.A1(clknet_1_0__leaf_net862),
    .A2(net90),
    .B1_N(net866),
    .X(net94));
 sky130_fd_sc_hd__a21bo_1 c231 (.A1(net772),
    .A2(clknet_1_0__leaf_net94),
    .B1_N(net866),
    .X(net836));
 sky130_fd_sc_hd__mux4_1 c232 (.A0(net767),
    .A1(net90),
    .A2(net802),
    .A3(net92),
    .S0(clknet_1_0__leaf_net836),
    .S1(clknet_1_1__leaf_net604),
    .X(net95));
 sky130_fd_sc_hd__sdfbbn_1 c233 (.CLK_N(clknet_4_15_0_clk),
    .D(net51),
    .RESET_B(net0),
    .SCD(clknet_1_0__leaf_net836),
    .SCE(net857),
    .SET_B(net897),
    .Q(net835),
    .Q_N(net96));
 sky130_fd_sc_hd__buf_1 c234 (.A(net851),
    .X(net97));
 sky130_fd_sc_hd__dlymetal6s2s_1 c235 (.A(net851),
    .X(net846));
 sky130_fd_sc_hd__a21bo_1 c236 (.A1(net97),
    .A2(net866),
    .B1_N(net851),
    .X(net98));
 sky130_fd_sc_hd__mux4_1 c237 (.A0(net98),
    .A1(clknet_1_1__leaf_net94),
    .A2(clknet_1_1__leaf_net862),
    .A3(net800),
    .S0(clknet_1_1__leaf_net836),
    .S1(net96),
    .X(net99));
 sky130_fd_sc_hd__a21bo_1 c238 (.A1(net0),
    .A2(clknet_1_1__leaf_net604),
    .B1_N(net859),
    .X(net838));
 sky130_fd_sc_hd__a21bo_1 c239 (.A1(net92),
    .A2(net96),
    .B1_N(net897),
    .X(net854));
 sky130_fd_sc_hd__a41o_1 c240 (.A1(net854),
    .A2(clknet_1_0__leaf_net838),
    .A3(clknet_1_0__leaf_net836),
    .A4(net837),
    .B1(net851),
    .X(net100));
 sky130_fd_sc_hd__sdfbbn_2 c241 (.CLK_N(clknet_4_15_0_clk),
    .D(net796),
    .RESET_B(clknet_1_0__leaf_net94),
    .SCD(net854),
    .SCE(net846),
    .SET_B(net598),
    .Q(net834),
    .Q_N(net101));
 sky130_fd_sc_hd__xnor2_4 c264 (.A(net20),
    .B(net963),
    .Y(net102));
 sky130_fd_sc_hd__xnor2_4 c265 (.A(net715),
    .B(net21),
    .Y(net103));
 sky130_fd_sc_hd__a21bo_4 c266 (.A1(net102),
    .A2(net103),
    .B1_N(net905),
    .X(net104));
 sky130_fd_sc_hd__a21bo_1 c267 (.A1(net739),
    .A2(net22),
    .B1_N(net728),
    .X(net105));
 sky130_fd_sc_hd__xnor2_4 c268 (.A(net104),
    .B(net792),
    .Y(net106));
 sky130_fd_sc_hd__xnor2_1 c269 (.A(net716),
    .B(net104),
    .Y(net107));
 sky130_fd_sc_hd__xnor2_4 c270 (.A(net23),
    .B(net106),
    .Y(net108));
 sky130_fd_sc_hd__xnor2_2 c271 (.A(net108),
    .B(net106),
    .Y(net109));
 sky130_fd_sc_hd__a21bo_1 c272 (.A1(net109),
    .A2(net102),
    .B1_N(net108),
    .X(net110));
 sky130_fd_sc_hd__a41o_1 c273 (.A1(net105),
    .A2(net21),
    .A3(net792),
    .A4(net890),
    .B1(net22),
    .X(net111));
 sky130_fd_sc_hd__a21bo_4 c274 (.A1(net750),
    .A2(net106),
    .B1_N(net905),
    .X(net112));
 sky130_fd_sc_hd__a21bo_1 c275 (.A1(net111),
    .A2(net707),
    .B1_N(net105),
    .X(net113));
 sky130_fd_sc_hd__xnor2_2 c276 (.A(net113),
    .B(net12),
    .Y(net114));
 sky130_fd_sc_hd__xnor2_4 c277 (.A(net112),
    .B(net17),
    .Y(net115));
 sky130_fd_sc_hd__xnor2_4 c278 (.A(net890),
    .B(net115),
    .Y(net116));
 sky130_fd_sc_hd__a21bo_1 c279 (.A1(net111),
    .A2(net115),
    .B1_N(net905),
    .X(net117));
 sky130_fd_sc_hd__a41o_1 c280 (.A1(net117),
    .A2(net884),
    .A3(net15),
    .A4(net557),
    .B1(net108),
    .X(net118));
 sky130_fd_sc_hd__a41o_1 c281 (.A1(net114),
    .A2(net118),
    .A3(net112),
    .A4(net884),
    .B1(net104),
    .X(net119));
 sky130_fd_sc_hd__a41o_1 c282 (.A1(net119),
    .A2(net118),
    .A3(net884),
    .A4(net105),
    .B1(net108),
    .X(net120));
 sky130_fd_sc_hd__mux4_1 c283 (.A0(net118),
    .A1(net119),
    .A2(net739),
    .A3(net112),
    .S0(net884),
    .S1(net109),
    .X(net121));
 sky130_fd_sc_hd__a41o_2 c284 (.A1(net115),
    .A2(net118),
    .A3(net883),
    .A4(net108),
    .B1(net112),
    .X(net122));
 sky130_fd_sc_hd__mux4_2 c285 (.A0(net120),
    .A1(net122),
    .A2(net121),
    .A3(net103),
    .S0(net728),
    .S1(net118),
    .X(net123));
 sky130_fd_sc_hd__a21bo_2 c286 (.A1(net107),
    .A2(net104),
    .B1_N(net22),
    .X(net124));
 sky130_fd_sc_hd__a31o_1 c287 (.A1(net722),
    .A2(net887),
    .A3(net37),
    .B1(net31),
    .X(net125));
 sky130_fd_sc_hd__a21bo_2 c288 (.A1(net43),
    .A2(net109),
    .B1_N(net808),
    .X(net126));
 sky130_fd_sc_hd__a21bo_1 c289 (.A1(net113),
    .A2(net112),
    .B1_N(net889),
    .X(net127));
 sky130_fd_sc_hd__a21bo_1 c290 (.A1(net34),
    .A2(net120),
    .B1_N(net941),
    .X(net128));
 sky130_fd_sc_hd__a31o_1 c291 (.A1(net120),
    .A2(net128),
    .A3(net125),
    .B1(net901),
    .X(net129));
 sky130_fd_sc_hd__clkbuf_2 c292 (.A(net830),
    .X(net130));
 sky130_fd_sc_hd__a31o_4 c293 (.A1(net46),
    .A2(net125),
    .A3(net113),
    .B1(net889),
    .X(net131));
 sky130_fd_sc_hd__a41o_2 c294 (.A1(net39),
    .A2(net124),
    .A3(net750),
    .A4(net108),
    .B1(net127),
    .X(net850));
 sky130_fd_sc_hd__mux4_2 c295 (.A0(net41),
    .A1(net892),
    .A2(net130),
    .A3(net34),
    .S0(net39),
    .S1(net102),
    .X(net132));
 sky130_fd_sc_hd__a31o_4 c296 (.A1(net879),
    .A2(net130),
    .A3(net22),
    .B1(net726),
    .X(net133));
 sky130_fd_sc_hd__a31o_4 c297 (.A1(net130),
    .A2(net133),
    .A3(net879),
    .B1(net931),
    .X(net134));
 sky130_fd_sc_hd__sdfbbp_1 c298 (.CLK(clknet_4_7_0_clk),
    .D(net108),
    .RESET_B(net47),
    .SCD(net935),
    .SCE(net933),
    .SET_B(net130),
    .Q(net136),
    .Q_N(net135));
 sky130_fd_sc_hd__a31o_4 c299 (.A1(net770),
    .A2(net882),
    .A3(net905),
    .B1(net39),
    .X(net137));
 sky130_fd_sc_hd__a41o_1 c300 (.A1(net935),
    .A2(net102),
    .A3(net934),
    .A4(net135),
    .B1(net575),
    .X(net138));
 sky130_fd_sc_hd__a41o_1 c301 (.A1(net136),
    .A2(net130),
    .A3(net892),
    .A4(net730),
    .B1(net599),
    .X(net139));
 sky130_fd_sc_hd__mux4_2 c302 (.A0(net117),
    .A1(net46),
    .A2(net957),
    .A3(net935),
    .S0(net108),
    .S1(net599),
    .X(net140));
 sky130_fd_sc_hd__sdfrbp_1 c303 (.CLK(clknet_4_7_0_clk),
    .D(net127),
    .RESET_B(net140),
    .SCD(net137),
    .SCE(net134),
    .Q(net142),
    .Q_N(net141));
 sky130_fd_sc_hd__a31o_4 c304 (.A1(net850),
    .A2(net132),
    .A3(net736),
    .B1(net135),
    .X(net143));
 sky130_fd_sc_hd__mux4_2 c305 (.A0(net125),
    .A1(net143),
    .A2(net136),
    .A3(net141),
    .S0(net134),
    .X(net599));
 sky130_fd_sc_hd__a41o_1 c306 (.A1(net109),
    .A2(net41),
    .A3(net143),
    .A4(net128),
    .B1(net721),
    .X(net145));
 sky130_fd_sc_hd__mux4_2 c307 (.A0(net107),
    .A1(net127),
    .A2(net130),
    .A3(net143),
    .S0(net575),
    .S1(net928),
    .X(net146));
 sky130_fd_sc_hd__buf_1 c308 (.A(net607),
    .X(net147));
 sky130_fd_sc_hd__a21bo_1 c309 (.A1(net48),
    .A2(net885),
    .B1_N(net749),
    .X(net148));
 sky130_fd_sc_hd__a21bo_1 c310 (.A1(net49),
    .A2(net885),
    .B1_N(net941),
    .X(net149));
 sky130_fd_sc_hd__a31o_1 c311 (.A1(net148),
    .A2(net149),
    .A3(net124),
    .B1(net899),
    .X(net150));
 sky130_fd_sc_hd__clkbuf_2 c312 (.A(net607),
    .X(net151));
 sky130_fd_sc_hd__mux4_1 c313 (.A0(net60),
    .A1(net741),
    .A2(net883),
    .A3(net140),
    .S0(net37),
    .S1(net752),
    .X(net152));
 sky130_fd_sc_hd__mux4_1 c314 (.A0(net142),
    .A1(net762),
    .A2(net149),
    .A3(net879),
    .S0(net906),
    .S1(net899),
    .X(net153));
 sky130_fd_sc_hd__mux4_1 c315 (.A0(net746),
    .A1(net146),
    .A2(net148),
    .A3(net141),
    .S0(net902),
    .S1(net896),
    .X(net154));
 sky130_fd_sc_hd__a31o_1 c316 (.A1(net133),
    .A2(net762),
    .A3(net148),
    .B1(net153),
    .X(net155));
 sky130_fd_sc_hd__a21bo_2 c317 (.A1(net148),
    .A2(net52),
    .B1_N(net147),
    .X(net156));
 sky130_fd_sc_hd__sdfbbn_1 c318 (.CLK_N(clknet_4_7_0_clk),
    .D(net741),
    .RESET_B(net124),
    .SCD(net123),
    .SCE(net877),
    .SET_B(net899),
    .Q(net158),
    .Q_N(net157));
 sky130_fd_sc_hd__clkbuf_1 c319 (.A(net830),
    .X(net159));
 sky130_fd_sc_hd__a21bo_2 c320 (.A1(net153),
    .A2(net142),
    .B1_N(net899),
    .X(net160));
 sky130_fd_sc_hd__a21bo_1 c321 (.A1(net149),
    .A2(net157),
    .B1_N(net578),
    .X(net161));
 sky130_fd_sc_hd__mux4_1 c322 (.A0(net132),
    .A1(net37),
    .A2(net157),
    .A3(net156),
    .S0(net160),
    .S1(net877),
    .X(net162));
 sky130_fd_sc_hd__a21bo_1 c323 (.A1(net55),
    .A2(net158),
    .B1_N(net888),
    .X(net163));
 sky130_fd_sc_hd__clkbuf_1 c324 (.A(net630),
    .X(net164));
 sky130_fd_sc_hd__mux4_1 c325 (.A0(net164),
    .A1(net39),
    .A2(net160),
    .A3(net158),
    .S0(net745),
    .S1(net151),
    .X(net165));
 sky130_fd_sc_hd__a31o_1 c326 (.A1(net161),
    .A2(net163),
    .A3(net151),
    .B1(net899),
    .X(net166));
 sky130_fd_sc_hd__mux4_1 c327 (.A0(net154),
    .A1(net158),
    .A2(net166),
    .A3(net56),
    .S0(net142),
    .S1(net634),
    .X(net167));
 sky130_fd_sc_hd__mux4_1 c328 (.A0(net166),
    .A1(net160),
    .A2(net148),
    .A3(net50),
    .S0(net633),
    .S1(net635),
    .X(net168));
 sky130_fd_sc_hd__mux4_1 c329 (.A0(net159),
    .A1(net160),
    .A2(net133),
    .A3(net166),
    .S0(net579),
    .S1(net635),
    .X(net169));
 sky130_fd_sc_hd__mux4_1 c330 (.A0(net150),
    .A1(net752),
    .A2(net63),
    .A3(net80),
    .S0(net773),
    .S1(net28),
    .X(net170));
 sky130_fd_sc_hd__buf_1 c331 (.A(net626),
    .X(net171));
 sky130_fd_sc_hd__a41o_1 c332 (.A1(net80),
    .A2(net160),
    .A3(net877),
    .A4(net137),
    .B1(net48),
    .X(net172));
 sky130_fd_sc_hd__clkbuf_2 c333 (.A(net626),
    .X(net173));
 sky130_fd_sc_hd__a21bo_1 c334 (.A1(net771),
    .A2(net173),
    .B1_N(net840),
    .X(net174));
 sky130_fd_sc_hd__mux4_1 c335 (.A0(net747),
    .A1(net156),
    .A2(net22),
    .A3(net160),
    .S0(net80),
    .S1(net625),
    .X(net175));
 sky130_fd_sc_hd__a31o_1 c336 (.A1(net174),
    .A2(net879),
    .A3(net173),
    .B1(net591),
    .X(net176));
 sky130_fd_sc_hd__a21bo_1 c337 (.A1(net736),
    .A2(net176),
    .B1_N(net151),
    .X(net177));
 sky130_fd_sc_hd__sdfbbn_2 c338 (.CLK_N(clknet_4_12_0_clk),
    .D(net22),
    .RESET_B(net156),
    .SCD(net173),
    .SCE(net177),
    .SET_B(net747),
    .Q(net179),
    .Q_N(net178));
 sky130_fd_sc_hd__a31o_1 c339 (.A1(net747),
    .A2(net171),
    .A3(net850),
    .B1(net600),
    .X(net180));
 sky130_fd_sc_hd__a41o_1 c340 (.A1(net137),
    .A2(net180),
    .A3(net837),
    .A4(net178),
    .B1(net856),
    .X(net181));
 sky130_fd_sc_hd__a21bo_1 c341 (.A1(net52),
    .A2(net181),
    .B1_N(net817),
    .X(net182));
 sky130_fd_sc_hd__a21bo_2 c342 (.A1(net176),
    .A2(net48),
    .B1_N(net950),
    .X(net183));
 sky130_fd_sc_hd__a21bo_1 c343 (.A1(net179),
    .A2(net180),
    .B1_N(net625),
    .X(net184));
 sky130_fd_sc_hd__mux4_1 c344 (.A0(net173),
    .A1(net179),
    .A2(net180),
    .A3(net183),
    .S0(net181),
    .S1(net579),
    .X(net185));
 sky130_fd_sc_hd__sdfrbp_1 c345 (.CLK(clknet_4_14_0_clk),
    .D(net180),
    .RESET_B(net183),
    .SCD(net817),
    .SCE(net636),
    .Q(net187),
    .Q_N(net186));
 sky130_fd_sc_hd__mux4_1 c346 (.A0(net86),
    .A1(net182),
    .A2(net183),
    .A3(net186),
    .S0(net817),
    .S1(net636),
    .X(net188));
 sky130_fd_sc_hd__mux4_1 c347 (.A0(net181),
    .A1(net173),
    .A2(net183),
    .A3(net186),
    .S0(clknet_1_0__leaf_net604),
    .S1(clknet_1_1__leaf_net852),
    .X(net189));
 sky130_fd_sc_hd__mux4_1 c348 (.A0(net56),
    .A1(net174),
    .A2(net183),
    .A3(net598),
    .S1(clknet_1_0__leaf_net604),
    .X(net190));
 sky130_fd_sc_hd__a41o_1 c349 (.A1(net180),
    .A2(net598),
    .A3(net632),
    .A4(net636),
    .B1(clknet_1_0__leaf_net852),
    .X(net191));
 sky130_fd_sc_hd__mux4_1 c350 (.A0(net182),
    .A1(clknet_1_0__leaf_net191),
    .A2(net181),
    .A3(net160),
    .S0(net600),
    .S1(clknet_1_0__leaf_net852),
    .X(net192));
 sky130_fd_sc_hd__mux4_1 c351 (.A0(clknet_1_1__leaf_net191),
    .A1(net181),
    .A2(net156),
    .A3(net80),
    .S0(clknet_1_0__leaf_net852),
    .S1(clknet_1_1__leaf_net637),
    .X(net193));
 sky130_fd_sc_hd__a31o_1 c352 (.A1(net187),
    .A2(net835),
    .A3(net179),
    .B1(net801),
    .X(net844));
 sky130_fd_sc_hd__a41o_2 c353 (.A1(net844),
    .A2(net766),
    .A3(net726),
    .A4(net770),
    .B1(net882),
    .X(net819));
 sky130_fd_sc_hd__sdfbbp_1 c354 (.CLK(clknet_4_14_0_clk),
    .D(net171),
    .RESET_B(net801),
    .SCD(net907),
    .SCE(net183),
    .SET_B(clknet_1_0__leaf_net852),
    .Q(net195),
    .Q_N(net194));
 sky130_fd_sc_hd__sdfbbn_1 c355 (.CLK_N(clknet_4_14_0_clk),
    .D(net67),
    .RESET_B(net184),
    .SCD(net801),
    .SCE(clknet_1_0__leaf_net838),
    .SET_B(net897),
    .Q(net197),
    .Q_N(net196));
 sky130_fd_sc_hd__a31o_1 c356 (.A1(net87),
    .A2(net197),
    .A3(net849),
    .B1(net801),
    .X(net198));
 sky130_fd_sc_hd__sdfbbn_1 c357 (.CLK_N(clknet_4_14_0_clk),
    .D(net184),
    .RESET_B(net87),
    .SCD(net846),
    .SCE(net194),
    .SET_B(net198),
    .Q(net200),
    .Q_N(net199));
 sky130_fd_sc_hd__a31o_1 c358 (.A1(net768),
    .A2(net195),
    .A3(net92),
    .B1(net13),
    .X(net201));
 sky130_fd_sc_hd__mux4_1 c359 (.A0(net837),
    .A1(net903),
    .A2(net879),
    .A3(net768),
    .S0(net635),
    .S1(clknet_1_0__leaf_net852),
    .X(net841));
 sky130_fd_sc_hd__a31o_1 c360 (.A1(net183),
    .A2(net67),
    .A3(net101),
    .B1(net633),
    .X(net202));
 sky130_fd_sc_hd__a31o_1 c361 (.A1(net195),
    .A2(net885),
    .A3(net766),
    .B1(net851),
    .X(net822));
 sky130_fd_sc_hd__mux4_1 c362 (.A0(net160),
    .A1(net882),
    .A2(net67),
    .A3(net819),
    .S0(net184),
    .S1(net97),
    .X(net203));
 sky130_fd_sc_hd__a31o_1 c363 (.A1(net881),
    .A2(net773),
    .A3(net847),
    .B1(clknet_1_0__leaf_net638),
    .X(net204));
 sky130_fd_sc_hd__mux4_1 c364 (.A0(net758),
    .A1(clknet_1_1__leaf_net204),
    .A2(net801),
    .A3(net96),
    .S0(clknet_1_0__leaf_net841),
    .S1(clknet_1_0__leaf_net638),
    .X(net824));
 sky130_fd_sc_hd__mux4_1 c365 (.A0(net201),
    .A1(net196),
    .A2(clknet_1_0__leaf_net841),
    .A3(net101),
    .S0(net910),
    .S1(clknet_1_1__leaf_net638),
    .X(net205));
 sky130_fd_sc_hd__a41o_1 c366 (.A1(clknet_1_0__leaf_net204),
    .A2(net844),
    .A3(net881),
    .A4(net744),
    .B1(net630),
    .X(net816));
 sky130_fd_sc_hd__sdfrtn_1 c367 (.CLK_N(clknet_4_15_0_clk),
    .D(net771),
    .RESET_B(net945),
    .SCD(clknet_1_1__leaf_net824),
    .SCE(clknet_1_1__leaf_net816),
    .Q(net805));
 sky130_fd_sc_hd__mux4_1 c368 (.A0(net785),
    .A1(net909),
    .A2(net903),
    .A3(net771),
    .S0(net847),
    .S1(net630),
    .X(net206));
 sky130_fd_sc_hd__a41o_1 c369 (.A1(net784),
    .A2(net835),
    .A3(net881),
    .A4(net843),
    .B1(net630),
    .X(net845));
 sky130_fd_sc_hd__mux4_1 c370 (.A0(clknet_1_0__leaf_net816),
    .A1(net846),
    .A2(clknet_1_1__leaf_net838),
    .A3(net206),
    .S0(net843),
    .S1(clknet_1_1__leaf_net638),
    .X(net207));
 sky130_fd_sc_hd__mux4_1 c371 (.A0(net911),
    .A1(clknet_1_1__leaf_net841),
    .A2(net171),
    .A3(net97),
    .S0(clknet_1_1__leaf_net207),
    .S1(net634),
    .X(net208));
 sky130_fd_sc_hd__mux4_1 c372 (.A0(net206),
    .A1(net187),
    .A2(net845),
    .A3(clknet_1_1__leaf_net207),
    .S0(clknet_1_0__leaf_net816),
    .S1(net843),
    .X(net209));
 sky130_fd_sc_hd__mux4_1 c373 (.A0(net197),
    .A1(net28),
    .A2(clknet_1_1__leaf_net207),
    .A3(net206),
    .S0(net845),
    .S1(net639),
    .X(net210));
 sky130_fd_sc_hd__mux4_2 c396 (.A0(net28),
    .A1(net17),
    .A2(net892),
    .A3(net713),
    .S0(net715),
    .S1(net883),
    .X(net211));
 sky130_fd_sc_hd__a21bo_1 c397 (.A1(net121),
    .A2(net15),
    .B1_N(net25),
    .X(net212));
 sky130_fd_sc_hd__xnor2_4 c398 (.A(net890),
    .B(net905),
    .Y(net213));
 sky130_fd_sc_hd__xnor2_4 c399 (.A(net557),
    .B(net211),
    .Y(net214));
 sky130_fd_sc_hd__a41o_1 c400 (.A1(net213),
    .A2(net211),
    .A3(net212),
    .A4(net103),
    .B1(net707),
    .X(net215));
 sky130_fd_sc_hd__xnor2_1 c401 (.A(net105),
    .B(net213),
    .Y(net216));
 sky130_fd_sc_hd__dlymetal6s2s_1 c402 (.A(net576),
    .X(net217));
 sky130_fd_sc_hd__a31o_4 c403 (.A1(net213),
    .A2(net103),
    .A3(net114),
    .B1(net214),
    .X(net218));
 sky130_fd_sc_hd__a21bo_1 c404 (.A1(net17),
    .A2(net878),
    .B1_N(net211),
    .X(net219));
 sky130_fd_sc_hd__xnor2_2 c405 (.A(net21),
    .B(net886),
    .Y(net220));
 sky130_fd_sc_hd__xnor2_1 c406 (.A(net220),
    .B(net219),
    .Y(net221));
 sky130_fd_sc_hd__xnor2_2 c407 (.A(net219),
    .B(net213),
    .Y(net222));
 sky130_fd_sc_hd__mux4_1 c408 (.A0(net222),
    .A1(net21),
    .A2(net123),
    .A3(net17),
    .S0(net217),
    .S1(net213),
    .X(net223));
 sky130_fd_sc_hd__buf_2 c409 (.A(net576),
    .X(net224));
 sky130_fd_sc_hd__a21bo_1 c410 (.A1(net219),
    .A2(net224),
    .B1_N(net211),
    .X(net225));
 sky130_fd_sc_hd__clkbuf_4 c411 (.A(net622),
    .X(net226));
 sky130_fd_sc_hd__a21bo_1 c412 (.A1(net216),
    .A2(net224),
    .B1_N(net214),
    .X(net227));
 sky130_fd_sc_hd__buf_1 c413 (.A(net623),
    .X(net228));
 sky130_fd_sc_hd__mux4_1 c414 (.A0(net224),
    .A1(net222),
    .A2(net227),
    .A3(net219),
    .S0(net218),
    .S1(net958),
    .X(net229));
 sky130_fd_sc_hd__xnor2_2 c415 (.A(net218),
    .B(net226),
    .Y(net230));
 sky130_fd_sc_hd__clkbuf_4 c416 (.A(net622),
    .X(net231));
 sky130_fd_sc_hd__sdfbbp_1 c417 (.CLK(clknet_4_4_0_clk),
    .D(net230),
    .RESET_B(net225),
    .SCD(net224),
    .SCE(net214),
    .SET_B(net946),
    .Q(net233),
    .Q_N(net232));
 sky130_fd_sc_hd__a31o_1 c418 (.A1(net146),
    .A2(net218),
    .A3(net715),
    .B1(net575),
    .X(net234));
 sky130_fd_sc_hd__a21bo_1 c419 (.A1(net724),
    .A2(net139),
    .B1_N(net124),
    .X(net235));
 sky130_fd_sc_hd__clkbuf_1 c420 (.A(net589),
    .X(net236));
 sky130_fd_sc_hd__sdfbbn_1 c421 (.CLK_N(clknet_4_5_0_clk),
    .D(net143),
    .RESET_B(net12),
    .SCD(net225),
    .SCE(net31),
    .SET_B(net738),
    .Q(net238),
    .Q_N(net237));
 sky130_fd_sc_hd__a31o_1 c422 (.A1(net235),
    .A2(net122),
    .A3(net47),
    .B1(net238),
    .X(net239));
 sky130_fd_sc_hd__a41o_1 c423 (.A1(net139),
    .A2(net13),
    .A3(net932),
    .A4(net227),
    .B1(net143),
    .X(net240));
 sky130_fd_sc_hd__sdfbbn_1 c424 (.CLK_N(clknet_4_5_0_clk),
    .D(net37),
    .RESET_B(net235),
    .SCD(net146),
    .SCE(net876),
    .SET_B(net13),
    .Q(net242),
    .Q_N(net241));
 sky130_fd_sc_hd__a21bo_2 c425 (.A1(net236),
    .A2(net218),
    .B1_N(net224),
    .X(net848));
 sky130_fd_sc_hd__clkbuf_2 c426 (.A(net589),
    .X(net243));
 sky130_fd_sc_hd__sdfrtp_4 c427 (.CLK(clknet_4_5_0_clk),
    .D(net225),
    .RESET_B(net876),
    .SCD(net243),
    .SCE(net12),
    .Q(net244));
 sky130_fd_sc_hd__a21bo_1 c428 (.A1(net239),
    .A2(net143),
    .B1_N(net244),
    .X(net245));
 sky130_fd_sc_hd__sdfbbp_1 c429 (.CLK(clknet_4_7_0_clk),
    .D(net245),
    .RESET_B(net28),
    .SCD(net217),
    .SCE(net123),
    .SET_B(net240),
    .Q(net247),
    .Q_N(net246));
 sky130_fd_sc_hd__a31o_4 c430 (.A1(net235),
    .A2(net227),
    .A3(net104),
    .B1(net243),
    .X(net818));
 sky130_fd_sc_hd__sdfbbn_1 c431 (.CLK_N(clknet_4_7_0_clk),
    .D(net12),
    .RESET_B(net217),
    .SCD(net243),
    .SCE(net246),
    .SET_B(net245),
    .Q(net249),
    .Q_N(net248));
 sky130_fd_sc_hd__buf_1 c432 (.A(net620),
    .X(net250));
 sky130_fd_sc_hd__buf_1 c433 (.A(net611),
    .X(net251));
 sky130_fd_sc_hd__sdfbbn_1 c434 (.CLK_N(clknet_4_5_0_clk),
    .D(net216),
    .RESET_B(net953),
    .SCD(net217),
    .SCE(net247),
    .SET_B(net848),
    .Q(net253),
    .Q_N(net252));
 sky130_fd_sc_hd__a41o_2 c435 (.A1(net251),
    .A2(net252),
    .A3(net102),
    .A4(net239),
    .B1(net250),
    .X(net254));
 sky130_fd_sc_hd__mux4_1 c436 (.A0(net818),
    .A1(net254),
    .A2(net102),
    .A3(net243),
    .S0(net252),
    .S1(net576),
    .X(net255));
 sky130_fd_sc_hd__a41o_1 c437 (.A1(net250),
    .A2(net249),
    .A3(net251),
    .A4(net254),
    .B1(net645),
    .X(net256));
 sky130_fd_sc_hd__sdfbbp_1 c438 (.CLK(clknet_4_7_0_clk),
    .D(net738),
    .RESET_B(net250),
    .SCD(net248),
    .SCE(net818),
    .SET_B(net952),
    .Q(net258),
    .Q_N(net257));
 sky130_fd_sc_hd__mux4_2 c439 (.A0(net242),
    .A1(net253),
    .A2(net247),
    .A3(net248),
    .S0(net244),
    .S1(net257),
    .X(net259));
 sky130_fd_sc_hd__buf_1 c440 (.A(net705),
    .X(net260));
 sky130_fd_sc_hd__a31o_1 c441 (.A1(net713),
    .A2(net258),
    .A3(net37),
    .B1(net50),
    .X(net261));
 sky130_fd_sc_hd__clkbuf_4 c442 (.A(net705),
    .X(net262));
 sky130_fd_sc_hd__mux4_1 c443 (.A0(net243),
    .A1(net28),
    .A2(net230),
    .A3(net261),
    .S0(net248),
    .S1(net633),
    .X(net263));
 sky130_fd_sc_hd__clkbuf_1 c444 (.A(net619),
    .X(net264));
 sky130_fd_sc_hd__buf_1 c445 (.A(net629),
    .X(net265));
 sky130_fd_sc_hd__clkbuf_1 c446 (.A(net619),
    .X(net266));
 sky130_fd_sc_hd__mux4_1 c447 (.A0(net243),
    .A1(net151),
    .A2(net234),
    .A3(net259),
    .S0(net155),
    .S1(net608),
    .X(net267));
 sky130_fd_sc_hd__a21bo_1 c448 (.A1(net932),
    .A2(net251),
    .B1_N(net646),
    .X(net826));
 sky130_fd_sc_hd__sdfrtp_1 c449 (.CLK(clknet_4_12_0_clk),
    .D(net124),
    .RESET_B(net230),
    .SCD(net879),
    .SCE(net147),
    .Q(net268));
 sky130_fd_sc_hd__a21bo_1 c450 (.A1(net792),
    .A2(net882),
    .B1_N(net266),
    .X(net269));
 sky130_fd_sc_hd__a41o_2 c451 (.A1(net238),
    .A2(net726),
    .A3(net880),
    .A4(net265),
    .B1(net50),
    .X(net270));
 sky130_fd_sc_hd__mux4_2 c452 (.A0(net266),
    .A1(net270),
    .A2(net882),
    .A3(net572),
    .S0(net608),
    .S1(net646),
    .X(net271));
 sky130_fd_sc_hd__mux4_1 c453 (.A0(net224),
    .A1(net270),
    .A2(net155),
    .A3(net880),
    .S1(net635),
    .X(net272));
 sky130_fd_sc_hd__mux4_1 c454 (.A0(net217),
    .A1(net261),
    .A2(net271),
    .A3(net237),
    .S0(net124),
    .S1(net269),
    .X(net273));
 sky130_fd_sc_hd__mux4_1 c455 (.A0(net260),
    .A1(net261),
    .A2(net273),
    .A3(net268),
    .S0(net271),
    .S1(net264),
    .X(net274));
 sky130_fd_sc_hd__mux4_2 c456 (.A0(net249),
    .A1(net258),
    .A2(net762),
    .A3(net271),
    .S0(net246),
    .S1(net262),
    .X(net275));
 sky130_fd_sc_hd__mux4_1 c457 (.A0(net271),
    .A1(net37),
    .A2(net269),
    .A3(net155),
    .S0(net633),
    .S1(net954),
    .X(net276));
 sky130_fd_sc_hd__clkbuf_1 c458 (.A(net611),
    .X(net277));
 sky130_fd_sc_hd__a21bo_1 c459 (.A1(net260),
    .A2(net647),
    .B1_N(net648),
    .X(net278));
 sky130_fd_sc_hd__mux4_1 c460 (.A0(net147),
    .A1(net902),
    .A2(net254),
    .A3(net880),
    .S0(net275),
    .S1(net571),
    .X(net279));
 sky130_fd_sc_hd__mux4_1 c461 (.A0(net277),
    .A1(net826),
    .A2(net260),
    .A3(net278),
    .S0(net648),
    .S1(net649),
    .X(net280));
 sky130_fd_sc_hd__a21bo_1 c462 (.A1(net868),
    .A2(net233),
    .B1_N(net788),
    .X(net281));
 sky130_fd_sc_hd__a21bo_1 c463 (.A1(net137),
    .A2(net896),
    .B1_N(clknet_1_1__leaf_net637),
    .X(net282));
 sky130_fd_sc_hd__a21bo_1 c464 (.A1(clknet_1_0__leaf_net282),
    .A2(net903),
    .B1_N(net636),
    .X(net283));
 sky130_fd_sc_hd__buf_1 c465 (.A(net704),
    .X(net284));
 sky130_fd_sc_hd__a21bo_1 c466 (.A1(net281),
    .A2(net788),
    .B1_N(clknet_1_0__leaf_net637),
    .X(net285));
 sky130_fd_sc_hd__a21bo_1 c467 (.A1(net278),
    .A2(clknet_1_0__leaf_net282),
    .B1_N(net151),
    .X(net286));
 sky130_fd_sc_hd__a21bo_1 c468 (.A1(clknet_1_0__leaf_net282),
    .A2(net600),
    .B1_N(net636),
    .X(net287));
 sky130_fd_sc_hd__a21bo_1 c469 (.A1(net788),
    .A2(net880),
    .B1_N(net646),
    .X(net288));
 sky130_fd_sc_hd__mux4_1 c470 (.A0(net762),
    .A1(net224),
    .A2(net288),
    .A3(clknet_1_1__leaf_net286),
    .S0(net636),
    .S1(clknet_1_0__leaf_net637),
    .X(net289));
 sky130_fd_sc_hd__a21bo_1 c471 (.A1(clknet_1_0__leaf_net286),
    .A2(net281),
    .B1_N(net246),
    .X(net290));
 sky130_fd_sc_hd__a21bo_1 c472 (.A1(net283),
    .A2(net868),
    .B1_N(net646),
    .X(net291));
 sky130_fd_sc_hd__mux4_1 c473 (.A0(net173),
    .A1(clknet_1_1__leaf_net286),
    .A2(net275),
    .A3(net257),
    .S0(clknet_1_1__leaf_net282),
    .S1(net896),
    .X(net292));
 sky130_fd_sc_hd__a21bo_1 c474 (.A1(net247),
    .A2(net880),
    .B1_N(net288),
    .X(net293));
 sky130_fd_sc_hd__mux4_1 c475 (.A0(clknet_1_0__leaf_net290),
    .A1(clknet_1_1__leaf_net285),
    .A2(net257),
    .A3(clknet_1_0__leaf_net291),
    .S0(clknet_1_1__leaf_net286),
    .S1(net856),
    .X(net294));
 sky130_fd_sc_hd__mux4_1 c476 (.A0(net151),
    .A1(net284),
    .A2(clknet_1_0__leaf_net286),
    .A3(net262),
    .S0(clknet_1_0__leaf_net291),
    .S1(net896),
    .X(net295));
 sky130_fd_sc_hd__mux4_1 c477 (.A0(net259),
    .A1(clknet_1_1__leaf_net289),
    .A2(net773),
    .A3(clknet_1_1__leaf_net282),
    .S0(net284),
    .S1(net650),
    .X(net296));
 sky130_fd_sc_hd__mux4_1 c478 (.A0(net288),
    .A1(net726),
    .A2(net744),
    .A3(clknet_1_0__leaf_net291),
    .S0(net650),
    .S1(net652),
    .X(net297));
 sky130_fd_sc_hd__mux4_1 c479 (.A0(net293),
    .A1(clknet_1_1__leaf_net285),
    .A2(net173),
    .A3(clknet_1_0__leaf_net291),
    .S0(net651),
    .S1(net652),
    .X(net298));
 sky130_fd_sc_hd__clkbuf_1 c480 (.A(net703),
    .X(net299));
 sky130_fd_sc_hd__a41o_1 c481 (.A1(net299),
    .A2(net288),
    .A3(net13),
    .A4(net650),
    .B1(net653),
    .X(net300));
 sky130_fd_sc_hd__mux4_1 c482 (.A0(net273),
    .A1(net300),
    .A2(net856),
    .A3(net648),
    .S0(net652),
    .S1(net829),
    .X(net301));
 sky130_fd_sc_hd__mux4_1 c483 (.A0(clknet_1_0__leaf_net289),
    .A1(net787),
    .A2(net300),
    .A3(net830),
    .S0(net651),
    .S1(net832),
    .X(net302));
 sky130_fd_sc_hd__mux4_1 c484 (.A0(net881),
    .A1(net178),
    .A2(net868),
    .A3(net640),
    .S0(net641),
    .S1(net653),
    .X(net828));
 sky130_fd_sc_hd__mux4_2 c485 (.A0(net226),
    .A1(net200),
    .A2(net868),
    .A3(net881),
    .S0(net936),
    .S1(net817),
    .X(net303));
 sky130_fd_sc_hd__mux4_1 c486 (.A0(net92),
    .A1(net178),
    .A2(net903),
    .A3(net634),
    .S0(net817),
    .S1(net641),
    .X(net304));
 sky130_fd_sc_hd__mux4_1 c487 (.A0(net726),
    .A1(net773),
    .A2(clknet_1_0__leaf_net207),
    .A3(net304),
    .S0(net92),
    .S1(net823),
    .X(net305));
 sky130_fd_sc_hd__a41o_1 c488 (.A1(net938),
    .A2(net868),
    .A3(net818),
    .A4(net634),
    .B1(net639),
    .X(net306));
 sky130_fd_sc_hd__mux4_1 c489 (.A0(net303),
    .A1(net224),
    .A2(clknet_1_0__leaf_net816),
    .A3(net907),
    .S0(net787),
    .S1(net726),
    .X(net812));
 sky130_fd_sc_hd__mux4_1 c490 (.A0(clknet_1_0__leaf_net207),
    .A1(net834),
    .A2(clknet_1_1__leaf_net282),
    .A3(net28),
    .S0(net275),
    .S1(net610),
    .X(net307));
 sky130_fd_sc_hd__mux4_1 c491 (.A0(net201),
    .A1(clknet_1_1__leaf_net812),
    .A2(net101),
    .A3(net881),
    .S0(net640),
    .S1(clknet_1_1__leaf_net654),
    .X(net308));
 sky130_fd_sc_hd__mux4_1 c492 (.A0(net304),
    .A1(net92),
    .A2(net5),
    .A3(net937),
    .S0(net817),
    .S1(net832),
    .X(net309));
 sky130_fd_sc_hd__mux4_1 c493 (.A0(net818),
    .A1(clknet_1_1__leaf_net812),
    .A2(net868),
    .A3(net856),
    .S0(clknet_1_1__leaf_net654),
    .S1(clknet_1_1__leaf_net655),
    .X(net310));
 sky130_fd_sc_hd__mux4_1 c494 (.A0(net179),
    .A1(net97),
    .A2(net303),
    .A3(net819),
    .S0(net198),
    .S1(net627),
    .X(net311));
 sky130_fd_sc_hd__mux4_1 c495 (.A0(net198),
    .A1(net819),
    .A2(net627),
    .A3(net817),
    .S0(net833),
    .S1(clknet_1_1__leaf_net654),
    .X(net312));
 sky130_fd_sc_hd__mux4_1 c496 (.A0(net201),
    .A1(net198),
    .A2(net881),
    .A3(net5),
    .S0(net627),
    .S1(clknet_1_0__leaf_net656),
    .X(net313));
 sky130_fd_sc_hd__mux4_1 c497 (.A0(net773),
    .A1(net179),
    .A2(net199),
    .A3(net897),
    .S0(net610),
    .S1(clknet_1_0__leaf_net656),
    .X(net314));
 sky130_fd_sc_hd__mux4_1 c498 (.A0(net178),
    .A1(net201),
    .A2(net938),
    .A3(net571),
    .S0(net627),
    .S1(clknet_1_1__leaf_net656),
    .X(net315));
 sky130_fd_sc_hd__mux4_1 c499 (.A0(net303),
    .A1(net819),
    .A2(net178),
    .A3(net304),
    .S0(net787),
    .S1(net649),
    .X(net316));
 sky130_fd_sc_hd__mux4_1 c500 (.A0(net258),
    .A1(net834),
    .A2(net199),
    .A3(net897),
    .S0(net610),
    .S1(clknet_1_1__leaf_net655),
    .X(net317));
 sky130_fd_sc_hd__a41o_1 c501 (.A1(clknet_1_1__leaf_net317),
    .A2(net101),
    .A3(net881),
    .A4(clknet_1_0__leaf_net821),
    .B1(net817),
    .X(net318));
 sky130_fd_sc_hd__mux4_1 c502 (.A0(clknet_1_1__leaf_net282),
    .A1(clknet_1_1__leaf_net318),
    .A2(clknet_1_1__leaf_net317),
    .A3(net881),
    .S0(net856),
    .S1(clknet_1_1__leaf_net656),
    .X(net825));
 sky130_fd_sc_hd__mux4_1 c503 (.A0(net917),
    .A1(clknet_1_0__leaf_net314),
    .A2(clknet_1_0__leaf_net318),
    .A3(net787),
    .S0(net641),
    .S1(clknet_1_0__leaf_net654),
    .X(net319));
 sky130_fd_sc_hd__mux4_1 c504 (.A0(clknet_1_0__leaf_net314),
    .A1(clknet_1_0__leaf_net318),
    .A2(net881),
    .A3(clknet_1_1__leaf_net317),
    .S0(clknet_1_0__leaf_net654),
    .S1(clknet_1_1__leaf_net655),
    .X(net320));
 sky130_fd_sc_hd__mux4_1 c505 (.A0(net320),
    .A1(net319),
    .A2(clknet_1_1__leaf_net314),
    .A3(clknet_1_0__leaf_net824),
    .S0(clknet_1_1__leaf_net318),
    .S1(net770),
    .X(net321));
 sky130_fd_sc_hd__xnor2_1 c528 (.A(net25),
    .B(net232),
    .Y(net322));
 sky130_fd_sc_hd__xnor2_4 c529 (.A(net886),
    .B(net878),
    .Y(net323));
 sky130_fd_sc_hd__dlymetal6s2s_1 c530 (.A(net593),
    .X(net324));
 sky130_fd_sc_hd__xnor2_4 c531 (.A(net728),
    .B(net883),
    .Y(net325));
 sky130_fd_sc_hd__a21bo_4 c532 (.A1(net228),
    .A2(net214),
    .B1_N(net325),
    .X(net326));
 sky130_fd_sc_hd__buf_4 c533 (.A(net593),
    .X(net814));
 sky130_fd_sc_hd__a21bo_1 c534 (.A1(net322),
    .A2(net324),
    .B1_N(net326),
    .X(net327));
 sky130_fd_sc_hd__a31o_1 c535 (.A1(net707),
    .A2(net326),
    .A3(net322),
    .B1(net211),
    .X(net328));
 sky130_fd_sc_hd__dlymetal6s2s_1 c536 (.A(net592),
    .X(net329));
 sky130_fd_sc_hd__dlymetal6s2s_1 c537 (.A(net581),
    .X(net330));
 sky130_fd_sc_hd__sdfrtp_1 c538 (.CLK(clknet_4_4_0_clk),
    .D(net114),
    .RESET_B(net327),
    .SCD(net326),
    .SCE(net330),
    .Q(net331));
 sky130_fd_sc_hd__clkbuf_4 c539 (.A(net592),
    .X(net332));
 sky130_fd_sc_hd__mux4_1 c540 (.A0(net330),
    .A1(net327),
    .A2(net322),
    .A3(net323),
    .S0(net329),
    .S1(net218),
    .X(net333));
 sky130_fd_sc_hd__mux4_1 c541 (.A0(net323),
    .A1(net327),
    .A2(net15),
    .A3(net332),
    .S0(net231),
    .S1(net657),
    .X(net334));
 sky130_fd_sc_hd__a21bo_1 c542 (.A1(net330),
    .A2(net332),
    .B1_N(net644),
    .X(net335));
 sky130_fd_sc_hd__a21bo_1 c543 (.A1(net324),
    .A2(net326),
    .B1_N(net335),
    .X(net336));
 sky130_fd_sc_hd__mux4_1 c544 (.A0(net326),
    .A1(net330),
    .A2(net327),
    .A3(net335),
    .S0(net231),
    .S1(net660),
    .X(net337));
 sky130_fd_sc_hd__a21bo_2 c545 (.A1(net335),
    .A2(net814),
    .B1_N(net662),
    .X(net338));
 sky130_fd_sc_hd__mux4_2 c546 (.A0(net211),
    .A1(net323),
    .A2(net228),
    .A3(net891),
    .S0(net25),
    .S1(net332),
    .X(net339));
 sky130_fd_sc_hd__sdfbbn_1 c547 (.CLK_N(clknet_4_4_0_clk),
    .D(net103),
    .RESET_B(net956),
    .SCD(net336),
    .SCE(net339),
    .SET_B(net891),
    .Q(net341),
    .Q_N(net340));
 sky130_fd_sc_hd__a31o_1 c548 (.A1(net332),
    .A2(net231),
    .A3(net891),
    .B1(net340),
    .X(net342));
 sky130_fd_sc_hd__mux4_1 c549 (.A0(net328),
    .A1(net341),
    .A2(net339),
    .A3(net13),
    .S0(net342),
    .S1(net661),
    .X(net343));
 sky130_fd_sc_hd__a21bo_1 c550 (.A1(net964),
    .A2(net645),
    .B1_N(net658),
    .X(net344));
 sky130_fd_sc_hd__xnor2_4 c551 (.A(net326),
    .B(net721),
    .Y(net345));
 sky130_fd_sc_hd__clkbuf_2 c552 (.A(net613),
    .X(net346));
 sky130_fd_sc_hd__clkbuf_2 c553 (.A(net613),
    .X(net347));
 sky130_fd_sc_hd__xnor2_4 c554 (.A(net242),
    .B(net599),
    .Y(net348));
 sky130_fd_sc_hd__clkbuf_2 c555 (.A(net613),
    .X(net349));
 sky130_fd_sc_hd__a41o_1 c556 (.A1(net253),
    .A2(net226),
    .A3(net331),
    .A4(net964),
    .B1(net244),
    .X(net350));
 sky130_fd_sc_hd__a21bo_2 c557 (.A1(net102),
    .A2(net902),
    .B1_N(net232),
    .X(net351));
 sky130_fd_sc_hd__a21bo_1 c558 (.A1(net915),
    .A2(net351),
    .B1_N(net906),
    .X(net352));
 sky130_fd_sc_hd__sdfbbn_1 c559 (.CLK_N(clknet_4_4_0_clk),
    .D(net350),
    .RESET_B(net959),
    .SCD(net345),
    .SCE(net231),
    .SET_B(net122),
    .Q(net354),
    .Q_N(net353));
 sky130_fd_sc_hd__a21bo_1 c560 (.A1(net347),
    .A2(net244),
    .B1_N(net904),
    .X(net355));
 sky130_fd_sc_hd__xnor2_2 c561 (.A(net231),
    .B(net348),
    .Y(net356));
 sky130_fd_sc_hd__buf_1 c562 (.A(net706),
    .X(net357));
 sky130_fd_sc_hd__a41o_1 c563 (.A1(net356),
    .A2(net242),
    .A3(net31),
    .A4(net329),
    .B1(net942),
    .X(net358));
 sky130_fd_sc_hd__a31o_1 c564 (.A1(net354),
    .A2(net122),
    .A3(net347),
    .B1(net351),
    .X(net359));
 sky130_fd_sc_hd__clkbuf_2 c565 (.A(net613),
    .X(net360));
 sky130_fd_sc_hd__a41o_1 c566 (.A1(net359),
    .A2(net358),
    .A3(net350),
    .A4(net908),
    .B1(net351),
    .X(net361));
 sky130_fd_sc_hd__a21bo_1 c567 (.A1(net358),
    .A2(net349),
    .B1_N(net355),
    .X(net362));
 sky130_fd_sc_hd__mux4_2 c568 (.A0(net357),
    .A1(net244),
    .A2(net358),
    .A3(net908),
    .S0(net362),
    .S1(net929),
    .X(net363));
 sky130_fd_sc_hd__sdfbbp_1 c569 (.CLK(clknet_4_1_0_clk),
    .D(net362),
    .RESET_B(net913),
    .SCD(net955),
    .SCE(net347),
    .SET_B(net361),
    .Q(net804),
    .Q_N(net364));
 sky130_fd_sc_hd__a41o_1 c570 (.A1(net122),
    .A2(net361),
    .A3(net362),
    .A4(net804),
    .B1(net358),
    .X(net365));
 sky130_fd_sc_hd__a41o_1 c571 (.A1(net353),
    .A2(net363),
    .A3(net361),
    .A4(net358),
    .B1(net947),
    .X(net366));
 sky130_fd_sc_hd__mux4_1 c572 (.A0(net58),
    .A1(net914),
    .A2(net848),
    .A3(net891),
    .S0(net880),
    .S1(net648),
    .X(net367));
 sky130_fd_sc_hd__clkbuf_1 c573 (.A(net631),
    .X(net368));
 sky130_fd_sc_hd__a31o_1 c574 (.A1(net335),
    .A2(net814),
    .A3(net123),
    .B1(net664),
    .X(net369));
 sky130_fd_sc_hd__a21bo_1 c575 (.A1(net231),
    .A2(net280),
    .B1_N(net900),
    .X(net370));
 sky130_fd_sc_hd__buf_1 c576 (.A(net631),
    .X(net371));
 sky130_fd_sc_hd__clkbuf_1 c577 (.A(net620),
    .X(net372));
 sky130_fd_sc_hd__mux4_1 c578 (.A0(net814),
    .A1(net371),
    .A2(net921),
    .A3(net368),
    .S0(clknet_1_1__leaf_net605),
    .S1(net648),
    .X(net373));
 sky130_fd_sc_hd__sdfbbn_1 c579 (.CLK_N(clknet_4_3_0_clk),
    .D(net352),
    .RESET_B(net918),
    .SCD(net370),
    .SCE(net218),
    .SET_B(net894),
    .Q(net375),
    .Q_N(net374));
 sky130_fd_sc_hd__a21bo_1 c580 (.A1(net354),
    .A2(net324),
    .B1_N(net894),
    .X(net376));
 sky130_fd_sc_hd__mux4_1 c581 (.A0(net268),
    .A1(net376),
    .A2(net721),
    .A3(net137),
    .S0(clknet_1_0__leaf_net605),
    .S1(net894),
    .X(net377));
 sky130_fd_sc_hd__a31o_1 c582 (.A1(net331),
    .A2(net372),
    .A3(net370),
    .B1(net894),
    .X(net378));
 sky130_fd_sc_hd__a31o_1 c583 (.A1(net930),
    .A2(net715),
    .A3(net268),
    .B1(net894),
    .X(net379));
 sky130_fd_sc_hd__a31o_1 c584 (.A1(net378),
    .A2(net377),
    .A3(net376),
    .B1(net894),
    .X(net380));
 sky130_fd_sc_hd__mux4_2 c585 (.A0(net344),
    .A1(net352),
    .A2(clknet_1_1__leaf_net380),
    .A3(net363),
    .S0(net378),
    .S1(net894),
    .X(net381));
 sky130_fd_sc_hd__mux4_1 c586 (.A0(net379),
    .A1(net371),
    .A2(net378),
    .A3(net275),
    .S0(net347),
    .S1(clknet_1_1__leaf_net380),
    .X(net382));
 sky130_fd_sc_hd__mux4_1 c587 (.A0(net376),
    .A1(net375),
    .A2(net371),
    .A3(net912),
    .S0(clknet_1_1__leaf_net380),
    .S1(net666),
    .X(net383));
 sky130_fd_sc_hd__mux4_1 c588 (.A0(net848),
    .A1(net137),
    .A2(net218),
    .A3(net374),
    .S0(clknet_1_1__leaf_net380),
    .S1(net667),
    .X(net384));
 sky130_fd_sc_hd__a41o_1 c589 (.A1(net376),
    .A2(clknet_1_1__leaf_net380),
    .A3(net894),
    .A4(net668),
    .B1(net671),
    .X(net385));
 sky130_fd_sc_hd__mux4_1 c590 (.A0(net231),
    .A1(net268),
    .A2(net900),
    .A3(net590),
    .S0(net667),
    .S1(net670),
    .X(net386));
 sky130_fd_sc_hd__mux4_1 c591 (.A0(net877),
    .A1(net386),
    .A2(clknet_1_1__leaf_net380),
    .A3(net664),
    .S0(net669),
    .S1(net671),
    .X(net387));
 sky130_fd_sc_hd__mux4_1 c592 (.A0(net749),
    .A1(net336),
    .A2(clknet_1_1__leaf_net380),
    .A3(net848),
    .S0(net590),
    .S1(net670),
    .X(net388));
 sky130_fd_sc_hd__mux4_2 c593 (.A0(net371),
    .A1(net378),
    .A2(net811),
    .A3(net664),
    .S0(net667),
    .S1(net671),
    .X(net839));
 sky130_fd_sc_hd__clkbuf_1 c594 (.A(net702),
    .X(net389));
 sky130_fd_sc_hd__sdfbbn_1 c595 (.CLK_N(clknet_4_3_0_clk),
    .D(net918),
    .RESET_B(clknet_1_0__leaf_net285),
    .SCD(net848),
    .SCE(net374),
    .SET_B(net364),
    .Q(net391),
    .Q_N(net390));
 sky130_fd_sc_hd__a41o_1 c596 (.A1(net347),
    .A2(clknet_1_0__leaf_net285),
    .A3(net804),
    .A4(net346),
    .B1(net651),
    .X(net392));
 sky130_fd_sc_hd__clkbuf_4 c597 (.A(net701),
    .X(net393));
 sky130_fd_sc_hd__a21bo_1 c598 (.A1(net907),
    .A2(net346),
    .B1_N(net651),
    .X(net394));
 sky130_fd_sc_hd__a21bo_1 c599 (.A1(net300),
    .A2(net393),
    .B1_N(net770),
    .X(net395));
 sky130_fd_sc_hd__a31o_1 c600 (.A1(net233),
    .A2(clknet_1_0__leaf_net285),
    .A3(clknet_1_1__leaf_net392),
    .B1(net648),
    .X(net396));
 sky130_fd_sc_hd__a21bo_1 c601 (.A1(net368),
    .A2(net393),
    .B1_N(clknet_1_1__leaf_net396),
    .X(net397));
 sky130_fd_sc_hd__buf_1 c602 (.A(clknet_1_1__leaf_net605),
    .X(net398));
 sky130_fd_sc_hd__a21bo_1 c603 (.A1(net397),
    .A2(net923),
    .B1_N(net300),
    .X(net399));
 sky130_fd_sc_hd__a31o_1 c604 (.A1(clknet_1_0__leaf_net396),
    .A2(net13),
    .A3(net393),
    .B1(clknet_1_1__leaf_net392),
    .X(net400));
 sky130_fd_sc_hd__mux4_1 c605 (.A0(clknet_1_0__leaf_net285),
    .A1(net375),
    .A2(net749),
    .A3(net393),
    .S0(net808),
    .S1(net648),
    .X(net401));
 sky130_fd_sc_hd__a41o_1 c606 (.A1(net386),
    .A2(net848),
    .A3(net876),
    .A4(net904),
    .B1(net920),
    .X(net402));
 sky130_fd_sc_hd__mux4_1 c607 (.A0(net375),
    .A1(net884),
    .A2(net814),
    .A3(net391),
    .S0(net364),
    .S1(net651),
    .X(net403));
 sky130_fd_sc_hd__mux4_1 c608 (.A0(net403),
    .A1(net752),
    .A2(clknet_1_0__leaf_net291),
    .A3(net232),
    .S0(net393),
    .S1(net635),
    .X(net404));
 sky130_fd_sc_hd__buf_1 c609 (.A(clknet_1_0__leaf_net605),
    .X(net405));
 sky130_fd_sc_hd__dlymetal6s2s_1 c610 (.A(net706),
    .X(net803));
 sky130_fd_sc_hd__a41o_1 c611 (.A1(net339),
    .A2(net877),
    .A3(net393),
    .A4(net374),
    .B1(net635),
    .X(net406));
 sky130_fd_sc_hd__a21bo_1 c612 (.A1(net390),
    .A2(net810),
    .B1_N(net616),
    .X(net407));
 sky130_fd_sc_hd__mux4_1 c613 (.A0(net400),
    .A1(net407),
    .A2(net803),
    .A3(clknet_1_0__leaf_net291),
    .S0(net393),
    .S1(net895),
    .X(net408));
 sky130_fd_sc_hd__mux4_1 c614 (.A0(net405),
    .A1(clknet_1_1__leaf_net392),
    .A2(net752),
    .A3(clknet_1_0__leaf_net285),
    .S0(net349),
    .S1(net394),
    .X(net806));
 sky130_fd_sc_hd__mux4_1 c615 (.A0(net393),
    .A1(clknet_1_1__leaf_net392),
    .A2(net912),
    .A3(net803),
    .S0(net602),
    .S1(net616),
    .X(net807));
 sky130_fd_sc_hd__mux4_1 c616 (.A0(net908),
    .A1(net5),
    .A2(net346),
    .A3(net349),
    .S0(net390),
    .S1(net666),
    .X(net409));
 sky130_fd_sc_hd__a41o_1 c617 (.A1(clknet_1_1__leaf_net291),
    .A2(net200),
    .A3(net805),
    .A4(clknet_1_1__leaf_net317),
    .B1(net641),
    .X(net410));
 sky130_fd_sc_hd__a31o_1 c618 (.A1(net226),
    .A2(clknet_1_0__leaf_net317),
    .A3(clknet_1_1__leaf_net398),
    .B1(net642),
    .X(net411));
 sky130_fd_sc_hd__a41o_1 c619 (.A1(net233),
    .A2(clknet_1_0__leaf_net398),
    .A3(net642),
    .A4(clknet_1_0__leaf_net655),
    .B1(net666),
    .X(net809));
 sky130_fd_sc_hd__mux4_1 c620 (.A0(net349),
    .A1(net805),
    .A2(net346),
    .A3(net770),
    .S0(clknet_1_0__leaf_net809),
    .S1(clknet_1_0__leaf_net655),
    .X(net412));
 sky130_fd_sc_hd__mux4_1 c621 (.A0(net275),
    .A1(clknet_1_0__leaf_net317),
    .A2(net338),
    .A3(net349),
    .S0(clknet_1_0__leaf_net412),
    .S1(net635),
    .X(net413));
 sky130_fd_sc_hd__mux4_1 c622 (.A0(net908),
    .A1(clknet_1_0__leaf_net824),
    .A2(net5),
    .A3(clknet_1_1__leaf_net412),
    .S0(net882),
    .S1(net642),
    .X(net414));
 sky130_fd_sc_hd__mux4_1 c623 (.A0(net13),
    .A1(net922),
    .A2(net745),
    .A3(clknet_1_1__leaf_net812),
    .S0(net805),
    .S1(clknet_1_1__leaf_net655),
    .X(net415));
 sky130_fd_sc_hd__sdfbbp_1 c624 (.CLK(clknet_4_10_0_clk),
    .D(net5),
    .RESET_B(clknet_1_0__leaf_net412),
    .SCD(clknet_1_0__leaf_net812),
    .SCE(clknet_1_0__leaf_net317),
    .SET_B(net943),
    .Q(net417),
    .Q_N(net416));
 sky130_fd_sc_hd__mux4_1 c625 (.A0(net5),
    .A1(net882),
    .A2(clknet_1_0__leaf_net412),
    .A3(clknet_1_1__leaf_net291),
    .S0(net631),
    .S1(net943),
    .X(net418));
 sky130_fd_sc_hd__mux4_1 c626 (.A0(net200),
    .A1(net411),
    .A2(clknet_1_0__leaf_net809),
    .A3(net883),
    .S0(clknet_1_0__leaf_net412),
    .S1(net962),
    .X(net419));
 sky130_fd_sc_hd__mux4_1 c627 (.A0(clknet_1_0__leaf_net317),
    .A1(net5),
    .A2(clknet_1_1__leaf_net412),
    .A3(clknet_1_1__leaf_net809),
    .S0(net813),
    .S1(clknet_1_0__leaf_net655),
    .X(net420));
 sky130_fd_sc_hd__mux4_1 c628 (.A0(net419),
    .A1(clknet_1_1__leaf_net412),
    .A2(clknet_1_1__leaf_net812),
    .A3(clknet_1_0__leaf_net317),
    .S0(net814),
    .S1(net642),
    .X(net421));
 sky130_fd_sc_hd__mux4_1 c629 (.A0(clknet_1_0__leaf_net398),
    .A1(net417),
    .A2(net883),
    .A3(clknet_1_0__leaf_net317),
    .S0(clknet_1_0__leaf_net655),
    .S1(net666),
    .X(net422));
 sky130_fd_sc_hd__mux4_1 c630 (.A0(clknet_1_0__leaf_net412),
    .A1(net417),
    .A2(net883),
    .A3(net226),
    .S0(net5),
    .S1(clknet_1_1__leaf_net291),
    .X(net423));
 sky130_fd_sc_hd__mux4_1 c631 (.A0(net422),
    .A1(clknet_1_0__leaf_net809),
    .A2(clknet_1_0__leaf_net812),
    .A3(clknet_1_1__leaf_net291),
    .S0(net126),
    .S1(clknet_1_0__leaf_net317),
    .X(net424));
 sky130_fd_sc_hd__mux4_1 c632 (.A0(net346),
    .A1(net882),
    .A2(clknet_1_1__leaf_net809),
    .A3(net883),
    .S0(net615),
    .S1(net673),
    .X(net855));
 sky130_fd_sc_hd__mux4_1 c633 (.A0(net116),
    .A1(net416),
    .A2(clknet_1_0__leaf_net855),
    .A3(net815),
    .S0(net631),
    .S1(clknet_1_0__leaf_net655),
    .X(net425));
 sky130_fd_sc_hd__mux4_1 c634 (.A0(net425),
    .A1(clknet_1_0__leaf_net855),
    .A2(clknet_1_1__leaf_net420),
    .A3(clknet_1_0__leaf_net812),
    .S0(clknet_1_1__leaf_net412),
    .S1(net673),
    .X(net426));
 sky130_fd_sc_hd__mux4_1 c635 (.A0(clknet_1_0__leaf_net420),
    .A1(clknet_1_1__leaf_net291),
    .A2(clknet_1_1__leaf_net412),
    .A3(clknet_1_1__leaf_net855),
    .S0(clknet_1_0__leaf_net655),
    .S1(net674),
    .X(net427));
 sky130_fd_sc_hd__mux4_1 c636 (.A0(net389),
    .A1(net409),
    .A2(net808),
    .A3(clknet_1_0__leaf_net412),
    .S0(net226),
    .S1(net674),
    .X(net428));
 sky130_fd_sc_hd__mux4_1 c637 (.A0(net391),
    .A1(clknet_1_1__leaf_net412),
    .A2(clknet_1_0__leaf_net812),
    .A3(clknet_1_0__leaf_net824),
    .S0(net615),
    .S1(net674),
    .X(net429));
 sky130_fd_sc_hd__xnor2_1 c660 (.A(net233),
    .B(net15),
    .Y(net430));
 sky130_fd_sc_hd__xnor2_2 c661 (.A(net323),
    .B(net878),
    .Y(net431));
 sky130_fd_sc_hd__a21bo_2 c662 (.A1(net15),
    .A2(net878),
    .B1_N(net657),
    .X(net432));
 sky130_fd_sc_hd__a31o_1 c663 (.A1(net432),
    .A2(net884),
    .A3(net430),
    .B1(net925),
    .X(net433));
 sky130_fd_sc_hd__xnor2_4 c664 (.A(net332),
    .B(net432),
    .Y(net434));
 sky130_fd_sc_hd__buf_1 c665 (.A(net582),
    .X(net435));
 sky130_fd_sc_hd__clkbuf_4 c666 (.A(net582),
    .X(net436));
 sky130_fd_sc_hd__a21bo_4 c667 (.A1(net884),
    .A2(net323),
    .B1_N(net662),
    .X(net437));
 sky130_fd_sc_hd__clkbuf_2 c668 (.A(net581),
    .X(net438));
 sky130_fd_sc_hd__a21bo_1 c669 (.A1(net435),
    .A2(net436),
    .B1_N(net658),
    .X(net439));
 sky130_fd_sc_hd__buf_2 c670 (.A(net629),
    .X(net440));
 sky130_fd_sc_hd__a21bo_1 c671 (.A1(net430),
    .A2(net432),
    .B1_N(net435),
    .X(net441));
 sky130_fd_sc_hd__sdfbbn_1 c672 (.CLK_N(clknet_4_1_0_clk),
    .D(net435),
    .RESET_B(net441),
    .SCD(net438),
    .SCE(net432),
    .SET_B(net440),
    .Q(net443),
    .Q_N(net442));
 sky130_fd_sc_hd__sdfsbp_1 c673 (.CLK(clknet_4_0_0_clk),
    .D(net441),
    .SCD(net439),
    .SCE(net433),
    .SET_B(net442),
    .Q(net445),
    .Q_N(net444));
 sky130_fd_sc_hd__sdfsbp_1 c674 (.CLK(clknet_4_1_0_clk),
    .D(net443),
    .SCD(net438),
    .SCE(net436),
    .SET_B(net431),
    .Q(net447),
    .Q_N(net446));
 sky130_fd_sc_hd__a31o_1 c675 (.A1(net878),
    .A2(net446),
    .A3(net442),
    .B1(net444),
    .X(net448));
 sky130_fd_sc_hd__sdfstp_2 c676 (.CLK(clknet_4_0_0_clk),
    .D(net448),
    .SCD(net441),
    .SCE(net440),
    .SET_B(net332),
    .Q(net449));
 sky130_fd_sc_hd__sdfbbn_1 c677 (.CLK_N(clknet_4_0_0_clk),
    .D(net440),
    .RESET_B(net438),
    .SCD(net449),
    .SCE(net437),
    .SET_B(net960),
    .Q(net451),
    .Q_N(net450));
 sky130_fd_sc_hd__a41o_1 c678 (.A1(net451),
    .A2(net448),
    .A3(net449),
    .A4(net325),
    .B1(net663),
    .X(net452));
 sky130_fd_sc_hd__mux4_1 c679 (.A0(net452),
    .A1(net445),
    .A2(net450),
    .A3(net891),
    .S0(net449),
    .S1(net658),
    .X(net453));
 sky130_fd_sc_hd__mux4_1 c680 (.A0(net443),
    .A1(net451),
    .A2(net448),
    .A3(net438),
    .S0(net452),
    .S1(net657),
    .X(net454));
 sky130_fd_sc_hd__mux4_1 c681 (.A0(net452),
    .A1(net443),
    .A2(net325),
    .A3(net341),
    .S0(net450),
    .S1(clknet_1_0__leaf_net677),
    .X(net455));
 sky130_fd_sc_hd__mux4_1 c682 (.A0(net449),
    .A1(net137),
    .A2(net439),
    .A3(net876),
    .S0(net434),
    .S1(net906),
    .X(net456));
 sky130_fd_sc_hd__a41o_1 c683 (.A1(net434),
    .A2(net112),
    .A3(net137),
    .A4(net663),
    .B1(clknet_1_1__leaf_net676),
    .X(net457));
 sky130_fd_sc_hd__a31o_1 c684 (.A1(net445),
    .A2(net351),
    .A3(net439),
    .B1(net434),
    .X(net458));
 sky130_fd_sc_hd__a31o_1 c685 (.A1(net439),
    .A2(net628),
    .A3(net659),
    .B1(clknet_1_0__leaf_net676),
    .X(net459));
 sky130_fd_sc_hd__sdfstp_1 c686 (.CLK(clknet_4_0_0_clk),
    .D(net437),
    .SCD(clknet_1_1__leaf_net459),
    .SCE(net947),
    .SET_B(net944),
    .Q(net460));
 sky130_fd_sc_hd__a31o_1 c687 (.A1(net351),
    .A2(net434),
    .A3(net876),
    .B1(clknet_1_0__leaf_net459),
    .X(net461));
 sky130_fd_sc_hd__mux4_1 c688 (.A0(net345),
    .A1(net444),
    .A2(net438),
    .A3(net340),
    .S0(net663),
    .S1(clknet_1_0__leaf_net676),
    .X(net462));
 sky130_fd_sc_hd__a21bo_1 c689 (.A1(net439),
    .A2(net445),
    .B1_N(clknet_1_0__leaf_net677),
    .X(net463));
 sky130_fd_sc_hd__mux4_1 c690 (.A0(net218),
    .A1(net436),
    .A2(net876),
    .A3(net345),
    .S0(net628),
    .S1(clknet_1_1__leaf_net677),
    .X(net464));
 sky130_fd_sc_hd__buf_1 c691 (.A(net552),
    .X(net465));
 sky130_fd_sc_hd__a21bo_1 c692 (.A1(net325),
    .A2(clknet_1_0__leaf_net459),
    .B1_N(net438),
    .X(net466));
 sky130_fd_sc_hd__a21bo_1 c693 (.A1(clknet_1_1__leaf_net466),
    .A2(net360),
    .B1_N(net658),
    .X(net467));
 sky130_fd_sc_hd__mux4_2 c694 (.A0(net884),
    .A1(net112),
    .A2(net891),
    .A3(net446),
    .S0(net436),
    .S1(net660),
    .X(net468));
 sky130_fd_sc_hd__a31o_1 c695 (.A1(net951),
    .A2(net876),
    .A3(net351),
    .B1(net678),
    .X(net469));
 sky130_fd_sc_hd__buf_1 c696 (.A(net551),
    .X(net470));
 sky130_fd_sc_hd__mux4_2 c697 (.A0(net465),
    .A1(net436),
    .A2(net468),
    .A3(net341),
    .S0(net629),
    .S1(net680),
    .X(net471));
 sky130_fd_sc_hd__a21bo_1 c698 (.A1(net465),
    .A2(net468),
    .B1_N(net574),
    .X(net472));
 sky130_fd_sc_hd__mux4_1 c699 (.A0(net467),
    .A1(net470),
    .A2(net439),
    .A3(net471),
    .S0(net612),
    .S1(net663),
    .X(net473));
 sky130_fd_sc_hd__mux4_1 c700 (.A0(net341),
    .A1(net472),
    .A2(net449),
    .A3(clknet_1_0__leaf_net473),
    .S0(net437),
    .S1(net434),
    .X(net474));
 sky130_fd_sc_hd__mux4_1 c701 (.A0(net355),
    .A1(net470),
    .A2(net472),
    .A3(net449),
    .S0(clknet_1_0__leaf_net473),
    .S1(clknet_1_0__leaf_net466),
    .X(net475));
 sky130_fd_sc_hd__mux4_1 c702 (.A0(net470),
    .A1(clknet_1_0__leaf_net473),
    .A2(clknet_1_1__leaf_net459),
    .A3(net472),
    .S0(net465),
    .S1(net682),
    .X(net476));
 sky130_fd_sc_hd__mux4_1 c703 (.A0(net471),
    .A1(net470),
    .A2(net437),
    .A3(net472),
    .S0(net683),
    .S1(net684),
    .X(net477));
 sky130_fd_sc_hd__mux4_1 c704 (.A0(net137),
    .A1(net906),
    .A2(net900),
    .A3(clknet_1_1__leaf_net380),
    .S0(net573),
    .S1(net894),
    .X(net478));
 sky130_fd_sc_hd__sdfbbp_1 c705 (.CLK(clknet_4_2_0_clk),
    .D(net360),
    .RESET_B(net900),
    .SCD(clknet_1_0__leaf_net380),
    .SCE(net678),
    .SET_B(net684),
    .Q(net480),
    .Q_N(net479));
 sky130_fd_sc_hd__a41o_1 c706 (.A1(clknet_1_1__leaf_net380),
    .A2(net218),
    .A3(net471),
    .A4(net900),
    .B1(net894),
    .X(net481));
 sky130_fd_sc_hd__mux4_1 c707 (.A0(net460),
    .A1(clknet_1_0__leaf_net463),
    .A2(net472),
    .A3(net891),
    .S0(net360),
    .S1(net436),
    .X(net482));
 sky130_fd_sc_hd__sdfbbn_1 c708 (.CLK_N(clknet_4_3_0_clk),
    .D(net270),
    .RESET_B(net440),
    .SCD(clknet_1_1__leaf_net380),
    .SCE(net28),
    .SET_B(net893),
    .Q(net484),
    .Q_N(net483));
 sky130_fd_sc_hd__clkbuf_1 c709 (.A(net623),
    .X(net485));
 sky130_fd_sc_hd__mux4_1 c710 (.A0(clknet_1_1__leaf_net459),
    .A1(net880),
    .A2(net900),
    .A3(clknet_1_1__leaf_net482),
    .S0(clknet_1_0__leaf_net380),
    .S1(net218),
    .X(net486));
 sky130_fd_sc_hd__mux4_1 c711 (.A0(net436),
    .A1(net882),
    .A2(net876),
    .A3(net460),
    .S0(net904),
    .S1(net684),
    .X(net487));
 sky130_fd_sc_hd__a41o_1 c712 (.A1(net472),
    .A2(clknet_1_0__leaf_net482),
    .A3(net577),
    .A4(net681),
    .B1(net687),
    .X(net488));
 sky130_fd_sc_hd__mux4_2 c713 (.A0(net440),
    .A1(net360),
    .A2(net635),
    .A3(net679),
    .S0(net685),
    .S1(net687),
    .X(net489));
 sky130_fd_sc_hd__mux4_1 c714 (.A0(net471),
    .A1(net440),
    .A2(net489),
    .A3(clknet_1_1__leaf_net473),
    .S0(net262),
    .S1(net893),
    .X(net490));
 sky130_fd_sc_hd__mux4_1 c715 (.A0(net342),
    .A1(clknet_1_1__leaf_net488),
    .A2(net468),
    .A3(clknet_1_1__leaf_net380),
    .S0(net900),
    .S1(net686),
    .X(net491));
 sky130_fd_sc_hd__mux4_1 c716 (.A0(net900),
    .A1(net360),
    .A2(net483),
    .A3(clknet_1_0__leaf_net488),
    .S0(net436),
    .S1(clknet_1_0__leaf_net380),
    .X(net492));
 sky130_fd_sc_hd__mux4_1 c717 (.A0(net465),
    .A1(net484),
    .A2(net468),
    .A3(clknet_1_1__leaf_net488),
    .S0(net436),
    .S1(net691),
    .X(net493));
 sky130_fd_sc_hd__sdfbbn_1 c718 (.CLK_N(clknet_4_2_0_clk),
    .D(net265),
    .RESET_B(clknet_1_0__leaf_net380),
    .SCD(net489),
    .SCE(net687),
    .SET_B(net693),
    .Q(net495),
    .Q_N(net494));
 sky130_fd_sc_hd__mux4_1 c719 (.A0(net900),
    .A1(net904),
    .A2(clknet_1_0__leaf_net380),
    .A3(net577),
    .S0(net687),
    .S1(net692),
    .X(net496));
 sky130_fd_sc_hd__mux4_1 c720 (.A0(net495),
    .A1(clknet_1_0__leaf_net482),
    .A2(net436),
    .A3(clknet_1_0__leaf_net380),
    .S0(net685),
    .S1(net694),
    .X(net497));
 sky130_fd_sc_hd__mux4_1 c721 (.A0(net485),
    .A1(clknet_1_0__leaf_net380),
    .A2(net495),
    .A3(net880),
    .S0(net646),
    .S1(net695),
    .X(net498));
 sky130_fd_sc_hd__mux4_1 c722 (.A0(net270),
    .A1(net494),
    .A2(net628),
    .A3(net893),
    .S0(net693),
    .S1(net695),
    .X(net499));
 sky130_fd_sc_hd__mux4_1 c723 (.A0(net360),
    .A1(net628),
    .A2(net686),
    .A3(net687),
    .S0(net694),
    .S1(net695),
    .X(net500));
 sky130_fd_sc_hd__mux4_1 c724 (.A0(clknet_1_0__leaf_net488),
    .A1(net500),
    .A2(net499),
    .A3(net440),
    .S0(clknet_1_0__leaf_net380),
    .S1(net679),
    .X(net501));
 sky130_fd_sc_hd__mux4_1 c725 (.A0(net499),
    .A1(net500),
    .A2(net494),
    .A3(net612),
    .S0(net679),
    .S1(clknet_1_0__leaf_net696),
    .X(net502));
 sky130_fd_sc_hd__a41o_1 c726 (.A1(net489),
    .A2(net437),
    .A3(net877),
    .A4(net646),
    .B1(net690),
    .X(net503));
 sky130_fd_sc_hd__a41o_1 c727 (.A1(clknet_1_1__leaf_net401),
    .A2(net143),
    .A3(net394),
    .A4(net904),
    .B1(net895),
    .X(net504));
 sky130_fd_sc_hd__mux4_1 c728 (.A0(net876),
    .A1(net721),
    .A2(net446),
    .A3(net882),
    .S0(net688),
    .S1(clknet_1_0__leaf_net696),
    .X(net505));
 sky130_fd_sc_hd__mux4_1 c729 (.A0(net468),
    .A1(net447),
    .A2(net28),
    .A3(net232),
    .S0(net893),
    .S1(net684),
    .X(net506));
 sky130_fd_sc_hd__mux4_1 c730 (.A0(net123),
    .A1(net484),
    .A2(clknet_1_1__leaf_net463),
    .A3(net232),
    .S0(net262),
    .S1(clknet_1_0__leaf_net504),
    .X(net507));
 sky130_fd_sc_hd__a41o_1 c731 (.A1(net394),
    .A2(clknet_1_1__leaf_net473),
    .A3(net884),
    .A4(net262),
    .B1(net893),
    .X(net508));
 sky130_fd_sc_hd__a41o_1 c732 (.A1(net472),
    .A2(net721),
    .A3(net483),
    .A4(net479),
    .B1(net893),
    .X(net509));
 sky130_fd_sc_hd__a41o_1 c733 (.A1(net447),
    .A2(net440),
    .A3(net907),
    .A4(net893),
    .B1(net688),
    .X(net510));
 sky130_fd_sc_hd__mux4_1 c734 (.A0(clknet_1_1__leaf_net504),
    .A1(net814),
    .A2(net891),
    .A3(net510),
    .S0(net602),
    .S1(net895),
    .X(net511));
 sky130_fd_sc_hd__a41o_1 c735 (.A1(clknet_1_0__leaf_net504),
    .A2(net876),
    .A3(net646),
    .A4(net893),
    .B1(net684),
    .X(net512));
 sky130_fd_sc_hd__a41o_1 c736 (.A1(net489),
    .A2(net510),
    .A3(net908),
    .A4(net880),
    .B1(net689),
    .X(net513));
 sky130_fd_sc_hd__a41o_1 c737 (.A1(net262),
    .A2(net764),
    .A3(clknet_1_0__leaf_net511),
    .A4(net595),
    .B1(net689),
    .X(net514));
 sky130_fd_sc_hd__sdfbbp_1 c738 (.CLK(clknet_4_8_0_clk),
    .D(net721),
    .RESET_B(net123),
    .SCD(clknet_1_0__leaf_net392),
    .SCE(net618),
    .SET_B(net895),
    .Q(net516),
    .Q_N(net515));
 sky130_fd_sc_hd__a41o_1 c739 (.A1(net880),
    .A2(net506),
    .A3(net510),
    .A4(net489),
    .B1(clknet_1_0__leaf_net401),
    .X(net517));
 sky130_fd_sc_hd__sdfbbn_1 c740 (.CLK_N(clknet_4_2_0_clk),
    .D(clknet_1_0__leaf_net502),
    .RESET_B(net517),
    .SCD(net515),
    .SCE(clknet_1_1__leaf_net473),
    .SET_B(net893),
    .Q(net519),
    .Q_N(net518));
 sky130_fd_sc_hd__a41o_1 c741 (.A1(net516),
    .A2(clknet_1_1__leaf_net502),
    .A3(net518),
    .A4(clknet_1_0__leaf_net392),
    .B1(net685),
    .X(net520));
 sky130_fd_sc_hd__mux4_1 c742 (.A0(net484),
    .A1(net447),
    .A2(net510),
    .A3(net907),
    .S0(net893),
    .S1(clknet_1_0__leaf_net696),
    .X(net521));
 sky130_fd_sc_hd__mux4_1 c743 (.A0(net884),
    .A1(net519),
    .A2(net468),
    .A3(net516),
    .S0(clknet_1_0__leaf_net521),
    .S1(net695),
    .X(net522));
 sky130_fd_sc_hd__mux4_1 c744 (.A0(clknet_1_1__leaf_net473),
    .A1(clknet_1_1__leaf_net522),
    .A2(net233),
    .A3(net515),
    .S0(clknet_1_0__leaf_net521),
    .S1(net646),
    .X(net523));
 sky130_fd_sc_hd__mux4_1 c745 (.A0(clknet_1_1__leaf_net463),
    .A1(net509),
    .A2(clknet_1_0__leaf_net522),
    .A3(net440),
    .S0(clknet_1_0__leaf_net521),
    .S1(clknet_1_0__leaf_net696),
    .X(net524));
 sky130_fd_sc_hd__mux4_1 c746 (.A0(net524),
    .A1(clknet_1_0__leaf_net522),
    .A2(net468),
    .A3(net594),
    .S0(net685),
    .S1(net695),
    .X(net525));
 sky130_fd_sc_hd__mux4_1 c747 (.A0(clknet_1_0__leaf_net401),
    .A1(clknet_1_0__leaf_net392),
    .A2(clknet_1_1__leaf_net522),
    .A3(net617),
    .S0(net618),
    .S1(net629),
    .X(net526));
 sky130_fd_sc_hd__mux4_1 c748 (.A0(clknet_1_0__leaf_net526),
    .A1(net480),
    .A2(clknet_1_0__leaf_net392),
    .A3(net617),
    .S0(net688),
    .S1(net695),
    .X(net527));
 sky130_fd_sc_hd__mux4_1 c749 (.A0(clknet_1_1__leaf_net521),
    .A1(net527),
    .A2(net437),
    .A3(clknet_1_0__leaf_net526),
    .S0(clknet_1_0__leaf_net675),
    .S1(clknet_1_1__leaf_net696),
    .X(net528));
 sky130_fd_sc_hd__mux4_1 c750 (.A0(clknet_1_1__leaf_net511),
    .A1(net416),
    .A2(net635),
    .A3(net674),
    .S0(net690),
    .S1(net695),
    .X(net529));
 sky130_fd_sc_hd__mux4_1 c751 (.A0(net480),
    .A1(clknet_1_1__leaf_net392),
    .A2(clknet_1_1__leaf_net526),
    .A3(clknet_1_1__leaf_net521),
    .S0(net674),
    .S1(net690),
    .X(net530));
 sky130_fd_sc_hd__mux4_1 c752 (.A0(net940),
    .A1(clknet_1_0__leaf_net392),
    .A2(clknet_1_0__leaf_net675),
    .A3(net695),
    .S0(clknet_1_1__leaf_net696),
    .S1(clknet_1_1__leaf_net697),
    .X(net531));
 sky130_fd_sc_hd__mux4_1 c753 (.A0(net530),
    .A1(clknet_1_0__leaf_net392),
    .A2(net814),
    .A3(net877),
    .S0(clknet_1_1__leaf_net526),
    .S1(clknet_1_1__leaf_net696),
    .X(net532));
 sky130_fd_sc_hd__mux4_1 c754 (.A0(net126),
    .A1(net764),
    .A2(net13),
    .A3(net904),
    .S0(clknet_1_0__leaf_net697),
    .S1(clknet_1_0__leaf_net698),
    .X(net533));
 sky130_fd_sc_hd__mux4_1 c755 (.A0(net437),
    .A1(net428),
    .A2(net480),
    .A3(clknet_1_0__leaf_net526),
    .S0(clknet_1_1__leaf_net697),
    .S1(clknet_1_1__leaf_net698),
    .X(net534));
 sky130_fd_sc_hd__mux4_1 c756 (.A0(net533),
    .A1(net891),
    .A2(net597),
    .A3(clknet_1_1__leaf_net675),
    .S0(net695),
    .S1(clknet_1_0__leaf_net698),
    .X(net535));
 sky130_fd_sc_hd__mux4_1 c757 (.A0(net531),
    .A1(net764),
    .A2(clknet_1_1__leaf_net526),
    .A3(clknet_1_0__leaf_net392),
    .S0(clknet_1_1__leaf_net698),
    .S1(net700),
    .X(net536));
 sky130_fd_sc_hd__mux4_1 c758 (.A0(clknet_1_0__leaf_net392),
    .A1(net417),
    .A2(clknet_1_1__leaf_net696),
    .A3(clknet_1_1__leaf_net697),
    .S0(clknet_1_0__leaf_net698),
    .S1(net699),
    .X(net537));
 sky130_fd_sc_hd__mux4_1 c759 (.A0(net877),
    .A1(net513),
    .A2(net770),
    .A3(clknet_1_1__leaf_net526),
    .S0(net823),
    .S1(clknet_1_1__leaf_net698),
    .X(net538));
 sky130_fd_sc_hd__mux4_1 c760 (.A0(net536),
    .A1(clknet_1_0__leaf_net392),
    .A2(net479),
    .A3(net823),
    .S0(clknet_1_1__leaf_net675),
    .S1(clknet_1_0__leaf_net698),
    .X(net539));
 sky130_fd_sc_hd__mux4_1 c761 (.A0(net764),
    .A1(net535),
    .A2(clknet_1_1__leaf_net521),
    .A3(net596),
    .S0(clknet_1_0__leaf_net697),
    .S1(clknet_1_0__leaf_net698),
    .X(net540));
 sky130_fd_sc_hd__mux4_1 c762 (.A0(net891),
    .A1(net537),
    .A2(net540),
    .A3(clknet_1_0__leaf_net392),
    .S0(clknet_1_1__leaf_net675),
    .S1(clknet_1_0__leaf_net698));
 sky130_fd_sc_hd__a41o_1 merge763 (.A1(net220),
    .A2(net123),
    .A3(net47),
    .A4(net241),
    .B1(net949),
    .X(net541));
 sky130_fd_sc_hd__a41o_1 merge764 (.A1(net156),
    .A2(net48),
    .A3(net883),
    .A4(net63),
    .B1(net747),
    .X(net542));
 sky130_fd_sc_hd__mux4_1 merge765 (.A0(net914),
    .A1(net234),
    .A2(net808),
    .A3(net370),
    .S0(net921),
    .S1(net110),
    .X(net543));
 sky130_fd_sc_hd__mux4_1 merge766 (.A0(net177),
    .A1(net173),
    .A2(clknet_1_0__leaf_net282),
    .A3(net287),
    .S0(clknet_1_1__leaf_net290),
    .S1(net749),
    .X(net544));
 sky130_fd_sc_hd__mux4_1 merge767 (.A0(net140),
    .A1(net763),
    .A2(net899),
    .A3(net742),
    .S0(net150),
    .S1(net148),
    .X(net545));
 sky130_fd_sc_hd__mux4_1 merge768 (.A0(net212),
    .A1(net231),
    .A2(net324),
    .A3(net878),
    .S0(net123),
    .S1(net643),
    .X(net546));
 sky130_fd_sc_hd__mux4_1 merge769 (.A0(net67),
    .A1(net796),
    .A2(clknet_1_1__leaf_net94),
    .A3(clknet_1_0__leaf_net862),
    .S0(clknet_1_1__leaf_net836),
    .S1(net897),
    .X(net547));
 sky130_fd_sc_hd__mux4_1 merge770 (.A0(net254),
    .A1(net58),
    .A2(net240),
    .A3(net230),
    .S0(net260),
    .S1(net726),
    .X(net548));
 sky130_fd_sc_hd__a31o_1 merge771 (.A1(net212),
    .A2(net216),
    .A3(net221),
    .B1(net621),
    .X(net549));
 sky130_fd_sc_hd__a41o_1 merge772 (.A1(net430),
    .A2(net433),
    .A3(net434),
    .A4(net435),
    .B1(net663),
    .X(net550));
 sky130_fd_sc_hd__sdfbbn_1 merge773 (.CLK_N(clknet_4_1_0_clk),
    .D(net112),
    .RESET_B(net434),
    .SCD(net345),
    .SCE(clknet_1_0__leaf_net463),
    .SET_B(net624),
    .Q(net552),
    .Q_N(net551));
 sky130_fd_sc_hd__a41o_1 merge774 (.A1(net123),
    .A2(net345),
    .A3(net340),
    .A4(net575),
    .B1(net663),
    .X(net553));
 sky130_fd_sc_hd__mux4_1 merge775 (.A0(net71),
    .A1(net777),
    .A2(net70),
    .A3(net907),
    .S0(clknet_1_0__leaf_net75),
    .S1(net896),
    .X(net554));
 sky130_fd_sc_hd__mux4_1 merge776 (.A0(net336),
    .A1(net902),
    .A2(net900),
    .A3(net877),
    .S0(net635),
    .S1(net961),
    .X(net555));
 sky130_fd_sc_hd__mux4_1 merge777 (.A0(clknet_1_0__leaf_net836),
    .A1(net76),
    .A2(net73),
    .A3(net72),
    .S0(net851),
    .S1(net632),
    .X(net556));
 sky130_fd_sc_hd__a31o_1 merge778 (.A1(net225),
    .A2(net222),
    .A3(net220),
    .X(net621));
 sky130_fd_sc_hd__mux4_1 merge779 (.A0(net393),
    .A1(net300),
    .A2(clknet_1_0__leaf_net291),
    .A3(net241),
    .S0(net345),
    .S1(net338),
    .X(net558));
 sky130_fd_sc_hd__mux4_1 merge780 (.A0(net227),
    .A1(net245),
    .A2(net104),
    .A3(net280),
    .S0(net919),
    .S1(net344),
    .X(net559));
 sky130_fd_sc_hd__mux4_1 merge781 (.A0(net128),
    .A1(net34),
    .A2(net123),
    .A3(net157),
    .S0(net132),
    .S1(net156),
    .X(net560));
 sky130_fd_sc_hd__a41o_1 merge782 (.A1(net399),
    .A2(net393),
    .A3(net839),
    .A4(net395),
    .B1(net650),
    .X(net561));
 sky130_fd_sc_hd__mux4_1 merge783 (.A0(net104),
    .A1(net250),
    .A2(net818),
    .A3(net261),
    .S0(net58),
    .S1(net275),
    .X(net562));
 sky130_fd_sc_hd__mux4_1 merge784 (.A0(net437),
    .A1(net431),
    .A2(net434),
    .A3(net328),
    .S0(net326),
    .S1(net329),
    .X(net563));
 sky130_fd_sc_hd__mux4_1 merge785 (.A0(net434),
    .A1(net342),
    .A2(net226),
    .A3(net707),
    .S0(net222),
    .S1(net577),
    .X(net564));
 sky130_fd_sc_hd__a41o_1 merge786 (.A1(net244),
    .A2(net359),
    .A3(net345),
    .A4(net241),
    .B1(net645),
    .X(net565));
 sky130_fd_sc_hd__mux4_1 merge787 (.A0(net163),
    .A1(net141),
    .A2(net154),
    .A3(net77),
    .S0(net783),
    .S1(net868),
    .X(net566));
 sky130_fd_sc_hd__mux4_1 merge788 (.A0(net146),
    .A1(net883),
    .A2(net254),
    .A3(net264),
    .S0(net877),
    .S1(net262),
    .X(net567));
 sky130_fd_sc_hd__mux4_1 merge789 (.A0(net221),
    .A1(net328),
    .A2(net330),
    .A3(net327),
    .S0(net814),
    .S1(net325),
    .X(net568));
 sky130_fd_sc_hd__mux4_1 merge790 (.A0(net431),
    .A1(net433),
    .A2(net437),
    .A3(net240),
    .S0(net254),
    .S1(net749),
    .X(net569));
 sky130_fd_sc_hd__xnor2_1 merge791 (.A(net295),
    .B(net301),
    .Y(net570));
 sky130_fd_sc_hd__dfrbp_1 merge792 (.CLK(clknet_4_12_0_clk),
    .D(net267),
    .Q(net272),
    .Q_N(net571));
 sky130_fd_sc_hd__dfrbp_1 merge793 (.CLK(clknet_4_1_0_clk),
    .D(net456),
    .RESET_B(net461),
    .Q(net574),
    .Q_N(net573));
 sky130_fd_sc_hd__dfrtn_1 merge794 (.CLK_N(clknet_4_5_0_clk),
    .D(net129),
    .RESET_B(net145),
    .Q(net575));
 sky130_fd_sc_hd__dfrtp_1 merge795 (.CLK(clknet_4_8_0_clk),
    .D(net402),
    .RESET_B(net404),
    .Q(net810));
 sky130_fd_sc_hd__dfrtp_1 merge796 (.CLK(clknet_4_4_0_clk),
    .D(net215),
    .RESET_B(net549),
    .Q(net576));
 sky130_fd_sc_hd__dfrtp_1 merge797 (.CLK(clknet_4_3_0_clk),
    .D(net478),
    .RESET_B(net481),
    .Q(net577));
 sky130_fd_sc_hd__dfsbp_1 merge798 (.CLK(clknet_4_12_0_clk),
    .D(net168),
    .SET_B(net152),
    .Q(net579),
    .Q_N(net578));
 sky130_fd_sc_hd__xnor2_1 merge799 (.A(net306),
    .B(net312),
    .Y(net580));
 sky130_fd_sc_hd__dfsbp_1 merge800 (.CLK(clknet_4_1_0_clk),
    .D(net550),
    .SET_B(net563),
    .Q(net582),
    .Q_N(net581));
 sky130_fd_sc_hd__xnor2_1 merge801 (.A(net85),
    .B(net554),
    .Y(net583));
 sky130_fd_sc_hd__xnor2_1 merge802 (.A(net529),
    .B(net538),
    .Y(net584));
 sky130_fd_sc_hd__xnor2_1 merge803 (.A(net100),
    .B(net89),
    .Y(net585));
 sky130_fd_sc_hd__xnor2_1 merge804 (.A(net414),
    .B(net415),
    .Y(net586));
 sky130_fd_sc_hd__xnor2_1 merge805 (.A(net365),
    .B(net366),
    .Y(net587));
 sky130_fd_sc_hd__xnor2_1 merge806 (.A(net66),
    .B(net65),
    .Y(net588));
 sky130_fd_sc_hd__dfstp_1 merge807 (.CLK(clknet_4_7_0_clk),
    .D(net256),
    .SET_B(net541),
    .Q(net589));
 sky130_fd_sc_hd__dfstp_1 merge808 (.CLK(clknet_4_14_0_clk),
    .D(net205),
    .SET_B(net208),
    .Q(net843));
 sky130_fd_sc_hd__dfstp_1 merge809 (.CLK(clknet_4_6_0_clk),
    .D(net385),
    .SET_B(net387),
    .Q(net590));
 sky130_fd_sc_hd__dlrbn_1 merge810 (.D(net193),
    .GATE_N(clknet_4_13_0_clk),
    .RESET_B(net170),
    .Q(net840),
    .Q_N(net591));
 sky130_fd_sc_hd__dlrbn_1 merge811 (.D(net546),
    .GATE_N(clknet_4_4_0_clk),
    .RESET_B(net568),
    .Q(net593),
    .Q_N(net592));
 sky130_fd_sc_hd__dlrbp_1 merge812 (.D(net503),
    .GATE(clknet_4_3_0_clk),
    .RESET_B(net505),
    .Q(net595),
    .Q_N(net594));
 sky130_fd_sc_hd__dlrbp_1 merge813 (.D(net520),
    .GATE(clknet_4_8_0_clk),
    .RESET_B(net539),
    .Q(net597),
    .Q_N(net596));
 sky130_fd_sc_hd__dlrtn_2 merge814 (.D(net570),
    .GATE_N(clknet_4_12_0_clk),
    .RESET_B(net560),
    .Q(net830));
 sky130_fd_sc_hd__dlrtn_1 merge815 (.D(net189),
    .GATE_N(clknet_4_15_0_clk),
    .RESET_B(net585),
    .Q(net598));
 sky130_fd_sc_hd__dlrtn_2 merge816 (.D(net138),
    .GATE_N(clknet_4_5_0_clk),
    .Q(net599));
 sky130_fd_sc_hd__dlrtp_1 merge817 (.GATE(clknet_4_13_0_clk),
    .RESET_B(net162),
    .Q(net190));
 sky130_fd_sc_hd__dlrtp_1 merge818 (.D(net388),
    .GATE(clknet_4_3_0_clk),
    .RESET_B(net427),
    .Q(net811));
 sky130_fd_sc_hd__xnor2_1 merge819 (.A(net547),
    .B(net556),
    .Y(net601));
 sky130_fd_sc_hd__dlrtp_1 merge820 (.D(net507),
    .GATE(clknet_4_8_0_clk),
    .RESET_B(net408),
    .Q(net602));
 sky130_fd_sc_hd__edfxbp_1 merge821 (.CLK(clknet_4_10_0_clk),
    .D(net315),
    .DE(net321),
    .Q(net827),
    .Q_N(net831));
 sky130_fd_sc_hd__edfxtp_1 merge822 (.CLK(clknet_4_13_0_clk),
    .D(net588),
    .DE(net68),
    .Q(net820));
 sky130_fd_sc_hd__xnor2_1 merge823 (.A(net423),
    .B(net418),
    .Y(net603));
 sky130_fd_sc_hd__sdlclkp_1 merge824 (.CLK(clknet_4_11_0_clk),
    .GATE(net580),
    .SCE(net316),
    .GCLK(net821));
 sky130_fd_sc_hd__sdlclkp_2 merge825 (.CLK(clknet_4_15_0_clk),
    .GATE(net74),
    .SCE(net93),
    .GCLK(net604));
 sky130_fd_sc_hd__sdlclkp_4 merge826 (.CLK(clknet_4_11_0_clk),
    .GATE(net369),
    .SCE(net561),
    .GCLK(net605));
 sky130_fd_sc_hd__dfrbp_2 merge827 (.CLK(clknet_4_13_0_clk),
    .D(net583),
    .RESET_B(net83),
    .Q(net859),
    .Q_N(net606));
 sky130_fd_sc_hd__dfrbp_1 merge828 (.CLK(clknet_4_12_0_clk),
    .D(net169),
    .RESET_B(net545),
    .Q(net608),
    .Q_N(net607));
 sky130_fd_sc_hd__xnor2_1 merge829 (.A(net95),
    .B(net99),
    .Y(net609));
 sky130_fd_sc_hd__dfrtn_1 merge830 (.CLK_N(clknet_4_14_0_clk),
    .D(net313),
    .RESET_B(net305),
    .Q(net610));
 sky130_fd_sc_hd__dfrtp_2 merge831 (.CLK(clknet_4_6_0_clk),
    .D(net562),
    .RESET_B(net587),
    .Q(net611));
 sky130_fd_sc_hd__dfrtp_1 merge832 (.CLK(clknet_4_0_0_clk),
    .D(net474),
    .RESET_B(net469),
    .Q(net612));
 sky130_fd_sc_hd__dfrtp_1 merge833 (.CLK(clknet_4_4_0_clk),
    .D(net565),
    .RESET_B(net553),
    .Q(net613));
 sky130_fd_sc_hd__xnor2_1 merge834 (.A(net462),
    .B(net525),
    .Y(net614));
 sky130_fd_sc_hd__dfsbp_1 merge835 (.CLK(clknet_4_10_0_clk),
    .D(net410),
    .SET_B(net421),
    .Q(net815),
    .Q_N(net615));
 sky130_fd_sc_hd__dfsbp_2 merge836 (.CLK(clknet_4_8_0_clk),
    .D(net406),
    .SET_B(net603),
    .Q(net616),
    .Q_N(net813));
 sky130_fd_sc_hd__dfstp_1 merge837 (.CLK(clknet_4_8_0_clk),
    .D(net523),
    .SET_B(net508),
    .Q(net617));
 sky130_fd_sc_hd__dfstp_1 merge838 (.CLK(clknet_4_8_0_clk),
    .D(net512),
    .SET_B(net514),
    .Q(net618));
 sky130_fd_sc_hd__dfstp_2 merge839 (.CLK(clknet_4_11_0_clk),
    .D(net292),
    .SET_B(net584),
    .Q(net823));
 sky130_fd_sc_hd__dlrbn_1 merge840 (.D(net559),
    .GATE_N(clknet_4_6_0_clk),
    .RESET_B(net567),
    .Q(net620),
    .Q_N(net619));
 sky130_fd_sc_hd__dlrbn_1 merge841 (.GATE_N(clknet_4_5_0_clk),
    .RESET_B(net223),
    .Q(net622),
    .Q_N(net621));
 sky130_fd_sc_hd__dlrbp_1 merge842 (.D(net457),
    .GATE(clknet_4_1_0_clk),
    .RESET_B(net564),
    .Q(net624),
    .Q_N(net623));
 sky130_fd_sc_hd__dlrbp_1 merge843 (.D(net542),
    .GATE(clknet_4_12_0_clk),
    .RESET_B(net172),
    .Q(net626),
    .Q_N(net625));
 sky130_fd_sc_hd__dlrtn_1 merge844 (.D(net308),
    .GATE_N(clknet_4_14_0_clk),
    .RESET_B(net310),
    .Q(net627));
 sky130_fd_sc_hd__dlrtn_1 merge845 (.D(net458),
    .GATE_N(clknet_4_0_0_clk),
    .RESET_B(net498),
    .Q(net628));
 sky130_fd_sc_hd__dlrtn_2 merge846 (.D(net601),
    .GATE_N(clknet_4_15_0_clk),
    .RESET_B(net609),
    .Q(net851));
 sky130_fd_sc_hd__dlrtp_2 merge847 (.D(net569),
    .GATE(clknet_4_1_0_clk),
    .RESET_B(net614),
    .Q(net629));
 sky130_fd_sc_hd__dlrtp_2 merge848 (.D(net566),
    .GATE(clknet_4_13_0_clk),
    .RESET_B(net202),
    .Q(net630));
 sky130_fd_sc_hd__dlrtp_1 merge849 (.D(net555),
    .GATE(clknet_4_11_0_clk),
    .RESET_B(net586),
    .Q(net631));
 sky130_fd_sc_hd__dfxbp_2 s850 (.CLK(clknet_4_13_0_clk),
    .D(net82),
    .Q(net856),
    .Q_N(net632));
 sky130_fd_sc_hd__dfxbp_2 s851 (.CLK(clknet_4_13_0_clk),
    .D(net165),
    .Q(net634),
    .Q_N(net633));
 sky130_fd_sc_hd__dfxtp_4 s852 (.CLK(clknet_4_12_0_clk),
    .D(net167),
    .Q(net635));
 sky130_fd_sc_hd__dfxtp_4 s853 (.CLK(clknet_4_12_0_clk),
    .D(net175),
    .Q(net817));
 sky130_fd_sc_hd__dfxtp_2 s854 (.CLK(clknet_4_14_0_clk),
    .D(net185),
    .Q(net636));
 sky130_fd_sc_hd__dlclkp_1 s855 (.CLK(clknet_4_15_0_clk),
    .GATE(net188),
    .GCLK(net852));
 sky130_fd_sc_hd__dlclkp_2 s856 (.CLK(clknet_4_14_0_clk),
    .GATE(net192),
    .GCLK(net637));
 sky130_fd_sc_hd__dlclkp_4 s857 (.CLK(clknet_4_15_0_clk),
    .GATE(net203),
    .GCLK(net638));
 sky130_fd_sc_hd__dlxbn_1 s858 (.D(net209),
    .GATE_N(clknet_4_14_0_clk),
    .Q(net640),
    .Q_N(net639));
 sky130_fd_sc_hd__dlxbn_1 s859 (.D(net210),
    .GATE_N(clknet_4_10_0_clk),
    .Q(net642),
    .Q_N(net641));
 sky130_fd_sc_hd__dlxbp_1 s860 (.D(net229),
    .GATE(clknet_4_4_0_clk),
    .Q(net644),
    .Q_N(net643));
 sky130_fd_sc_hd__dlxtn_1 s861 (.D(net255),
    .GATE_N(clknet_4_6_0_clk),
    .Q(net645));
 sky130_fd_sc_hd__dlxtn_4 s862 (.D(net263),
    .GATE_N(clknet_4_7_0_clk),
    .Q(net646));
 sky130_fd_sc_hd__dlxtn_1 s863 (.D(net274),
    .GATE_N(clknet_4_12_0_clk),
    .Q(net647));
 sky130_fd_sc_hd__dlxtp_1 s864 (.D(net276),
    .GATE(clknet_4_12_0_clk),
    .Q(net648));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s865 (.D(net279),
    .SLEEP_B(clknet_4_12_0_clk),
    .Q(net649));
 sky130_fd_sc_hd__dfxbp_2 s866 (.CLK(clknet_4_9_0_clk),
    .D(net294),
    .Q(net651),
    .Q_N(net650));
 sky130_fd_sc_hd__dfxbp_1 s867 (.CLK(clknet_4_11_0_clk),
    .D(net296),
    .Q(net832),
    .Q_N(net652));
 sky130_fd_sc_hd__dfxtp_1 s868 (.CLK(clknet_4_11_0_clk),
    .D(net297),
    .Q(net653));
 sky130_fd_sc_hd__dfxtp_1 s869 (.CLK(clknet_4_9_0_clk),
    .D(net298),
    .Q(net829));
 sky130_fd_sc_hd__dfxtp_1 s870 (.CLK(clknet_4_11_0_clk),
    .D(net302),
    .Q(net833));
 sky130_fd_sc_hd__dlclkp_1 s871 (.CLK(clknet_4_11_0_clk),
    .GATE(net307),
    .GCLK(net654));
 sky130_fd_sc_hd__dlclkp_2 s872 (.CLK(clknet_4_11_0_clk),
    .GATE(net309),
    .GCLK(net655));
 sky130_fd_sc_hd__dlclkp_4 s873 (.CLK(clknet_4_14_0_clk),
    .GATE(net311),
    .GCLK(net656));
 sky130_fd_sc_hd__dlxbn_1 s874 (.D(net333),
    .GATE_N(clknet_4_4_0_clk),
    .Q(net658),
    .Q_N(net657));
 sky130_fd_sc_hd__dlxbn_1 s875 (.D(net334),
    .GATE_N(clknet_4_1_0_clk),
    .Q(net660),
    .Q_N(net659));
 sky130_fd_sc_hd__dlxbp_1 s876 (.D(net337),
    .GATE(clknet_4_1_0_clk),
    .Q(net662),
    .Q_N(net661));
 sky130_fd_sc_hd__dlxtn_2 s877 (.D(net343),
    .GATE_N(clknet_4_1_0_clk),
    .Q(net663));
 sky130_fd_sc_hd__dlxtn_1 s878 (.D(net367),
    .GATE_N(clknet_4_6_0_clk),
    .Q(net664));
 sky130_fd_sc_hd__dlxtn_1 s879 (.D(net373),
    .GATE_N(clknet_4_9_0_clk),
    .Q(net665));
 sky130_fd_sc_hd__dlxtp_1 s880 (.D(net381),
    .GATE(clknet_4_6_0_clk),
    .Q(net666));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s881 (.D(net382),
    .SLEEP_B(clknet_4_6_0_clk),
    .Q(net667));
 sky130_fd_sc_hd__dfxbp_1 s882 (.CLK(clknet_4_6_0_clk),
    .D(net383),
    .Q(net669),
    .Q_N(net668));
 sky130_fd_sc_hd__dfxbp_1 s883 (.CLK(clknet_4_3_0_clk),
    .D(net384),
    .Q(net671),
    .Q_N(net670));
 sky130_fd_sc_hd__dfxtp_1 s884 (.CLK(clknet_4_10_0_clk),
    .D(net413),
    .Q(net672));
 sky130_fd_sc_hd__dfxtp_1 s885 (.CLK(clknet_4_10_0_clk),
    .D(net424),
    .Q(net673));
 sky130_fd_sc_hd__dfxtp_1 s886 (.CLK(clknet_4_10_0_clk),
    .D(net426),
    .Q(net674));
 sky130_fd_sc_hd__dlclkp_1 s887 (.CLK(clknet_4_10_0_clk),
    .GATE(net429),
    .GCLK(net675));
 sky130_fd_sc_hd__dlclkp_2 s888 (.CLK(clknet_4_0_0_clk),
    .GATE(net453),
    .GCLK(net676));
 sky130_fd_sc_hd__dlclkp_4 s889 (.CLK(clknet_4_0_0_clk),
    .GATE(net454),
    .GCLK(net677));
 sky130_fd_sc_hd__dlxbn_1 s890 (.D(net455),
    .GATE_N(clknet_4_0_0_clk),
    .Q(net679),
    .Q_N(net678));
 sky130_fd_sc_hd__dlxbn_1 s891 (.D(net464),
    .GATE_N(clknet_4_0_0_clk),
    .Q(net681),
    .Q_N(net680));
 sky130_fd_sc_hd__dlxbp_1 s892 (.D(net475),
    .GATE(clknet_4_0_0_clk),
    .Q(net683),
    .Q_N(net682));
 sky130_fd_sc_hd__dlxtn_1 s893 (.D(net476),
    .GATE_N(clknet_4_2_0_clk),
    .Q(net684));
 sky130_fd_sc_hd__dlxtn_2 s894 (.D(net477),
    .GATE_N(clknet_4_2_0_clk),
    .Q(net685));
 sky130_fd_sc_hd__dlxtn_1 s895 (.D(net486),
    .GATE_N(clknet_4_3_0_clk),
    .Q(net686));
 sky130_fd_sc_hd__dlxtp_1 s896 (.D(net487),
    .GATE(clknet_4_2_0_clk),
    .Q(net687));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s897 (.D(net490),
    .SLEEP_B(clknet_4_3_0_clk),
    .Q(net688));
 sky130_fd_sc_hd__dfxbp_1 s898 (.CLK(clknet_4_3_0_clk),
    .D(net491),
    .Q(net690),
    .Q_N(net689));
 sky130_fd_sc_hd__dfxbp_1 s899 (.CLK(clknet_4_2_0_clk),
    .D(net492),
    .Q(net692),
    .Q_N(net691));
 sky130_fd_sc_hd__dfxtp_1 s900 (.CLK(clknet_4_2_0_clk),
    .D(net493),
    .Q(net693));
 sky130_fd_sc_hd__dfxtp_1 s901 (.CLK(clknet_4_2_0_clk),
    .D(net496),
    .Q(net694));
 sky130_fd_sc_hd__dfxtp_2 s902 (.CLK(clknet_4_2_0_clk),
    .D(net497),
    .Q(net695));
 sky130_fd_sc_hd__dlclkp_1 s903 (.CLK(clknet_4_2_0_clk),
    .GATE(net501),
    .GCLK(net696));
 sky130_fd_sc_hd__dlclkp_2 s904 (.CLK(clknet_4_8_0_clk),
    .GATE(net528),
    .GCLK(net697));
 sky130_fd_sc_hd__dlclkp_4 s905 (.CLK(clknet_4_10_0_clk),
    .GATE(net532),
    .GCLK(net698));
 sky130_fd_sc_hd__dlxbn_1 s906 (.D(net534),
    .GATE_N(clknet_4_8_0_clk),
    .Q(net700),
    .Q_N(net699));
 sky130_fd_sc_hd__dlxbn_1 s907 (.D(net543),
    .GATE_N(clknet_4_9_0_clk),
    .Q(net702),
    .Q_N(net701));
 sky130_fd_sc_hd__dlxbp_1 s908 (.D(net544),
    .GATE(clknet_4_14_0_clk),
    .Q(net704),
    .Q_N(net703));
 sky130_fd_sc_hd__dlxtn_1 s909 (.D(net548),
    .GATE_N(clknet_4_9_0_clk),
    .Q(net705));
 sky130_fd_sc_hd__dlxtn_1 s910 (.D(net558),
    .GATE_N(clknet_4_9_0_clk),
    .Q(net706));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Right_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Right_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Right_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Right_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Right_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Right_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Right_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Right_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Right_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Right_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Right_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Right_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Right_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Right_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Right_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Right_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Right_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Right_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Right_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Right_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Right_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_161 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_162 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_163 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_164 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_165 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_166 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_167 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_168 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_169 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_170 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_171 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_172 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_173 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_174 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_175 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_176 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_177 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_178 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_179 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_180 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_181 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_182 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Left_183 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Left_184 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Left_185 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Left_186 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Left_187 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Left_188 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Left_189 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Left_190 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Left_191 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Left_192 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Left_193 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Left_194 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Left_195 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Left_196 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Left_197 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Left_198 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Left_199 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Left_200 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Left_201 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Left_202 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Left_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1347 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(in0),
    .X(net144));
 sky130_fd_sc_hd__buf_2 input2 (.A(in1),
    .X(net557));
 sky130_fd_sc_hd__buf_6 input3 (.A(in10),
    .X(net707));
 sky130_fd_sc_hd__buf_2 input4 (.A(in11),
    .X(net708));
 sky130_fd_sc_hd__dlymetal6s2s_1 input5 (.A(in12),
    .X(net709));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(in13),
    .X(net710));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(in14),
    .X(net711));
 sky130_fd_sc_hd__clkbuf_2 input8 (.A(in15),
    .X(net712));
 sky130_fd_sc_hd__clkbuf_2 input9 (.A(in16),
    .X(net713));
 sky130_fd_sc_hd__buf_1 input10 (.A(in17),
    .X(net714));
 sky130_fd_sc_hd__clkbuf_8 input11 (.A(in18),
    .X(net715));
 sky130_fd_sc_hd__buf_1 input12 (.A(in19),
    .X(net716));
 sky130_fd_sc_hd__buf_2 input13 (.A(in2),
    .X(net717));
 sky130_fd_sc_hd__buf_1 input14 (.A(in20),
    .X(net718));
 sky130_fd_sc_hd__buf_2 input15 (.A(in21),
    .X(net719));
 sky130_fd_sc_hd__buf_1 input16 (.A(in22),
    .X(net720));
 sky130_fd_sc_hd__buf_4 input17 (.A(in23),
    .X(net721));
 sky130_fd_sc_hd__buf_1 input18 (.A(in24),
    .X(net722));
 sky130_fd_sc_hd__clkbuf_2 input19 (.A(in25),
    .X(net723));
 sky130_fd_sc_hd__clkbuf_2 input20 (.A(in26),
    .X(net724));
 sky130_fd_sc_hd__buf_2 input21 (.A(in27),
    .X(net725));
 sky130_fd_sc_hd__buf_4 input22 (.A(in28),
    .X(net726));
 sky130_fd_sc_hd__buf_1 input23 (.A(in29),
    .X(net727));
 sky130_fd_sc_hd__buf_2 input24 (.A(in3),
    .X(net728));
 sky130_fd_sc_hd__buf_1 input25 (.A(in30),
    .X(net729));
 sky130_fd_sc_hd__buf_1 input26 (.A(in31),
    .X(net730));
 sky130_fd_sc_hd__dlymetal6s2s_1 input27 (.A(in32),
    .X(net731));
 sky130_fd_sc_hd__buf_1 input28 (.A(in33),
    .X(net732));
 sky130_fd_sc_hd__clkbuf_1 input29 (.A(in34),
    .X(net733));
 sky130_fd_sc_hd__clkbuf_1 input30 (.A(in35),
    .X(net734));
 sky130_fd_sc_hd__buf_1 input31 (.A(in36),
    .X(net735));
 sky130_fd_sc_hd__dlymetal6s2s_1 input32 (.A(in37),
    .X(net736));
 sky130_fd_sc_hd__buf_1 input33 (.A(in38),
    .X(net737));
 sky130_fd_sc_hd__clkbuf_2 input34 (.A(in39),
    .X(net738));
 sky130_fd_sc_hd__buf_1 input35 (.A(in4),
    .X(net739));
 sky130_fd_sc_hd__clkbuf_2 input36 (.A(in40),
    .X(net740));
 sky130_fd_sc_hd__buf_1 input37 (.A(in41),
    .X(net741));
 sky130_fd_sc_hd__buf_1 input38 (.A(in42),
    .X(net742));
 sky130_fd_sc_hd__buf_1 input39 (.A(in43),
    .X(net743));
 sky130_fd_sc_hd__buf_2 input40 (.A(in44),
    .X(net744));
 sky130_fd_sc_hd__clkbuf_2 input41 (.A(in45),
    .X(net745));
 sky130_fd_sc_hd__clkbuf_1 input42 (.A(in46),
    .X(net746));
 sky130_fd_sc_hd__clkbuf_2 input43 (.A(in47),
    .X(net747));
 sky130_fd_sc_hd__clkbuf_1 input44 (.A(in48),
    .X(net748));
 sky130_fd_sc_hd__clkbuf_4 input45 (.A(in49),
    .X(net749));
 sky130_fd_sc_hd__buf_12 input46 (.A(in5),
    .X(net750));
 sky130_fd_sc_hd__clkbuf_2 input47 (.A(in50),
    .X(net751));
 sky130_fd_sc_hd__buf_2 input48 (.A(in51),
    .X(net752));
 sky130_fd_sc_hd__clkbuf_1 input49 (.A(in52),
    .X(net753));
 sky130_fd_sc_hd__clkbuf_1 input50 (.A(in54),
    .X(net754));
 sky130_fd_sc_hd__buf_1 input51 (.A(in55),
    .X(net755));
 sky130_fd_sc_hd__clkbuf_2 input52 (.A(in56),
    .X(net756));
 sky130_fd_sc_hd__buf_1 input53 (.A(in57),
    .X(net757));
 sky130_fd_sc_hd__clkbuf_2 input54 (.A(in58),
    .X(net758));
 sky130_fd_sc_hd__buf_1 input55 (.A(in59),
    .X(net759));
 sky130_fd_sc_hd__clkbuf_2 input56 (.A(in6),
    .X(net760));
 sky130_fd_sc_hd__clkbuf_2 input57 (.A(in60),
    .X(net761));
 sky130_fd_sc_hd__clkbuf_2 input58 (.A(in61),
    .X(net762));
 sky130_fd_sc_hd__clkbuf_2 input59 (.A(in62),
    .X(net763));
 sky130_fd_sc_hd__clkbuf_2 input60 (.A(in63),
    .X(net764));
 sky130_fd_sc_hd__buf_1 input61 (.A(in65),
    .X(net765));
 sky130_fd_sc_hd__dlymetal6s2s_1 input62 (.A(in66),
    .X(net766));
 sky130_fd_sc_hd__buf_1 input63 (.A(in67),
    .X(net767));
 sky130_fd_sc_hd__buf_1 input64 (.A(in68),
    .X(net768));
 sky130_fd_sc_hd__buf_1 input65 (.A(in69),
    .X(net769));
 sky130_fd_sc_hd__buf_4 input66 (.A(in7),
    .X(net770));
 sky130_fd_sc_hd__clkbuf_2 input67 (.A(in70),
    .X(net771));
 sky130_fd_sc_hd__clkbuf_1 input68 (.A(in71),
    .X(net772));
 sky130_fd_sc_hd__clkbuf_4 input69 (.A(in72),
    .X(net773));
 sky130_fd_sc_hd__clkbuf_1 input70 (.A(in73),
    .X(net774));
 sky130_fd_sc_hd__clkbuf_1 input71 (.A(in74),
    .X(net775));
 sky130_fd_sc_hd__buf_1 input72 (.A(in75),
    .X(net776));
 sky130_fd_sc_hd__clkbuf_1 input73 (.A(in76),
    .X(net777));
 sky130_fd_sc_hd__clkbuf_1 input74 (.A(in77),
    .X(net778));
 sky130_fd_sc_hd__clkbuf_1 input75 (.A(in78),
    .X(net779));
 sky130_fd_sc_hd__clkbuf_1 input76 (.A(in79),
    .X(net780));
 sky130_fd_sc_hd__clkbuf_1 input77 (.A(in8),
    .X(net781));
 sky130_fd_sc_hd__buf_1 input78 (.A(in80),
    .X(net782));
 sky130_fd_sc_hd__clkbuf_1 input79 (.A(in81),
    .X(net783));
 sky130_fd_sc_hd__clkbuf_2 input80 (.A(in82),
    .X(net784));
 sky130_fd_sc_hd__buf_1 input81 (.A(in83),
    .X(net785));
 sky130_fd_sc_hd__clkbuf_1 input82 (.A(in84),
    .X(net786));
 sky130_fd_sc_hd__clkbuf_4 input83 (.A(in85),
    .X(net787));
 sky130_fd_sc_hd__clkbuf_2 input84 (.A(in86),
    .X(net788));
 sky130_fd_sc_hd__buf_1 input85 (.A(in87),
    .X(net789));
 sky130_fd_sc_hd__clkbuf_1 input86 (.A(in88),
    .X(net790));
 sky130_fd_sc_hd__dlymetal6s2s_1 input87 (.A(in89),
    .X(net791));
 sky130_fd_sc_hd__clkbuf_4 input88 (.A(in9),
    .X(net792));
 sky130_fd_sc_hd__clkbuf_1 input89 (.A(in90),
    .X(net793));
 sky130_fd_sc_hd__clkbuf_1 input90 (.A(in91),
    .X(net794));
 sky130_fd_sc_hd__clkbuf_1 input91 (.A(in92),
    .X(net795));
 sky130_fd_sc_hd__buf_2 input92 (.A(in93),
    .X(net796));
 sky130_fd_sc_hd__clkbuf_2 input93 (.A(in94),
    .X(net797));
 sky130_fd_sc_hd__buf_1 input94 (.A(in95),
    .X(net798));
 sky130_fd_sc_hd__clkbuf_1 input95 (.A(in96),
    .X(net799));
 sky130_fd_sc_hd__clkbuf_1 input96 (.A(in97),
    .X(net800));
 sky130_fd_sc_hd__buf_2 input97 (.A(in98),
    .X(net801));
 sky130_fd_sc_hd__buf_1 input98 (.A(in99),
    .X(net802));
 sky130_fd_sc_hd__buf_2 output99 (.A(net803),
    .X(out0));
 sky130_fd_sc_hd__buf_2 output100 (.A(net804),
    .X(out1));
 sky130_fd_sc_hd__buf_2 output101 (.A(net805),
    .X(out10));
 sky130_fd_sc_hd__clkbuf_1 output102 (.A(net806),
    .X(out11));
 sky130_fd_sc_hd__clkbuf_1 output103 (.A(net807),
    .X(out12));
 sky130_fd_sc_hd__clkbuf_4 output104 (.A(net808),
    .X(out13));
 sky130_fd_sc_hd__clkbuf_1 output105 (.A(clknet_1_1__leaf_net809),
    .X(out14));
 sky130_fd_sc_hd__buf_2 output106 (.A(net810),
    .X(out15));
 sky130_fd_sc_hd__buf_2 output107 (.A(net811),
    .X(out16));
 sky130_fd_sc_hd__clkbuf_1 output108 (.A(clknet_1_0__leaf_net812),
    .X(out17));
 sky130_fd_sc_hd__buf_2 output109 (.A(net813),
    .X(out19));
 sky130_fd_sc_hd__buf_2 output110 (.A(net814),
    .X(out2));
 sky130_fd_sc_hd__buf_2 output111 (.A(net815),
    .X(out21));
 sky130_fd_sc_hd__clkbuf_1 output112 (.A(clknet_1_1__leaf_net816),
    .X(out22));
 sky130_fd_sc_hd__buf_2 output113 (.A(net817),
    .X(out23));
 sky130_fd_sc_hd__buf_2 output114 (.A(net818),
    .X(out24));
 sky130_fd_sc_hd__buf_2 output115 (.A(net819),
    .X(out25));
 sky130_fd_sc_hd__clkbuf_4 output116 (.A(net897),
    .X(out26));
 sky130_fd_sc_hd__clkbuf_1 output117 (.A(clknet_1_1__leaf_net821),
    .X(out27));
 sky130_fd_sc_hd__buf_2 output118 (.A(net822),
    .X(out28));
 sky130_fd_sc_hd__buf_2 output119 (.A(net823),
    .X(out29));
 sky130_fd_sc_hd__clkbuf_1 output120 (.A(clknet_1_0__leaf_net824),
    .X(out3));
 sky130_fd_sc_hd__clkbuf_1 output121 (.A(net825),
    .X(out30));
 sky130_fd_sc_hd__buf_2 output122 (.A(net826),
    .X(out31));
 sky130_fd_sc_hd__buf_2 output123 (.A(net827),
    .X(out32));
 sky130_fd_sc_hd__buf_2 output124 (.A(net828),
    .X(out33));
 sky130_fd_sc_hd__buf_2 output125 (.A(net829),
    .X(out35));
 sky130_fd_sc_hd__clkbuf_4 output126 (.A(net830),
    .X(out36));
 sky130_fd_sc_hd__buf_2 output127 (.A(net831),
    .X(out38));
 sky130_fd_sc_hd__buf_2 output128 (.A(net832),
    .X(out40));
 sky130_fd_sc_hd__buf_2 output129 (.A(net833),
    .X(out41));
 sky130_fd_sc_hd__buf_2 output130 (.A(net834),
    .X(out42));
 sky130_fd_sc_hd__clkbuf_4 output131 (.A(net835),
    .X(out44));
 sky130_fd_sc_hd__clkbuf_1 output132 (.A(clknet_1_1__leaf_net836),
    .X(out45));
 sky130_fd_sc_hd__clkbuf_4 output133 (.A(net837),
    .X(out47));
 sky130_fd_sc_hd__clkbuf_1 output134 (.A(clknet_1_1__leaf_net838),
    .X(out48));
 sky130_fd_sc_hd__buf_2 output135 (.A(net839),
    .X(out5));
 sky130_fd_sc_hd__clkbuf_4 output136 (.A(net840),
    .X(out50));
 sky130_fd_sc_hd__clkbuf_1 output137 (.A(clknet_1_1__leaf_net841),
    .X(out51));
 sky130_fd_sc_hd__clkbuf_4 output138 (.A(net842),
    .X(out52));
 sky130_fd_sc_hd__buf_2 output139 (.A(net843),
    .X(out53));
 sky130_fd_sc_hd__clkbuf_4 output140 (.A(net844),
    .X(out55));
 sky130_fd_sc_hd__buf_2 output141 (.A(net845),
    .X(out56));
 sky130_fd_sc_hd__clkbuf_4 output142 (.A(net846),
    .X(out57));
 sky130_fd_sc_hd__clkbuf_4 output143 (.A(net885),
    .X(out58));
 sky130_fd_sc_hd__buf_2 output144 (.A(net848),
    .X(out6));
 sky130_fd_sc_hd__clkbuf_4 output145 (.A(net849),
    .X(out60));
 sky130_fd_sc_hd__clkbuf_4 output146 (.A(net850),
    .X(out63));
 sky130_fd_sc_hd__buf_2 output147 (.A(net851),
    .X(out64));
 sky130_fd_sc_hd__clkbuf_1 output148 (.A(clknet_1_1__leaf_net852),
    .X(out65));
 sky130_fd_sc_hd__clkbuf_4 output149 (.A(net853),
    .X(out68));
 sky130_fd_sc_hd__clkbuf_4 output150 (.A(net854),
    .X(out69));
 sky130_fd_sc_hd__clkbuf_1 output151 (.A(clknet_1_1__leaf_net855),
    .X(out7));
 sky130_fd_sc_hd__buf_2 output152 (.A(net856),
    .X(out70));
 sky130_fd_sc_hd__clkbuf_4 output153 (.A(net857),
    .X(out71));
 sky130_fd_sc_hd__clkbuf_4 output154 (.A(net858),
    .X(out73));
 sky130_fd_sc_hd__buf_2 output155 (.A(net859),
    .X(out75));
 sky130_fd_sc_hd__buf_2 output156 (.A(net860),
    .X(out76));
 sky130_fd_sc_hd__buf_2 output157 (.A(net861),
    .X(out78));
 sky130_fd_sc_hd__clkbuf_1 output158 (.A(clknet_1_1__leaf_net862),
    .X(out79));
 sky130_fd_sc_hd__buf_2 output159 (.A(net904),
    .X(out8));
 sky130_fd_sc_hd__buf_2 output160 (.A(net864),
    .X(out80));
 sky130_fd_sc_hd__buf_2 output161 (.A(net865),
    .X(out82));
 sky130_fd_sc_hd__buf_2 output162 (.A(net866),
    .X(out84));
 sky130_fd_sc_hd__buf_2 output163 (.A(net867),
    .X(out85));
 sky130_fd_sc_hd__buf_2 output164 (.A(net868),
    .X(out87));
 sky130_fd_sc_hd__buf_2 output165 (.A(net869),
    .X(out88));
 sky130_fd_sc_hd__buf_2 output166 (.A(net870),
    .X(out89));
 sky130_fd_sc_hd__buf_2 output167 (.A(net924),
    .X(out9));
 sky130_fd_sc_hd__buf_2 output168 (.A(net872),
    .X(out90));
 sky130_fd_sc_hd__buf_2 output169 (.A(net873),
    .X(out93));
 sky130_fd_sc_hd__buf_2 output170 (.A(net874),
    .X(out98));
 sky130_fd_sc_hd__buf_2 output171 (.A(net875),
    .X(out99));
 sky130_fd_sc_hd__clkbuf_4 fanout172 (.A(net234),
    .X(net876));
 sky130_fd_sc_hd__clkbuf_4 fanout173 (.A(net155),
    .X(net877));
 sky130_fd_sc_hd__buf_4 max_cap174 (.A(net214),
    .X(net878));
 sky130_fd_sc_hd__buf_8 fanout175 (.A(net131),
    .X(net879));
 sky130_fd_sc_hd__clkbuf_4 fanout176 (.A(net269),
    .X(net880));
 sky130_fd_sc_hd__buf_2 fanout177 (.A(net822),
    .X(net881));
 sky130_fd_sc_hd__buf_4 fanout178 (.A(net126),
    .X(net882));
 sky130_fd_sc_hd__buf_4 fanout179 (.A(net116),
    .X(net883));
 sky130_fd_sc_hd__buf_4 fanout180 (.A(net110),
    .X(net884));
 sky130_fd_sc_hd__clkbuf_4 fanout181 (.A(net847),
    .X(net885));
 sky130_fd_sc_hd__buf_4 max_cap182 (.A(net115),
    .X(net886));
 sky130_fd_sc_hd__buf_8 fanout183 (.A(net889),
    .X(net887));
 sky130_fd_sc_hd__clkbuf_2 fanout184 (.A(net889),
    .X(net888));
 sky130_fd_sc_hd__buf_8 fanout185 (.A(net44),
    .X(net889));
 sky130_fd_sc_hd__buf_4 max_cap186 (.A(net106),
    .X(net890));
 sky130_fd_sc_hd__buf_4 fanout187 (.A(net338),
    .X(net891));
 sky130_fd_sc_hd__buf_12 fanout188 (.A(net871),
    .X(net892));
 sky130_fd_sc_hd__clkbuf_4 fanout189 (.A(net895),
    .X(net893));
 sky130_fd_sc_hd__buf_2 fanout190 (.A(net895),
    .X(net894));
 sky130_fd_sc_hd__buf_2 fanout191 (.A(net665),
    .X(net895));
 sky130_fd_sc_hd__clkbuf_4 fanout192 (.A(net820),
    .X(net896));
 sky130_fd_sc_hd__buf_2 fanout193 (.A(net820),
    .X(net897));
 sky130_fd_sc_hd__buf_2 fanout194 (.A(net899),
    .X(net898));
 sky130_fd_sc_hd__clkbuf_2 fanout195 (.A(net50),
    .X(net899));
 sky130_fd_sc_hd__buf_2 fanout196 (.A(net50),
    .X(net900));
 sky130_fd_sc_hd__buf_8 fanout197 (.A(net902),
    .X(net901));
 sky130_fd_sc_hd__buf_8 fanout198 (.A(net903),
    .X(net902));
 sky130_fd_sc_hd__buf_8 fanout199 (.A(net904),
    .X(net903));
 sky130_fd_sc_hd__buf_12 fanout200 (.A(net863),
    .X(net904));
 sky130_fd_sc_hd__buf_4 fanout201 (.A(net906),
    .X(net905));
 sky130_fd_sc_hd__buf_4 fanout202 (.A(net907),
    .X(net906));
 sky130_fd_sc_hd__clkbuf_4 fanout203 (.A(net711),
    .X(net907));
 sky130_fd_sc_hd__clkbuf_8 fanout204 (.A(net730),
    .X(net908));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net698 (.A(net698),
    .X(clknet_0_net698));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net698 (.A(clknet_0_net698),
    .X(clknet_1_0__leaf_net698));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net698 (.A(clknet_0_net698),
    .X(clknet_1_1__leaf_net698));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net697 (.A(net697),
    .X(clknet_0_net697));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net697 (.A(clknet_0_net697),
    .X(clknet_1_0__leaf_net697));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net697 (.A(clknet_0_net697),
    .X(clknet_1_1__leaf_net697));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net696 (.A(net696),
    .X(clknet_0_net696));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net696 (.A(clknet_0_net696),
    .X(clknet_1_0__leaf_net696));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net696 (.A(clknet_0_net696),
    .X(clknet_1_1__leaf_net696));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net521 (.A(net521),
    .X(clknet_0_net521));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net521 (.A(clknet_0_net521),
    .X(clknet_1_0__leaf_net521));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net521 (.A(clknet_0_net521),
    .X(clknet_1_1__leaf_net521));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net522 (.A(net522),
    .X(clknet_0_net522));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net522 (.A(clknet_0_net522),
    .X(clknet_1_0__leaf_net522));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net522 (.A(clknet_0_net522),
    .X(clknet_1_1__leaf_net522));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net526 (.A(net526),
    .X(clknet_0_net526));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net526 (.A(clknet_0_net526),
    .X(clknet_1_0__leaf_net526));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net526 (.A(clknet_0_net526),
    .X(clknet_1_1__leaf_net526));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net502 (.A(net502),
    .X(clknet_0_net502));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net502 (.A(clknet_0_net502),
    .X(clknet_1_0__leaf_net502));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net502 (.A(clknet_0_net502),
    .X(clknet_1_1__leaf_net502));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net677 (.A(net677),
    .X(clknet_0_net677));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net677 (.A(clknet_0_net677),
    .X(clknet_1_0__leaf_net677));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net677 (.A(clknet_0_net677),
    .X(clknet_1_1__leaf_net677));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net463 (.A(net463),
    .X(clknet_0_net463));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net463 (.A(clknet_0_net463),
    .X(clknet_1_0__leaf_net463));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net463 (.A(clknet_0_net463),
    .X(clknet_1_1__leaf_net463));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net482 (.A(net482),
    .X(clknet_0_net482));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net482 (.A(clknet_0_net482),
    .X(clknet_1_0__leaf_net482));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net482 (.A(clknet_0_net482),
    .X(clknet_1_1__leaf_net482));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net488 (.A(net488),
    .X(clknet_0_net488));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net488 (.A(clknet_0_net488),
    .X(clknet_1_0__leaf_net488));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net488 (.A(clknet_0_net488),
    .X(clknet_1_1__leaf_net488));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net676 (.A(net676),
    .X(clknet_0_net676));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net676 (.A(clknet_0_net676),
    .X(clknet_1_0__leaf_net676));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net676 (.A(clknet_0_net676),
    .X(clknet_1_1__leaf_net676));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net459 (.A(net459),
    .X(clknet_0_net459));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net459 (.A(clknet_0_net459),
    .X(clknet_1_0__leaf_net459));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net459 (.A(clknet_0_net459),
    .X(clknet_1_1__leaf_net459));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net466 (.A(net466),
    .X(clknet_0_net466));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net466 (.A(clknet_0_net466),
    .X(clknet_1_0__leaf_net466));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net466 (.A(clknet_0_net466),
    .X(clknet_1_1__leaf_net466));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net473 (.A(net473),
    .X(clknet_0_net473));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net473 (.A(clknet_0_net473),
    .X(clknet_1_0__leaf_net473));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net473 (.A(clknet_0_net473),
    .X(clknet_1_1__leaf_net473));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net675 (.A(net675),
    .X(clknet_0_net675));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net675 (.A(clknet_0_net675),
    .X(clknet_1_0__leaf_net675));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net675 (.A(clknet_0_net675),
    .X(clknet_1_1__leaf_net675));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net656 (.A(net656),
    .X(clknet_0_net656));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net656 (.A(clknet_0_net656),
    .X(clknet_1_0__leaf_net656));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net656 (.A(clknet_0_net656),
    .X(clknet_1_1__leaf_net656));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net314 (.A(net314),
    .X(clknet_0_net314));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net314 (.A(clknet_0_net314),
    .X(clknet_1_0__leaf_net314));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net314 (.A(clknet_0_net314),
    .X(clknet_1_1__leaf_net314));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net655 (.A(net655),
    .X(clknet_0_net655));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net655 (.A(clknet_0_net655),
    .X(clknet_1_0__leaf_net655));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net655 (.A(clknet_0_net655),
    .X(clknet_1_1__leaf_net655));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net420 (.A(net420),
    .X(clknet_0_net420));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net420 (.A(clknet_0_net420),
    .X(clknet_1_0__leaf_net420));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net420 (.A(clknet_0_net420),
    .X(clknet_1_1__leaf_net420));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net412 (.A(net412),
    .X(clknet_0_net412));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net412 (.A(clknet_0_net412),
    .X(clknet_1_0__leaf_net412));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net412 (.A(clknet_0_net412),
    .X(clknet_1_1__leaf_net412));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net809 (.A(net809),
    .X(clknet_0_net809));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net809 (.A(clknet_0_net809),
    .X(clknet_1_0__leaf_net809));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net809 (.A(clknet_0_net809),
    .X(clknet_1_1__leaf_net809));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net855 (.A(net855),
    .X(clknet_0_net855));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net855 (.A(clknet_0_net855),
    .X(clknet_1_0__leaf_net855));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net855 (.A(clknet_0_net855),
    .X(clknet_1_1__leaf_net855));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net317 (.A(net317),
    .X(clknet_0_net317));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net317 (.A(clknet_0_net317),
    .X(clknet_1_0__leaf_net317));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net317 (.A(clknet_0_net317),
    .X(clknet_1_1__leaf_net317));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net318 (.A(net318),
    .X(clknet_0_net318));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net318 (.A(clknet_0_net318),
    .X(clknet_1_0__leaf_net318));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net318 (.A(clknet_0_net318),
    .X(clknet_1_1__leaf_net318));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net654 (.A(net654),
    .X(clknet_0_net654));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net654 (.A(clknet_0_net654),
    .X(clknet_1_0__leaf_net654));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net654 (.A(clknet_0_net654),
    .X(clknet_1_1__leaf_net654));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net821 (.A(net821),
    .X(clknet_0_net821));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net821 (.A(clknet_0_net821),
    .X(clknet_1_0__leaf_net821));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net821 (.A(clknet_0_net821),
    .X(clknet_1_1__leaf_net821));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net638 (.A(net638),
    .X(clknet_0_net638));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net638 (.A(clknet_0_net638),
    .X(clknet_1_0__leaf_net638));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net638 (.A(clknet_0_net638),
    .X(clknet_1_1__leaf_net638));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net207 (.A(net207),
    .X(clknet_0_net207));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net207 (.A(clknet_0_net207),
    .X(clknet_1_0__leaf_net207));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net207 (.A(clknet_0_net207),
    .X(clknet_1_1__leaf_net207));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net824 (.A(net824),
    .X(clknet_0_net824));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net824 (.A(clknet_0_net824),
    .X(clknet_1_0__leaf_net824));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net824 (.A(clknet_0_net824),
    .X(clknet_1_1__leaf_net824));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net204 (.A(net204),
    .X(clknet_0_net204));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net204 (.A(clknet_0_net204),
    .X(clknet_1_0__leaf_net204));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net204 (.A(clknet_0_net204),
    .X(clknet_1_1__leaf_net204));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net816 (.A(net816),
    .X(clknet_0_net816));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net816 (.A(clknet_0_net816),
    .X(clknet_1_0__leaf_net816));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net816 (.A(clknet_0_net816),
    .X(clknet_1_1__leaf_net816));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net812 (.A(net812),
    .X(clknet_0_net812));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net812 (.A(clknet_0_net812),
    .X(clknet_1_0__leaf_net812));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net812 (.A(clknet_0_net812),
    .X(clknet_1_1__leaf_net812));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net637 (.A(net637),
    .X(clknet_0_net637));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net637 (.A(clknet_0_net637),
    .X(clknet_1_0__leaf_net637));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net637 (.A(clknet_0_net637),
    .X(clknet_1_1__leaf_net637));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net289 (.A(net289),
    .X(clknet_0_net289));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net289 (.A(clknet_0_net289),
    .X(clknet_1_0__leaf_net289));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net289 (.A(clknet_0_net289),
    .X(clknet_1_1__leaf_net289));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net285 (.A(net285),
    .X(clknet_0_net285));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net285 (.A(clknet_0_net285),
    .X(clknet_1_0__leaf_net285));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net285 (.A(clknet_0_net285),
    .X(clknet_1_1__leaf_net285));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net401 (.A(net401),
    .X(clknet_0_net401));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net401 (.A(clknet_0_net401),
    .X(clknet_1_0__leaf_net401));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net401 (.A(clknet_0_net401),
    .X(clknet_1_1__leaf_net401));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net504 (.A(net504),
    .X(clknet_0_net504));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net504 (.A(clknet_0_net504),
    .X(clknet_1_0__leaf_net504));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net504 (.A(clknet_0_net504),
    .X(clknet_1_1__leaf_net504));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net511 (.A(net511),
    .X(clknet_0_net511));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net511 (.A(clknet_0_net511),
    .X(clknet_1_0__leaf_net511));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net511 (.A(clknet_0_net511),
    .X(clknet_1_1__leaf_net511));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net396 (.A(net396),
    .X(clknet_0_net396));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net396 (.A(clknet_0_net396),
    .X(clknet_1_0__leaf_net396));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net396 (.A(clknet_0_net396),
    .X(clknet_1_1__leaf_net396));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net605 (.A(net605),
    .X(clknet_0_net605));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net605 (.A(clknet_0_net605),
    .X(clknet_1_0__leaf_net605));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net605 (.A(clknet_0_net605),
    .X(clknet_1_1__leaf_net605));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net398 (.A(net398),
    .X(clknet_0_net398));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net398 (.A(clknet_0_net398),
    .X(clknet_1_0__leaf_net398));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net398 (.A(clknet_0_net398),
    .X(clknet_1_1__leaf_net398));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net380 (.A(net380),
    .X(clknet_0_net380));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net380 (.A(clknet_0_net380),
    .X(clknet_1_0__leaf_net380));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net380 (.A(clknet_0_net380),
    .X(clknet_1_1__leaf_net380));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net392 (.A(net392),
    .X(clknet_0_net392));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net392 (.A(clknet_0_net392),
    .X(clknet_1_0__leaf_net392));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net392 (.A(clknet_0_net392),
    .X(clknet_1_1__leaf_net392));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net282 (.A(net282),
    .X(clknet_0_net282));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net282 (.A(clknet_0_net282),
    .X(clknet_1_0__leaf_net282));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net282 (.A(clknet_0_net282),
    .X(clknet_1_1__leaf_net282));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net286 (.A(net286),
    .X(clknet_0_net286));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net286 (.A(clknet_0_net286),
    .X(clknet_1_0__leaf_net286));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net286 (.A(clknet_0_net286),
    .X(clknet_1_1__leaf_net286));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net290 (.A(net290),
    .X(clknet_0_net290));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net290 (.A(clknet_0_net290),
    .X(clknet_1_0__leaf_net290));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net290 (.A(clknet_0_net290),
    .X(clknet_1_1__leaf_net290));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net291 (.A(net291),
    .X(clknet_0_net291));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net291 (.A(clknet_0_net291),
    .X(clknet_1_0__leaf_net291));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net291 (.A(clknet_0_net291),
    .X(clknet_1_1__leaf_net291));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net852 (.A(net852),
    .X(clknet_0_net852));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net852 (.A(clknet_0_net852),
    .X(clknet_1_0__leaf_net852));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net852 (.A(clknet_0_net852),
    .X(clknet_1_1__leaf_net852));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net841 (.A(net841),
    .X(clknet_0_net841));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net841 (.A(clknet_0_net841),
    .X(clknet_1_0__leaf_net841));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net841 (.A(clknet_0_net841),
    .X(clknet_1_1__leaf_net841));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net191 (.A(net191),
    .X(clknet_0_net191));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net191 (.A(clknet_0_net191),
    .X(clknet_1_0__leaf_net191));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net191 (.A(clknet_0_net191),
    .X(clknet_1_1__leaf_net191));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net604 (.A(net604),
    .X(clknet_0_net604));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net604 (.A(clknet_0_net604),
    .X(clknet_1_0__leaf_net604));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net604 (.A(clknet_0_net604),
    .X(clknet_1_1__leaf_net604));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net838 (.A(net838),
    .X(clknet_0_net838));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net838 (.A(clknet_0_net838),
    .X(clknet_1_0__leaf_net838));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net838 (.A(clknet_0_net838),
    .X(clknet_1_1__leaf_net838));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net862 (.A(net862),
    .X(clknet_0_net862));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net862 (.A(clknet_0_net862),
    .X(clknet_1_0__leaf_net862));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net862 (.A(clknet_0_net862),
    .X(clknet_1_1__leaf_net862));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net94 (.A(net94),
    .X(clknet_0_net94));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net94 (.A(clknet_0_net94),
    .X(clknet_1_0__leaf_net94));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net94 (.A(clknet_0_net94),
    .X(clknet_1_1__leaf_net94));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net836 (.A(net836),
    .X(clknet_0_net836));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net836 (.A(clknet_0_net836),
    .X(clknet_1_0__leaf_net836));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net836 (.A(clknet_0_net836),
    .X(clknet_1_1__leaf_net836));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net75 (.A(net75),
    .X(clknet_0_net75));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net75 (.A(clknet_0_net75),
    .X(clknet_1_0__leaf_net75));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net75 (.A(clknet_0_net75),
    .X(clknet_1_1__leaf_net75));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer1 (.A(net27),
    .X(net909));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer2 (.A(net909),
    .X(net910));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer3 (.A(net910),
    .X(net911));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer4 (.A(net363),
    .X(net912));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer5 (.A(net912),
    .X(net913));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer6 (.A(net912),
    .X(net914));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer7 (.A(net348),
    .X(net915));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer8 (.A(net24),
    .X(net916));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer9 (.A(net131),
    .X(net917));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer10 (.A(net134),
    .X(net918));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer11 (.A(net918),
    .X(net919));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer12 (.A(net918),
    .X(net920));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer13 (.A(net918),
    .X(net921));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer14 (.A(net939),
    .X(net922));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer15 (.A(net922),
    .X(net923));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer16 (.A(net939),
    .X(net924));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer17 (.A(net939),
    .X(net925));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer18 (.A(net41),
    .X(net926));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer19 (.A(net926),
    .X(net927));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer20 (.A(net599),
    .X(net928));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer21 (.A(net599),
    .X(net929));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer22 (.A(net356),
    .X(net930));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer23 (.A(net889),
    .X(net931));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer24 (.A(net931),
    .X(net932));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer25 (.A(net134),
    .X(net933));
 sky130_fd_sc_hd__buf_2 rebuffer26 (.A(net933),
    .X(net934));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer27 (.A(net133),
    .X(net935));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer28 (.A(net879),
    .X(net936));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer29 (.A(net936),
    .X(net937));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer30 (.A(net936),
    .X(net938));
 sky130_fd_sc_hd__clkbuf_1 clone31 (.A(net871),
    .X(net939));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer32 (.A(net871),
    .X(net940));
 sky130_fd_sc_hd__clkbuf_1 clone33 (.A(net889),
    .X(net941));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(net962),
    .X(net943));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(net624),
    .X(net944));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(net834),
    .X(net945));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(net644),
    .X(net946));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(net611),
    .X(net947));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(net632),
    .X(net948));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(net576),
    .X(net949));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(net817),
    .X(net950));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(net438),
    .X(net951));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(net589),
    .X(net952));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(net249),
    .X(net953));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(net647),
    .X(net954));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(net331),
    .X(net955));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(net332),
    .X(net956));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(net136),
    .X(net957));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(net622),
    .X(net958));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(net329),
    .X(net959));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(net442),
    .X(net960));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(net664),
    .X(net961));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(net672),
    .X(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_A (.DIODE(clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(in0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(in1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(in10));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(in11));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(in12));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(in13));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(in14));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(in15));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(in16));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(in17));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(in18));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(in19));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(in2));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(in20));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(in21));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(in22));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(in23));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(in24));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(in25));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(in26));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(in27));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_A (.DIODE(in28));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_A (.DIODE(in29));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_A (.DIODE(in3));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_A (.DIODE(in30));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_A (.DIODE(in31));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_A (.DIODE(in32));
 sky130_fd_sc_hd__diode_2 ANTENNA_input28_A (.DIODE(in33));
 sky130_fd_sc_hd__diode_2 ANTENNA_input29_A (.DIODE(in34));
 sky130_fd_sc_hd__diode_2 ANTENNA_input30_A (.DIODE(in35));
 sky130_fd_sc_hd__diode_2 ANTENNA_input31_A (.DIODE(in36));
 sky130_fd_sc_hd__diode_2 ANTENNA_input32_A (.DIODE(in37));
 sky130_fd_sc_hd__diode_2 ANTENNA_input33_A (.DIODE(in38));
 sky130_fd_sc_hd__diode_2 ANTENNA_input34_A (.DIODE(in39));
 sky130_fd_sc_hd__diode_2 ANTENNA_input35_A (.DIODE(in4));
 sky130_fd_sc_hd__diode_2 ANTENNA_input36_A (.DIODE(in40));
 sky130_fd_sc_hd__diode_2 ANTENNA_input37_A (.DIODE(in41));
 sky130_fd_sc_hd__diode_2 ANTENNA_input38_A (.DIODE(in42));
 sky130_fd_sc_hd__diode_2 ANTENNA_input39_A (.DIODE(in43));
 sky130_fd_sc_hd__diode_2 ANTENNA_input40_A (.DIODE(in44));
 sky130_fd_sc_hd__diode_2 ANTENNA_input41_A (.DIODE(in45));
 sky130_fd_sc_hd__diode_2 ANTENNA_input42_A (.DIODE(in46));
 sky130_fd_sc_hd__diode_2 ANTENNA_input43_A (.DIODE(in47));
 sky130_fd_sc_hd__diode_2 ANTENNA_input44_A (.DIODE(in48));
 sky130_fd_sc_hd__diode_2 ANTENNA_input45_A (.DIODE(in49));
 sky130_fd_sc_hd__diode_2 ANTENNA_input46_A (.DIODE(in5));
 sky130_fd_sc_hd__diode_2 ANTENNA_input47_A (.DIODE(in50));
 sky130_fd_sc_hd__diode_2 ANTENNA_input48_A (.DIODE(in51));
 sky130_fd_sc_hd__diode_2 ANTENNA_input49_A (.DIODE(in52));
 sky130_fd_sc_hd__diode_2 ANTENNA_input50_A (.DIODE(in54));
 sky130_fd_sc_hd__diode_2 ANTENNA_input51_A (.DIODE(in55));
 sky130_fd_sc_hd__diode_2 ANTENNA_input52_A (.DIODE(in56));
 sky130_fd_sc_hd__diode_2 ANTENNA_input53_A (.DIODE(in57));
 sky130_fd_sc_hd__diode_2 ANTENNA_input54_A (.DIODE(in58));
 sky130_fd_sc_hd__diode_2 ANTENNA_input55_A (.DIODE(in59));
 sky130_fd_sc_hd__diode_2 ANTENNA_input56_A (.DIODE(in6));
 sky130_fd_sc_hd__diode_2 ANTENNA_input57_A (.DIODE(in60));
 sky130_fd_sc_hd__diode_2 ANTENNA_input58_A (.DIODE(in61));
 sky130_fd_sc_hd__diode_2 ANTENNA_input59_A (.DIODE(in62));
 sky130_fd_sc_hd__diode_2 ANTENNA_input60_A (.DIODE(in63));
 sky130_fd_sc_hd__diode_2 ANTENNA_input61_A (.DIODE(in65));
 sky130_fd_sc_hd__diode_2 ANTENNA_input62_A (.DIODE(in66));
 sky130_fd_sc_hd__diode_2 ANTENNA_input63_A (.DIODE(in67));
 sky130_fd_sc_hd__diode_2 ANTENNA_input64_A (.DIODE(in68));
 sky130_fd_sc_hd__diode_2 ANTENNA_input65_A (.DIODE(in69));
 sky130_fd_sc_hd__diode_2 ANTENNA_input66_A (.DIODE(in7));
 sky130_fd_sc_hd__diode_2 ANTENNA_input67_A (.DIODE(in70));
 sky130_fd_sc_hd__diode_2 ANTENNA_input68_A (.DIODE(in71));
 sky130_fd_sc_hd__diode_2 ANTENNA_input69_A (.DIODE(in72));
 sky130_fd_sc_hd__diode_2 ANTENNA_input70_A (.DIODE(in73));
 sky130_fd_sc_hd__diode_2 ANTENNA_input71_A (.DIODE(in74));
 sky130_fd_sc_hd__diode_2 ANTENNA_input72_A (.DIODE(in75));
 sky130_fd_sc_hd__diode_2 ANTENNA_input73_A (.DIODE(in76));
 sky130_fd_sc_hd__diode_2 ANTENNA_input74_A (.DIODE(in77));
 sky130_fd_sc_hd__diode_2 ANTENNA_input75_A (.DIODE(in78));
 sky130_fd_sc_hd__diode_2 ANTENNA_input76_A (.DIODE(in79));
 sky130_fd_sc_hd__diode_2 ANTENNA_input77_A (.DIODE(in8));
 sky130_fd_sc_hd__diode_2 ANTENNA_input78_A (.DIODE(in80));
 sky130_fd_sc_hd__diode_2 ANTENNA_input79_A (.DIODE(in81));
 sky130_fd_sc_hd__diode_2 ANTENNA_input80_A (.DIODE(in82));
 sky130_fd_sc_hd__diode_2 ANTENNA_input81_A (.DIODE(in83));
 sky130_fd_sc_hd__diode_2 ANTENNA_input82_A (.DIODE(in84));
 sky130_fd_sc_hd__diode_2 ANTENNA_input83_A (.DIODE(in85));
 sky130_fd_sc_hd__diode_2 ANTENNA_input84_A (.DIODE(in86));
 sky130_fd_sc_hd__diode_2 ANTENNA_input85_A (.DIODE(in87));
 sky130_fd_sc_hd__diode_2 ANTENNA_input86_A (.DIODE(in88));
 sky130_fd_sc_hd__diode_2 ANTENNA_input87_A (.DIODE(in89));
 sky130_fd_sc_hd__diode_2 ANTENNA_input88_A (.DIODE(in9));
 sky130_fd_sc_hd__diode_2 ANTENNA_input89_A (.DIODE(in90));
 sky130_fd_sc_hd__diode_2 ANTENNA_input90_A (.DIODE(in91));
 sky130_fd_sc_hd__diode_2 ANTENNA_input91_A (.DIODE(in92));
 sky130_fd_sc_hd__diode_2 ANTENNA_input92_A (.DIODE(in93));
 sky130_fd_sc_hd__diode_2 ANTENNA_input93_A (.DIODE(in94));
 sky130_fd_sc_hd__diode_2 ANTENNA_input94_A (.DIODE(in95));
 sky130_fd_sc_hd__diode_2 ANTENNA_input95_A (.DIODE(in96));
 sky130_fd_sc_hd__diode_2 ANTENNA_input96_A (.DIODE(in97));
 sky130_fd_sc_hd__diode_2 ANTENNA_input97_A (.DIODE(in98));
 sky130_fd_sc_hd__diode_2 ANTENNA_input98_A (.DIODE(in99));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_B (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_A3 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA_c190_A1 (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_S1 (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_A (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_A2 (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c134_X (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_A2 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_A2 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c365_A3 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_A3 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c241_Q_N (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c557_A1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_A2 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_A3 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_A2 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA_c295_S1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA_c272_A2 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA_c266_A1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA_c264_Y (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge783_A0 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge780_A2 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c430_A3 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c286_A2 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_B1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c269_B (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_A (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c266_X (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout180_A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge765_S1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c272_X (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge773_D (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_A1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_A2 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_A2 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_B1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c283_A3 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_A3 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c277_A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c274_X (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout179_A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c633_A0 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c278_Y (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c431_D (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_c427_SCE (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_RESET_B (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_c276_B (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_A1 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_B1 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_A0 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_c136_X (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_A1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c564_A2 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c559_SET_B (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_A2 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_A1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_X (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge781_A2 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge774_A1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge768_S0 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge763_A2 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_RESET_B (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_A0 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_A3 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_SCE (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c408_A2 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_SCD (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_X (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_S0 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_D (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_B1_N (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_RESET_B (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c311_A3 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_A2 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c286_X (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout178_A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A0 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_S0 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_X (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A2 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_A0 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_A2 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c549_A3 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_A3 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c424_SET_B (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_A2 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_B1 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_A4 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_A2 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_X (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_A0 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_A3 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_A1 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_A1 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_A3 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_A1 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_c340_A1 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_A4 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_SCD (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_X (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A2 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA_c428_A2 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_B1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_D (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_A3 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_A3 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_A1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_X (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge788_A0 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_c424_SCD (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_A1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_A1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_X (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_c662_A1 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_c660_B (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_c541_A2 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_c397_A2 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_A3 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_A0 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_c143_B (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_Y (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge781_S1 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge764_A1 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_A2 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_RESET_B (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_A1 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_A3 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_X (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_A0 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA_c350_A3 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_A3 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_A2 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_A1 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_A1 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_A2 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_S0 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_X (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge766_A1 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_A2 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_A0 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_A1 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA_c344_A0 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_SCD (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_A3 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_A2 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_X (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_A2 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_A0 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_A1 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_A1 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA_c340_A4 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_Q_N (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_A1 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_A2 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c198_B1_N (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_A3 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_B (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_A2 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c143_Y (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_S1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_A2 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_A0 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_A2 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_SCE (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA_c540_S1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_A2 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_A2 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA_c415_A (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA_c414_S0 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA_c403_X (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_D (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_A2 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_A3 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_c286_B1_N (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_c273_B1 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_c267_A2 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_X (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_A1 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_A1 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_A0 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_B1_N (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_SCD (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_c414_A0 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_c412_A2 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_c410_A2 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_c409_X (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge785_A2 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_S0 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_A3 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_A1 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA_c556_A2 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_A0 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA_c415_B (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA_c411_X (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge770_A3 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_RESET_B (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_A2 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_D (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA_c415_Y (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA_c561_A (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge768_A1 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_A0 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_A1 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_c559_SCE (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_c548_A2 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_c544_S0 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_c541_S0 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_c416_X (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_A3 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_A3 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_A3 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c557_B1_N (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c528_B (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_Q_N (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c744_A2 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA_c660_A (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_A1 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_A1 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_A2 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_Q (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout172_A (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_A2 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge765_A1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_X (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge790_A3 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge770_A2 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_SET_B (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_X (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge786_A4 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge779_A3 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge763_A4 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA_c424_Q_N (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_A0 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_A0 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_A3 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA_c431_SCD (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA_c430_B1 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA_c427_SCD (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_X (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_A1 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_A2 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c434_SCE (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_Q (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge790_S0 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge788_A2 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge770_A0 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_A2 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA_c437_A4 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_A1 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_X (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_A2 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_A3 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_S1 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_Q_N (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_A0 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_A1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_A2 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_Q (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_A0 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_A3 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_X (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge788_S1 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_A1 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_A4 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_S0 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_S0 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_A3 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_S1 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_X (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_D (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_A4 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_X (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_A1 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_A3 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_A0 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_A3 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_Q (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_A0 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_D (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_A1 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_A1 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_X (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge783_S1 (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_A0 (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA_c586_A3 (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_S0 (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_A2 (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_S0 (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_X (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_A2 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_SCE (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_A3 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_A1 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_RESET_B (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_A0 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c373_A1 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_S1 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_X (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c563_A3 (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c556_A4 (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_A1 (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_SCE (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_B1 (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_A0 (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_A1 (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c158_A3 (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_X (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge789_S1 (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_A1 (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA_c681_A2 (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA_c678_A4 (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA_c532_B1_N (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA_c531_Y (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold51_A (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA_c563_A4 (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge784_S1 (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA_c540_S0 (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA_c536_X (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold48_A (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA_c676_SET_B (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA_c664_A (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA_c548_A1 (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA_c546_S1 (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA_c542_A2 (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA_c541_A3 (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA_c539_X (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_A1 (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA_c545_A1 (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA_c544_A3 (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA_c543_B1_N (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA_c542_X (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge776_A0 (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_A1 (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA_c547_SCD (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA_c543_X (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout187_A (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_A2 (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge779_S1 (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA_c545_X (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA_c611_A1 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_c549_A2 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_c547_SCE (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_c546_X (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_c700_A0 (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_A3 (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA_c681_A3 (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA_c549_A1 (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA_c547_Q (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge786_A3 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge779_S0 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge774_A2 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge773_SCD (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_A3 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_A0 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA_c559_SCD (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_Y (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_A0 (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_A2 (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_A2 (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_A2 (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_A4 (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_X (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_A1 (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_A3 (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_A0 (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_A3 (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA_c614_S0 (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA_c555_X (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA_c695_A3 (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA_c687_A1 (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_A2 (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA_c566_B1 (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA_c564_B1 (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA_c558_A2 (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA_c557_X (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA_c723_A0 (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_A1 (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_A1 (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_S0 (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_D (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA_c693_A2 (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA_c565_X (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_A1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_A3 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c424_D (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_A1 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c313_S0 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_A3 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_A1 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_X (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_A1 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_B1 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_c295_S0 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_A1 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_A1 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_B1 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_A2 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_B1 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_X (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge785_A0 (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge784_A2 (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge773_RESET_B (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge772_A3 (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA_c700_S1 (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA_c687_A2 (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_B1 (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_A1 (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_S0 (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA_c664_Y (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA_c720_A2 (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_S0 (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_S0 (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_A0 (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_S1 (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_A1 (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_S0 (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_A1 (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA_c674_SCE (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA_c669_A2 (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA_c666_X (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge790_A2 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge784_A0 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A0 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_A2 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A2 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA_c703_A2 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA_c700_S0 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA_c686_D (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA_c677_SCE (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA_c667_X (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA_c745_A3 (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_A2 (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA_c724_A3 (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_A1 (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_A0 (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_RESET_B (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA_c677_D (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA_c676_SCE (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA_c672_SET_B (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA_c670_X (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_A2 (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_A3 (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA_c675_A2 (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA_c674_Q_N (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA_c746_A2 (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA_c743_A2 (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_A0 (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_A2 (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_A2 (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA_c698_A2 (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_A2 (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_X (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_A1 (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_A1 (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_A2 (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA_c703_A3 (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA_c702_A3 (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA_c701_A2 (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA_c700_A1 (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA_c698_X (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge764_A2 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_A2 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_B1 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_A1 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_c215_A0 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_X (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_S0 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_A1 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_A0 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_D (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_A2 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_A1 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_c496_A3 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_A2 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_c108_X (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout196_A (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout195_A (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_A3 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_B1 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_B1 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_X (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_D (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_B1 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_A2 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_X (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_A1 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_A2 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_X (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge834_B (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA_c746_X (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge792_Q_N (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_A3 (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_S1 (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge794_Q (.DIODE(net575));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge774_A4 (.DIODE(net575));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_B1 (.DIODE(net575));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_S0 (.DIODE(net575));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_B1 (.DIODE(net575));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge797_Q (.DIODE(net577));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge785_S1 (.DIODE(net577));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_A3 (.DIODE(net577));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_A3 (.DIODE(net577));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge783_S0 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge770_A1 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_A0 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_X (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge845_Q (.DIODE(net628));
 sky130_fd_sc_hd__diode_2 ANTENNA_c723_A1 (.DIODE(net628));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_A2 (.DIODE(net628));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_S0 (.DIODE(net628));
 sky130_fd_sc_hd__diode_2 ANTENNA_c685_A2 (.DIODE(net628));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge847_Q (.DIODE(net629));
 sky130_fd_sc_hd__diode_2 ANTENNA_c747_S1 (.DIODE(net629));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_S0 (.DIODE(net629));
 sky130_fd_sc_hd__diode_2 ANTENNA_c670_A (.DIODE(net629));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_A (.DIODE(net629));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge764_A4 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_A2 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_c205_A2 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_A2 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_c194_A2 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_X (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge848_Q (.DIODE(net630));
 sky130_fd_sc_hd__diode_2 ANTENNA_c369_B1 (.DIODE(net630));
 sky130_fd_sc_hd__diode_2 ANTENNA_c368_S1 (.DIODE(net630));
 sky130_fd_sc_hd__diode_2 ANTENNA_c366_B1 (.DIODE(net630));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_A (.DIODE(net630));
 sky130_fd_sc_hd__diode_2 ANTENNA_c212_A (.DIODE(net630));
 sky130_fd_sc_hd__diode_2 ANTENNA_s851_Q (.DIODE(net634));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_A4 (.DIODE(net634));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_A3 (.DIODE(net634));
 sky130_fd_sc_hd__diode_2 ANTENNA_c371_S1 (.DIODE(net634));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_S1 (.DIODE(net634));
 sky130_fd_sc_hd__diode_2 ANTENNA_s852_Q (.DIODE(net635));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge776_S0 (.DIODE(net635));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_A2 (.DIODE(net635));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_A2 (.DIODE(net635));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_S1 (.DIODE(net635));
 sky130_fd_sc_hd__diode_2 ANTENNA_c611_B1 (.DIODE(net635));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_S1 (.DIODE(net635));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_S1 (.DIODE(net635));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_S0 (.DIODE(net635));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_S1 (.DIODE(net635));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_S1 (.DIODE(net635));
 sky130_fd_sc_hd__diode_2 ANTENNA_s862_Q (.DIODE(net646));
 sky130_fd_sc_hd__diode_2 ANTENNA_c744_S1 (.DIODE(net646));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_A3 (.DIODE(net646));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A4 (.DIODE(net646));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_S0 (.DIODE(net646));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_B1_N (.DIODE(net646));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_B1_N (.DIODE(net646));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_S1 (.DIODE(net646));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_B1_N (.DIODE(net646));
 sky130_fd_sc_hd__diode_2 ANTENNA_s865_Q (.DIODE(net649));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_S1 (.DIODE(net649));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_S1 (.DIODE(net649));
 sky130_fd_sc_hd__diode_2 ANTENNA_s874_Q (.DIODE(net658));
 sky130_fd_sc_hd__diode_2 ANTENNA_c693_B1_N (.DIODE(net658));
 sky130_fd_sc_hd__diode_2 ANTENNA_c679_S1 (.DIODE(net658));
 sky130_fd_sc_hd__diode_2 ANTENNA_c669_B1_N (.DIODE(net658));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_B1_N (.DIODE(net658));
 sky130_fd_sc_hd__diode_2 ANTENNA_s877_Q (.DIODE(net663));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge774_B1 (.DIODE(net663));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge772_B1 (.DIODE(net663));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_S1 (.DIODE(net663));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_S0 (.DIODE(net663));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_A4 (.DIODE(net663));
 sky130_fd_sc_hd__diode_2 ANTENNA_c678_B1 (.DIODE(net663));
 sky130_fd_sc_hd__diode_2 ANTENNA_s880_Q (.DIODE(net666));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_S1 (.DIODE(net666));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_B1 (.DIODE(net666));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_S1 (.DIODE(net666));
 sky130_fd_sc_hd__diode_2 ANTENNA_c587_S1 (.DIODE(net666));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge769_A0 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_A2 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_A2 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_D (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_S1 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_X (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA_s893_Q (.DIODE(net684));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_B1 (.DIODE(net684));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_S1 (.DIODE(net684));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_S1 (.DIODE(net684));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_SET_B (.DIODE(net684));
 sky130_fd_sc_hd__diode_2 ANTENNA_c703_S1 (.DIODE(net684));
 sky130_fd_sc_hd__diode_2 ANTENNA_s902_Q (.DIODE(net695));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_S0 (.DIODE(net695));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_A3 (.DIODE(net695));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_S1 (.DIODE(net695));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_S1 (.DIODE(net695));
 sky130_fd_sc_hd__diode_2 ANTENNA_c746_S1 (.DIODE(net695));
 sky130_fd_sc_hd__diode_2 ANTENNA_c743_S1 (.DIODE(net695));
 sky130_fd_sc_hd__diode_2 ANTENNA_c723_S1 (.DIODE(net695));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_S1 (.DIODE(net695));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_S1 (.DIODE(net695));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_A1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_S0 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_A0 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_A3 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_c239_A1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_c232_A3 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_c226_X (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_X (.DIODE(net707));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge785_A3 (.DIODE(net707));
 sky130_fd_sc_hd__diode_2 ANTENNA_c535_A1 (.DIODE(net707));
 sky130_fd_sc_hd__diode_2 ANTENNA_c400_B1 (.DIODE(net707));
 sky130_fd_sc_hd__diode_2 ANTENNA_c275_A2 (.DIODE(net707));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_A2 (.DIODE(net707));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_A1 (.DIODE(net707));
 sky130_fd_sc_hd__diode_2 ANTENNA_c134_A2 (.DIODE(net707));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_X (.DIODE(net708));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_A2 (.DIODE(net708));
 sky130_fd_sc_hd__diode_2 ANTENNA_c182_A1 (.DIODE(net708));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_B (.DIODE(net708));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_X (.DIODE(net713));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_A1 (.DIODE(net713));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_A3 (.DIODE(net713));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_A3 (.DIODE(net713));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_X (.DIODE(net715));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_A2 (.DIODE(net715));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_A3 (.DIODE(net715));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_S0 (.DIODE(net715));
 sky130_fd_sc_hd__diode_2 ANTENNA_c265_A (.DIODE(net715));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_A1 (.DIODE(net715));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_B1_N (.DIODE(net715));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_A4 (.DIODE(net715));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_A4 (.DIODE(net715));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_S0 (.DIODE(net715));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_X (.DIODE(net719));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_A2 (.DIODE(net719));
 sky130_fd_sc_hd__diode_2 ANTENNA_c140_B (.DIODE(net719));
 sky130_fd_sc_hd__diode_2 ANTENNA_c103_A3 (.DIODE(net719));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_X (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_D (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_A2 (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_A1 (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_A2 (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_B (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_B1 (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA_c102_A3 (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_X (.DIODE(net723));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_A2 (.DIODE(net723));
 sky130_fd_sc_hd__diode_2 ANTENNA_c184_A0 (.DIODE(net723));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_S0 (.DIODE(net723));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_A3 (.DIODE(net723));
 sky130_fd_sc_hd__diode_2 ANTENNA_c108_A1 (.DIODE(net723));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_X (.DIODE(net724));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_A1 (.DIODE(net724));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_A3 (.DIODE(net724));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_X (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_B1_N (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA_c203_A1 (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_A2 (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_A2 (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_B1_N (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_X (.DIODE(net726));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge770_S1 (.DIODE(net726));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_S1 (.DIODE(net726));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_A0 (.DIODE(net726));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_A1 (.DIODE(net726));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_A2 (.DIODE(net726));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_A3 (.DIODE(net726));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_B1 (.DIODE(net726));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_A2 (.DIODE(net726));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_A2 (.DIODE(net726));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_X (.DIODE(net729));
 sky130_fd_sc_hd__diode_2 ANTENNA_c183_A1 (.DIODE(net729));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_A1 (.DIODE(net729));
 sky130_fd_sc_hd__diode_2 ANTENNA_input32_X (.DIODE(net736));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_A1 (.DIODE(net736));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_A3 (.DIODE(net736));
 sky130_fd_sc_hd__diode_2 ANTENNA_input34_X (.DIODE(net738));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_D (.DIODE(net738));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_SET_B (.DIODE(net738));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_A2 (.DIODE(net738));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_A1 (.DIODE(net738));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_A3 (.DIODE(net738));
 sky130_fd_sc_hd__diode_2 ANTENNA_input36_X (.DIODE(net740));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_B1_N (.DIODE(net740));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_A2 (.DIODE(net740));
 sky130_fd_sc_hd__diode_2 ANTENNA_c127_A0 (.DIODE(net740));
 sky130_fd_sc_hd__diode_2 ANTENNA_c108_A3 (.DIODE(net740));
 sky130_fd_sc_hd__diode_2 ANTENNA_c100_A4 (.DIODE(net740));
 sky130_fd_sc_hd__diode_2 ANTENNA_input38_X (.DIODE(net742));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge767_A3 (.DIODE(net742));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_A2 (.DIODE(net742));
 sky130_fd_sc_hd__diode_2 ANTENNA_input40_X (.DIODE(net744));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_A2 (.DIODE(net744));
 sky130_fd_sc_hd__diode_2 ANTENNA_c366_A4 (.DIODE(net744));
 sky130_fd_sc_hd__diode_2 ANTENNA_c180_A2 (.DIODE(net744));
 sky130_fd_sc_hd__diode_2 ANTENNA_c107_S0 (.DIODE(net744));
 sky130_fd_sc_hd__diode_2 ANTENNA_c104_A3 (.DIODE(net744));
 sky130_fd_sc_hd__diode_2 ANTENNA_input41_X (.DIODE(net745));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_A2 (.DIODE(net745));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_S0 (.DIODE(net745));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_B1_N (.DIODE(net745));
 sky130_fd_sc_hd__diode_2 ANTENNA_input43_X (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge764_B1 (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_A1 (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_SET_B (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_A0 (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA_input45_X (.DIODE(net749));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge790_S1 (.DIODE(net749));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge766_S1 (.DIODE(net749));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_A2 (.DIODE(net749));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_A0 (.DIODE(net749));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_B1_N (.DIODE(net749));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_A1 (.DIODE(net749));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_A3 (.DIODE(net749));
 sky130_fd_sc_hd__diode_2 ANTENNA_input46_X (.DIODE(net750));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_A3 (.DIODE(net750));
 sky130_fd_sc_hd__diode_2 ANTENNA_c274_A1 (.DIODE(net750));
 sky130_fd_sc_hd__diode_2 ANTENNA_c158_A1 (.DIODE(net750));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_A3 (.DIODE(net750));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_A1 (.DIODE(net750));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_B (.DIODE(net750));
 sky130_fd_sc_hd__diode_2 ANTENNA_c134_B1_N (.DIODE(net750));
 sky130_fd_sc_hd__diode_2 ANTENNA_input48_X (.DIODE(net752));
 sky130_fd_sc_hd__diode_2 ANTENNA_c614_A2 (.DIODE(net752));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_A1 (.DIODE(net752));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_A1 (.DIODE(net752));
 sky130_fd_sc_hd__diode_2 ANTENNA_c313_S1 (.DIODE(net752));
 sky130_fd_sc_hd__diode_2 ANTENNA_input52_X (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_A4 (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA_c194_S0 (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_B1 (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA_c104_A1 (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA_input54_X (.DIODE(net758));
 sky130_fd_sc_hd__diode_2 ANTENNA_c364_A0 (.DIODE(net758));
 sky130_fd_sc_hd__diode_2 ANTENNA_c226_A4 (.DIODE(net758));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_S0 (.DIODE(net758));
 sky130_fd_sc_hd__diode_2 ANTENNA_input55_X (.DIODE(net759));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_A1 (.DIODE(net759));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_B1_N (.DIODE(net759));
 sky130_fd_sc_hd__diode_2 ANTENNA_input57_X (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_A1 (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_B1_N (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_A1 (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_input58_X (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_A0 (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_A2 (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_A2 (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_A1 (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_A2 (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA_input59_X (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge767_A1 (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_A2 (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA_c206_A4 (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA_input60_X (.DIODE(net764));
 sky130_fd_sc_hd__diode_2 ANTENNA_c761_A0 (.DIODE(net764));
 sky130_fd_sc_hd__diode_2 ANTENNA_c757_A1 (.DIODE(net764));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A1 (.DIODE(net764));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_A2 (.DIODE(net764));
 sky130_fd_sc_hd__diode_2 ANTENNA_input62_X (.DIODE(net766));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_A3 (.DIODE(net766));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_A2 (.DIODE(net766));
 sky130_fd_sc_hd__diode_2 ANTENNA_c124_A1 (.DIODE(net766));
 sky130_fd_sc_hd__diode_2 ANTENNA_input64_X (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_A3 (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_A1 (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA_input66_X (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c759_A2 (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_A3 (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_B1_N (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_S1 (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_A4 (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_A1 (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_A2 (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_A3 (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_A1 (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_input67_X (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_c368_A3 (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_D (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_A1 (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_input69_X (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_A0 (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_A1 (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_A2 (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_A2 (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_S0 (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA_c203_A3 (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_B1_N (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA_c104_B1 (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA_input72_X (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c127_A2 (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c103_S1 (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_input80_X (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA_c369_A1 (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA_c215_A3 (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA_c206_A2 (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA_input81_X (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_c368_A0 (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_c226_A3 (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_input83_X (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_A3 (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_S0 (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_S0 (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_A1 (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c229_A1 (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_B1_N (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c205_B1 (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_input84_X (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_A1 (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_A2 (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_B1_N (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA_input88_X (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_A1 (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_c273_A3 (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_B (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_c158_A2 (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_c138_B (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_input92_X (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge769_A1 (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA_c241_D (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA_c123_A2 (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA_c122_A3 (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA_c107_A1 (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA_c106_B1 (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA_c100_A2 (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA_input97_X (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_c364_A2 (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_B1 (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_SCD (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_RESET_B (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_B1 (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_c124_B1 (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_c109_A2 (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_c102_B1 (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_output99_A (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA_c615_A3 (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA_c613_A2 (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA_c610_X (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA_output100_A (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_A3 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_A4 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_Q (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_output101_A (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_S0 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_A1 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_A3 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_Q (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_output102_A (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA_c614_X (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA_output103_A (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_c615_X (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_output104_A (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge765_A2 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_A2 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_S0 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_B1_N (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c228_A3 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_S0 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_A1 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_X (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_output106_A (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge795_Q (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_A2 (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_output107_A (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge818_Q (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_A2 (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net812_A (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_X (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_output109_A (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge836_Q_N (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_S0 (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_output110_A (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge789_S0 (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_A2 (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_A1 (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_S0 (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_A2 (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_A0 (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_A2 (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_c545_A2 (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_c533_X (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_output111_A (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge835_Q (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_c633_A3 (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold42_A (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_output113_A (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_s853_Q (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_B1 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_A3 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_S0 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_S0 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_S1 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c346_S0 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_SCD (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_B1_N (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_output114_A (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge783_A2 (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_A0 (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_A3 (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_SCE (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_A0 (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c430_X (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_output115_A (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_A1 (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_A1 (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_c494_A3 (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_A3 (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_X (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout177_A (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_output118_A (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_X (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_output119_A (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge839_Q (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_c760_A3 (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_c759_S0 (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_S1 (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net824_A (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_c364_X (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_output122_A (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_A1 (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_X (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_output125_A (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_s869_Q (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c482_S1 (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_output126_A (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge814_Q (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_A3 (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_A (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_A (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA_output128_A (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_s867_Q (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_S1 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_S1 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_output129_A (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_s870_Q (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_S0 (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold37_A (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_output130_A (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_A1 (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_A1 (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_c241_Q (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_output133_A (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_A0 (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c340_A3 (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c240_A4 (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c222_A4 (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c203_A2 (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c198_X (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_output135_A (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge782_A3 (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_X (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_output139_A (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge808_Q (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c372_S1 (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c370_S0 (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c369_A4 (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_output141_A (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_c373_S0 (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_c372_A2 (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_c369_X (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_output142_A (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_c370_A1 (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_SCD (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_c241_SCE (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_c235_X (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout181_A (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_c368_S0 (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_A3 (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_X (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_output144_A (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_A2 (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_SCD (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_A3 (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_A0 (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_A2 (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_c434_SET_B (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_X (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_output145_A (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_A3 (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_B1_N (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c215_A1 (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_B1_N (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c206_A3 (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c205_A3 (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c203_B1 (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_A2 (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_X (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_output146_A (.DIODE(net850));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_A3 (.DIODE(net850));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_A1 (.DIODE(net850));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_X (.DIODE(net850));
 sky130_fd_sc_hd__diode_2 ANTENNA_output147_A (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge846_Q (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge777_S0 (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_B1 (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_c240_B1 (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_c236_B1_N (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_c235_A (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_c234_A (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_c220_A (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_A (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_output150_A (.DIODE(net854));
 sky130_fd_sc_hd__diode_2 ANTENNA_c241_SCD (.DIODE(net854));
 sky130_fd_sc_hd__diode_2 ANTENNA_c240_A1 (.DIODE(net854));
 sky130_fd_sc_hd__diode_2 ANTENNA_c239_X (.DIODE(net854));
 sky130_fd_sc_hd__diode_2 ANTENNA_output152_A (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_s850_Q (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_c502_S0 (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_A3 (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_c482_A2 (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_S1 (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_c340_B1 (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_c218_S1 (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_output155_A (.DIODE(net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge827_Q (.DIODE(net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_c238_B1_N (.DIODE(net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_B1_N (.DIODE(net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_c208_A (.DIODE(net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_A (.DIODE(net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_output156_A (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_c131_A3 (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_c129_S0 (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_c128_S1 (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_c127_S0 (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_c126_A2 (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_c125_A2 (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_c124_A3 (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_c123_A3 (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_c122_X (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_output157_A (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_c191_A2 (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_A3 (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_X (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_output160_A (.DIODE(net864));
 sky130_fd_sc_hd__diode_2 ANTENNA_c109_A3 (.DIODE(net864));
 sky130_fd_sc_hd__diode_2 ANTENNA_c106_X (.DIODE(net864));
 sky130_fd_sc_hd__diode_2 ANTENNA_output162_A (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_c236_A2 (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_c231_B1_N (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_c230_B1_N (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_X (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_output163_A (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c228_A2 (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_A3 (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_X (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_output164_A (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge787_S1 (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_A2 (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_A2 (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_A2 (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_A2 (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_A2 (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_A1 (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_A2 (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_c208_X (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_output165_A (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_c105_A4 (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_c103_X (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_output169_A (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c107_S1 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c102_X (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout172_X (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA_c424_SCE (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA_c427_RESET_B (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_A3 (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_A2 (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_A0 (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_A2 (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA_c695_A2 (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_A2 (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA_c687_A3 (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_A3 (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout173_X (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_A3 (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_SCE (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_S1 (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_A3 (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_c759_A0 (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge776_A3 (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A3 (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_c611_A2 (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_A0 (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge788_S0 (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap174_X (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c675_A1 (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c662_A2 (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c661_B (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge768_A3 (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c529_B (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c404_A2 (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer28_A (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_A1 (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout175_X (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_A2 (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_SCD (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_A2 (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_A3 (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_c297_A3 (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout176_X (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_A3 (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_S0 (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_A2 (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_A2 (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_A3 (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_A3 (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c739_A1 (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_A3 (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_A1 (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_A4 (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout177_X (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c502_A3 (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_A2 (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_A3 (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c496_A2 (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_A3 (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_A3 (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_A0 (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c369_A3 (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c366_A3 (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_A1 (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout178_X (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_A1 (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_S0 (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_A1 (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_B1 (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_A1 (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_A3 (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_A1 (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_A2 (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_A2 (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_A2 (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout179_X (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_A3 (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_A2 (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_A2 (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_A3 (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge764_A3 (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge788_A1 (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c531_B (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_S1 (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c313_A2 (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_A3 (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout180_X (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_c283_S0 (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_A3 (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_A4 (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_A2 (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_c743_A0 (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_A3 (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_A1 (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_A0 (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_c667_A1 (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_c663_A2 (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout181_X (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_A2 (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_A2 (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_A2 (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_A3 (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_A2 (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_c184_A3 (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_output143_A (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_A2 (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_A2 (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_c183_B1_N (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout187_X (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c762_A0 (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_A2 (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_A1 (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_A3 (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_A2 (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_A3 (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c679_A3 (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c548_A3 (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c547_SET_B (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c546_A3 (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c182_B1_N (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout188_X (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_A2 (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_A3 (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_c295_A1 (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_S0 (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout191_X (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_B1 (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_c613_S1 (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout190_A (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_SET_B (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_S1 (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout189_A (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout192_X (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge775_S1 (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_S1 (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_S1 (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_A2 (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_S1 (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c222_B1 (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_B1_N (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_B1_N (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_B1 (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_S1 (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout193_X (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_output116_A (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge769_S1 (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_A3 (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_A3 (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_SET_B (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c239_B1_N (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_SET_B (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c226_B1 (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout196_X (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge776_A2 (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_A2 (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_B1_N (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_A0 (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_A0 (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_S0 (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_A2 (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_A4 (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_RESET_B (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_A2 (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout198_X (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout197_A (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_A2 (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_S0 (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge776_A1 (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_c557_A2 (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_A1 (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout199_X (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_A2 (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_A2 (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_c368_A2 (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_A1 (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout198_A (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout200_X (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout199_A (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_output159_A (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A3 (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A4 (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_A1 (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_S0 (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_A4 (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c560_B1_N (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout201_X (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_A3 (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c398_B (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c279_B1_N (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c274_B1_N (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c266_B1_N (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_B1 (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_B1_N (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_B1 (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_S1 (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_B1_N (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout202_X (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_S0 (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout201_A (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_A1 (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_S1 (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_c558_B1_N (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout203_X (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge775_A3 (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_c742_A3 (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_A3 (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_A1 (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_A3 (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_SCD (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout202_A (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout204_X (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c184_A2 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_A1 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_S0 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c128_S0 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c125_B1 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_A3 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_A0 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_A0 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_A3 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c566_A4 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_15_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_14_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_13_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_12_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_11_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_10_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_9_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_8_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_7_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_6_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_5_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_4_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_3_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_2_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_1_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_0_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_X (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c673_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c676_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c677_CLK_N (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c686_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge832_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge845_GATE_N (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s888_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s889_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s890_GATE_N (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s891_GATE_N (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s892_GATE (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_0_0_clk_X (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c672_CLK_N (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c674_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge773_CLK_N (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge793_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge800_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge842_GATE (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge847_GATE (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s875_GATE_N (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s876_GATE (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s877_GATE_N (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_1_0_clk_X (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge795_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge813_GATE (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge820_GATE (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge836_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge837_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge838_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s904_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s906_GATE_N (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_8_0_clk_X (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge821_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge835_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s859_GATE_N (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s884_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s885_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s886_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s887_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s905_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_10_0_clk_X (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge824_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge826_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge839_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge849_GATE (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s867_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s868_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s870_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s871_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s872_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_11_0_clk_X (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_CLK_N (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_CLK_N (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge808_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge830_CLK_N (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge844_GATE_N (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s854_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s856_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s858_GATE_N (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s873_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s908_GATE (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_14_0_clk_X (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_CLK_N (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c241_CLK_N (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_CLK_N (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge815_GATE_N (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge825_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge846_GATE_N (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s855_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s857_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_15_0_clk_X (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_A3 (.DIODE(clknet_1_1__leaf_net809));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_A2 (.DIODE(clknet_1_1__leaf_net809));
 sky130_fd_sc_hd__diode_2 ANTENNA_output105_A (.DIODE(clknet_1_1__leaf_net809));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net809_X (.DIODE(clknet_1_1__leaf_net809));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_A3 (.DIODE(clknet_1_0__leaf_net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_A1 (.DIODE(clknet_1_0__leaf_net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_A3 (.DIODE(clknet_1_0__leaf_net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_output120_A (.DIODE(clknet_1_0__leaf_net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net824_X (.DIODE(clknet_1_0__leaf_net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_SCD (.DIODE(clknet_1_0__leaf_net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_A2 (.DIODE(clknet_1_0__leaf_net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_A3 (.DIODE(clknet_1_0__leaf_net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_A2 (.DIODE(clknet_1_0__leaf_net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_output108_A (.DIODE(clknet_1_0__leaf_net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net812_X (.DIODE(clknet_1_0__leaf_net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_A3 (.DIODE(clknet_1_0__leaf_net291));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_S0 (.DIODE(clknet_1_0__leaf_net291));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_A3 (.DIODE(clknet_1_0__leaf_net291));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_A3 (.DIODE(clknet_1_0__leaf_net291));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_A2 (.DIODE(clknet_1_0__leaf_net291));
 sky130_fd_sc_hd__diode_2 ANTENNA_c613_A3 (.DIODE(clknet_1_0__leaf_net291));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge779_A2 (.DIODE(clknet_1_0__leaf_net291));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net291_X (.DIODE(clknet_1_0__leaf_net291));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer2_A (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_c368_A1 (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer1_X (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_c615_A2 (.DIODE(net912));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer6_A (.DIODE(net912));
 sky130_fd_sc_hd__diode_2 ANTENNA_c587_A3 (.DIODE(net912));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer5_A (.DIODE(net912));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer4_X (.DIODE(net912));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_A0 (.DIODE(net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer9_X (.DIODE(net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer13_A (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_D (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer12_A (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_RESET_B (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer11_A (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer10_X (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_A1 (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer15_A (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer14_X (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_S1 (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer17_A (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer14_A (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer16_A (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone31_X (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_A0 (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer32_X (.DIODE(net940));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer31 (.A(net348),
    .X(net942));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer33 (.A(net27),
    .X(net963));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer34 (.A(net31),
    .X(net964));
 sky130_fd_sc_hd__a21bo_1 clone35 (.A1(net30),
    .A2(net707),
    .B1_N(net901),
    .X(net965));
 sky130_fd_sc_hd__a21bo_1 clone36 (.A1(net144),
    .A2(net707),
    .B1_N(net750),
    .X(net966));
 sky130_fd_sc_hd__clkbuf_1 clone37 (.A(net863),
    .X(net967));
 sky130_fd_sc_hd__a31o_1 clone38 (.A1(net719),
    .A2(net35),
    .A3(net32),
    .B1(net901),
    .X(net968));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_283 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_301 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_283 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_394 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_62 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_355 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_395 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_115 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_274 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_356 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_67 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_189 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_366 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_199 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_359 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_394 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_394 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_497 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_244 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_327 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_186 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_112 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_270 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_172 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_413 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_338 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_143 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_163 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_224 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_140 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_478 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_387 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_67 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_144 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_247 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_267 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_383 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_103 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_155 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_299 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_516 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_491 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_412 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_103 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_87 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_135 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_239 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_499 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_143 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_357 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_115 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_143 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_102 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_423 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_428 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_525 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_491 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_189 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_497 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_479 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_525 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_497 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_283 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_357 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_14 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_20 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_282 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_507 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_611 ();
endmodule
