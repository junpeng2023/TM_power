module netlist_0 (clk,
    in0,
    in1,
    in10,
    in11,
    in12,
    in13,
    in14,
    in15,
    in16,
    in17,
    in18,
    in19,
    in2,
    in20,
    in21,
    in22,
    in23,
    in24,
    in25,
    in26,
    in27,
    in28,
    in29,
    in3,
    in30,
    in31,
    in32,
    in33,
    in34,
    in35,
    in36,
    in37,
    in38,
    in39,
    in4,
    in40,
    in41,
    in42,
    in43,
    in44,
    in45,
    in46,
    in47,
    in48,
    in49,
    in5,
    in50,
    in51,
    in52,
    in53,
    in54,
    in55,
    in56,
    in57,
    in58,
    in59,
    in6,
    in60,
    in61,
    in62,
    in63,
    in64,
    in65,
    in66,
    in67,
    in68,
    in69,
    in7,
    in70,
    in71,
    in72,
    in73,
    in74,
    in75,
    in76,
    in77,
    in78,
    in79,
    in8,
    in80,
    in81,
    in82,
    in83,
    in84,
    in85,
    in86,
    in87,
    in88,
    in89,
    in9,
    in90,
    in91,
    in92,
    in93,
    in94,
    in95,
    in96,
    in97,
    in98,
    in99,
    out0,
    out1,
    out10,
    out11,
    out12,
    out13,
    out14,
    out15,
    out16,
    out17,
    out18,
    out19,
    out2,
    out20,
    out21,
    out22,
    out23,
    out24,
    out25,
    out26,
    out27,
    out28,
    out29,
    out3,
    out30,
    out31,
    out32,
    out33,
    out34,
    out35,
    out36,
    out37,
    out38,
    out39,
    out4,
    out40,
    out41,
    out42,
    out43,
    out44,
    out45,
    out46,
    out47,
    out48,
    out49,
    out5,
    out50,
    out51,
    out52,
    out53,
    out54,
    out55,
    out56,
    out57,
    out58,
    out59,
    out6,
    out60,
    out61,
    out62,
    out63,
    out64,
    out65,
    out66,
    out67,
    out68,
    out69,
    out7,
    out70,
    out71,
    out72,
    out73,
    out74,
    out75,
    out76,
    out77,
    out78,
    out79,
    out8,
    out80,
    out81,
    out82,
    out83,
    out84,
    out85,
    out86,
    out87,
    out88,
    out89,
    out9,
    out90,
    out91,
    out92,
    out93,
    out94,
    out95,
    out96,
    out97,
    out98,
    out99,
    rst);
 input clk;
 input in0;
 input in1;
 input in10;
 input in11;
 input in12;
 input in13;
 input in14;
 input in15;
 input in16;
 input in17;
 input in18;
 input in19;
 input in2;
 input in20;
 input in21;
 input in22;
 input in23;
 input in24;
 input in25;
 input in26;
 input in27;
 input in28;
 input in29;
 input in3;
 input in30;
 input in31;
 input in32;
 input in33;
 input in34;
 input in35;
 input in36;
 input in37;
 input in38;
 input in39;
 input in4;
 input in40;
 input in41;
 input in42;
 input in43;
 input in44;
 input in45;
 input in46;
 input in47;
 input in48;
 input in49;
 input in5;
 input in50;
 input in51;
 input in52;
 input in53;
 input in54;
 input in55;
 input in56;
 input in57;
 input in58;
 input in59;
 input in6;
 input in60;
 input in61;
 input in62;
 input in63;
 input in64;
 input in65;
 input in66;
 input in67;
 input in68;
 input in69;
 input in7;
 input in70;
 input in71;
 input in72;
 input in73;
 input in74;
 input in75;
 input in76;
 input in77;
 input in78;
 input in79;
 input in8;
 input in80;
 input in81;
 input in82;
 input in83;
 input in84;
 input in85;
 input in86;
 input in87;
 input in88;
 input in89;
 input in9;
 input in90;
 input in91;
 input in92;
 input in93;
 input in94;
 input in95;
 input in96;
 input in97;
 input in98;
 input in99;
 output out0;
 output out1;
 output out10;
 output out11;
 output out12;
 output out13;
 output out14;
 output out15;
 output out16;
 output out17;
 output out18;
 output out19;
 output out2;
 output out20;
 output out21;
 output out22;
 output out23;
 output out24;
 output out25;
 output out26;
 output out27;
 output out28;
 output out29;
 output out3;
 output out30;
 output out31;
 output out32;
 output out33;
 output out34;
 output out35;
 output out36;
 output out37;
 output out38;
 output out39;
 output out4;
 output out40;
 output out41;
 output out42;
 output out43;
 output out44;
 output out45;
 output out46;
 output out47;
 output out48;
 output out49;
 output out5;
 output out50;
 output out51;
 output out52;
 output out53;
 output out54;
 output out55;
 output out56;
 output out57;
 output out58;
 output out59;
 output out6;
 output out60;
 output out61;
 output out62;
 output out63;
 output out64;
 output out65;
 output out66;
 output out67;
 output out68;
 output out69;
 output out7;
 output out70;
 output out71;
 output out72;
 output out73;
 output out74;
 output out75;
 output out76;
 output out77;
 output out78;
 output out79;
 output out8;
 output out80;
 output out81;
 output out82;
 output out83;
 output out84;
 output out85;
 output out86;
 output out87;
 output out88;
 output out89;
 output out9;
 output out90;
 output out91;
 output out92;
 output out93;
 output out94;
 output out95;
 output out96;
 output out97;
 output out98;
 output out99;
 input rst;

 wire net0;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net63;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net64;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net65;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net66;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net67;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net68;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net69;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net7;
 wire net70;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net71;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net72;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net73;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net74;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net75;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net76;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net77;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net165;
 wire net465;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_0_net775;
 wire clknet_1_0__leaf_net775;
 wire clknet_1_1__leaf_net775;
 wire clknet_0_net883;
 wire clknet_1_0__leaf_net883;
 wire clknet_1_1__leaf_net883;
 wire clknet_0_net533;
 wire clknet_1_0__leaf_net533;
 wire clknet_1_1__leaf_net533;
 wire clknet_0_net945;
 wire clknet_1_0__leaf_net945;
 wire clknet_1_1__leaf_net945;
 wire clknet_0_net758;
 wire clknet_1_0__leaf_net758;
 wire clknet_1_1__leaf_net758;
 wire clknet_0_net489;
 wire clknet_1_0__leaf_net489;
 wire clknet_1_1__leaf_net489;
 wire clknet_0_net487;
 wire clknet_1_0__leaf_net487;
 wire clknet_1_1__leaf_net487;
 wire clknet_0_net757;
 wire clknet_1_0__leaf_net757;
 wire clknet_1_1__leaf_net757;
 wire clknet_0_net484;
 wire clknet_1_0__leaf_net484;
 wire clknet_1_1__leaf_net484;
 wire clknet_0_net504;
 wire clknet_1_0__leaf_net504;
 wire clknet_1_1__leaf_net504;
 wire clknet_0_net506;
 wire clknet_1_0__leaf_net506;
 wire clknet_1_1__leaf_net506;
 wire clknet_0_net511;
 wire clknet_1_0__leaf_net511;
 wire clknet_1_1__leaf_net511;
 wire clknet_0_net481;
 wire clknet_1_0__leaf_net481;
 wire clknet_1_1__leaf_net481;
 wire clknet_0_net502;
 wire clknet_1_0__leaf_net502;
 wire clknet_1_1__leaf_net502;
 wire clknet_0_net497;
 wire clknet_1_0__leaf_net497;
 wire clknet_1_1__leaf_net497;
 wire clknet_0_net756;
 wire clknet_1_0__leaf_net756;
 wire clknet_1_1__leaf_net756;
 wire clknet_0_net527;
 wire clknet_1_0__leaf_net527;
 wire clknet_1_1__leaf_net527;
 wire clknet_0_net740;
 wire clknet_1_0__leaf_net740;
 wire clknet_1_1__leaf_net740;
 wire clknet_0_net399;
 wire clknet_1_0__leaf_net399;
 wire clknet_1_1__leaf_net399;
 wire clknet_0_net899;
 wire clknet_1_0__leaf_net899;
 wire clknet_1_1__leaf_net899;
 wire clknet_0_net428;
 wire clknet_1_0__leaf_net428;
 wire clknet_1_1__leaf_net428;
 wire clknet_0_net420;
 wire clknet_1_0__leaf_net420;
 wire clknet_1_1__leaf_net420;
 wire clknet_0_net421;
 wire clknet_1_0__leaf_net421;
 wire clknet_1_1__leaf_net421;
 wire clknet_0_net400;
 wire clknet_1_0__leaf_net400;
 wire clknet_1_1__leaf_net400;
 wire clknet_0_net739;
 wire clknet_1_0__leaf_net739;
 wire clknet_1_1__leaf_net739;
 wire clknet_0_net405;
 wire clknet_1_0__leaf_net405;
 wire clknet_1_1__leaf_net405;
 wire clknet_0_net404;
 wire clknet_1_0__leaf_net404;
 wire clknet_1_1__leaf_net404;
 wire clknet_0_net884;
 wire clknet_1_0__leaf_net884;
 wire clknet_1_1__leaf_net884;
 wire clknet_0_net495;
 wire clknet_1_0__leaf_net495;
 wire clknet_1_1__leaf_net495;
 wire clknet_0_net494;
 wire clknet_1_0__leaf_net494;
 wire clknet_1_1__leaf_net494;
 wire clknet_0_net446;
 wire clknet_1_0__leaf_net446;
 wire clknet_1_1__leaf_net446;
 wire clknet_0_net908;
 wire clknet_1_0__leaf_net908;
 wire clknet_1_1__leaf_net908;
 wire clknet_0_net892;
 wire clknet_1_0__leaf_net892;
 wire clknet_1_1__leaf_net892;
 wire clknet_0_net402;
 wire clknet_1_0__leaf_net402;
 wire clknet_1_1__leaf_net402;
 wire clknet_0_net738;
 wire clknet_1_0__leaf_net738;
 wire clknet_1_1__leaf_net738;
 wire clknet_0_net721;
 wire clknet_1_0__leaf_net721;
 wire clknet_1_1__leaf_net721;
 wire clknet_0_net355;
 wire clknet_1_0__leaf_net355;
 wire clknet_1_1__leaf_net355;
 wire clknet_0_net361;
 wire clknet_1_0__leaf_net361;
 wire clknet_1_1__leaf_net361;
 wire clknet_0_net486;
 wire clknet_1_0__leaf_net486;
 wire clknet_1_1__leaf_net486;
 wire clknet_0_net394;
 wire clknet_1_0__leaf_net394;
 wire clknet_1_1__leaf_net394;
 wire clknet_0_net365;
 wire clknet_1_0__leaf_net365;
 wire clknet_1_1__leaf_net365;
 wire clknet_0_net645;
 wire clknet_1_0__leaf_net645;
 wire clknet_1_1__leaf_net645;
 wire clknet_0_net391;
 wire clknet_1_0__leaf_net391;
 wire clknet_1_1__leaf_net391;
 wire clknet_0_net376;
 wire clknet_1_0__leaf_net376;
 wire clknet_1_1__leaf_net376;
 wire clknet_0_net375;
 wire clknet_1_0__leaf_net375;
 wire clknet_1_1__leaf_net375;
 wire clknet_0_net473;
 wire clknet_1_0__leaf_net473;
 wire clknet_1_1__leaf_net473;
 wire clknet_0_net476;
 wire clknet_1_0__leaf_net476;
 wire clknet_1_1__leaf_net476;
 wire clknet_0_net612;
 wire clknet_1_0__leaf_net612;
 wire clknet_1_1__leaf_net612;
 wire clknet_0_net387;
 wire clknet_1_0__leaf_net387;
 wire clknet_1_1__leaf_net387;
 wire clknet_0_net389;
 wire clknet_1_0__leaf_net389;
 wire clknet_1_1__leaf_net389;
 wire clknet_0_net366;
 wire clknet_1_0__leaf_net366;
 wire clknet_1_1__leaf_net366;
 wire clknet_0_net388;
 wire clknet_1_0__leaf_net388;
 wire clknet_1_1__leaf_net388;
 wire clknet_0_net909;
 wire clknet_1_0__leaf_net909;
 wire clknet_1_1__leaf_net909;
 wire clknet_0_net379;
 wire clknet_1_0__leaf_net379;
 wire clknet_1_1__leaf_net379;
 wire clknet_0_net368;
 wire clknet_1_0__leaf_net368;
 wire clknet_1_1__leaf_net368;
 wire clknet_0_net369;
 wire clknet_1_0__leaf_net369;
 wire clknet_1_1__leaf_net369;
 wire clknet_0_net358;
 wire clknet_1_0__leaf_net358;
 wire clknet_1_1__leaf_net358;
 wire clknet_0_net450;
 wire clknet_1_0__leaf_net450;
 wire clknet_1_1__leaf_net450;
 wire clknet_0_net720;
 wire clknet_1_0__leaf_net720;
 wire clknet_1_1__leaf_net720;
 wire clknet_0_net354;
 wire clknet_1_0__leaf_net354;
 wire clknet_1_1__leaf_net354;
 wire clknet_0_net392;
 wire clknet_1_0__leaf_net392;
 wire clknet_1_1__leaf_net392;
 wire clknet_0_net386;
 wire clknet_1_0__leaf_net386;
 wire clknet_1_1__leaf_net386;
 wire clknet_0_net351;
 wire clknet_1_0__leaf_net351;
 wire clknet_1_1__leaf_net351;
 wire clknet_0_net719;
 wire clknet_1_0__leaf_net719;
 wire clknet_1_1__leaf_net719;
 wire clknet_0_net701;
 wire clknet_1_0__leaf_net701;
 wire clknet_1_1__leaf_net701;
 wire clknet_0_net385;
 wire clknet_1_0__leaf_net385;
 wire clknet_1_1__leaf_net385;
 wire clknet_0_net925;
 wire clknet_1_0__leaf_net925;
 wire clknet_1_1__leaf_net925;
 wire clknet_0_net301;
 wire clknet_1_0__leaf_net301;
 wire clknet_1_1__leaf_net301;
 wire clknet_0_net700;
 wire clknet_1_0__leaf_net700;
 wire clknet_1_1__leaf_net700;
 wire clknet_0_net275;
 wire clknet_1_0__leaf_net275;
 wire clknet_1_1__leaf_net275;
 wire clknet_0_net271;
 wire clknet_1_0__leaf_net271;
 wire clknet_1_1__leaf_net271;
 wire clknet_0_net305;
 wire clknet_1_0__leaf_net305;
 wire clknet_1_1__leaf_net305;
 wire clknet_0_net299;
 wire clknet_1_0__leaf_net299;
 wire clknet_1_1__leaf_net299;
 wire clknet_0_net917;
 wire clknet_1_0__leaf_net917;
 wire clknet_1_1__leaf_net917;
 wire clknet_0_net283;
 wire clknet_1_0__leaf_net283;
 wire clknet_1_1__leaf_net283;
 wire clknet_0_net277;
 wire clknet_1_0__leaf_net277;
 wire clknet_1_1__leaf_net277;
 wire clknet_0_net699;
 wire clknet_1_0__leaf_net699;
 wire clknet_1_1__leaf_net699;
 wire clknet_0_net269;
 wire clknet_1_0__leaf_net269;
 wire clknet_1_1__leaf_net269;
 wire clknet_0_net933;
 wire clknet_1_0__leaf_net933;
 wire clknet_1_1__leaf_net933;
 wire clknet_0_net288;
 wire clknet_1_0__leaf_net288;
 wire clknet_1_1__leaf_net288;
 wire clknet_0_net291;
 wire clknet_1_0__leaf_net291;
 wire clknet_1_1__leaf_net291;
 wire clknet_0_net220;
 wire clknet_1_0__leaf_net220;
 wire clknet_1_1__leaf_net220;
 wire clknet_0_net942;
 wire clknet_1_0__leaf_net942;
 wire clknet_1_1__leaf_net942;
 wire clknet_0_net226;
 wire clknet_1_0__leaf_net226;
 wire clknet_1_1__leaf_net226;
 wire clknet_0_net222;
 wire clknet_1_0__leaf_net222;
 wire clknet_1_1__leaf_net222;
 wire clknet_0_net208;
 wire clknet_1_0__leaf_net208;
 wire clknet_1_1__leaf_net208;
 wire clknet_0_net914;
 wire clknet_1_0__leaf_net914;
 wire clknet_1_1__leaf_net914;
 wire clknet_0_net328;
 wire clknet_1_0__leaf_net328;
 wire clknet_1_1__leaf_net328;
 wire clknet_0_net320;
 wire clknet_1_0__leaf_net320;
 wire clknet_1_1__leaf_net320;
 wire clknet_0_net216;
 wire clknet_1_0__leaf_net216;
 wire clknet_1_1__leaf_net216;
 wire clknet_0_net214;
 wire clknet_1_0__leaf_net214;
 wire clknet_1_1__leaf_net214;
 wire clknet_0_net922;
 wire clknet_1_0__leaf_net922;
 wire clknet_1_1__leaf_net922;
 wire clknet_0_net330;
 wire clknet_1_0__leaf_net330;
 wire clknet_1_1__leaf_net330;
 wire clknet_0_net331;
 wire clknet_1_0__leaf_net331;
 wire clknet_1_1__leaf_net331;
 wire clknet_0_net918;
 wire clknet_1_0__leaf_net918;
 wire clknet_1_1__leaf_net918;
 wire clknet_0_net902;
 wire clknet_1_0__leaf_net902;
 wire clknet_1_1__leaf_net902;
 wire clknet_0_net680;
 wire clknet_1_0__leaf_net680;
 wire clknet_1_1__leaf_net680;
 wire clknet_0_net907;
 wire clknet_1_0__leaf_net907;
 wire clknet_1_1__leaf_net907;
 wire clknet_0_net911;
 wire clknet_1_0__leaf_net911;
 wire clknet_1_1__leaf_net911;
 wire clknet_0_net938;
 wire clknet_1_0__leaf_net938;
 wire clknet_1_1__leaf_net938;
 wire clknet_0_net664;
 wire clknet_1_0__leaf_net664;
 wire clknet_1_1__leaf_net664;
 wire clknet_0_net105;
 wire clknet_1_0__leaf_net105;
 wire clknet_1_1__leaf_net105;
 wire clknet_0_net325;
 wire clknet_1_0__leaf_net325;
 wire clknet_1_1__leaf_net325;
 wire clknet_0_net218;
 wire clknet_1_0__leaf_net218;
 wire clknet_1_1__leaf_net218;
 wire clknet_0_net114;
 wire clknet_1_0__leaf_net114;
 wire clknet_1_1__leaf_net114;
 wire clknet_0_net111;
 wire clknet_1_0__leaf_net111;
 wire clknet_1_1__leaf_net111;
 wire clknet_0_net948;
 wire clknet_1_0__leaf_net948;
 wire clknet_1_1__leaf_net948;
 wire clknet_0_net952;
 wire clknet_1_0__leaf_net952;
 wire clknet_1_1__leaf_net952;
 wire clknet_0_net928;
 wire clknet_1_0__leaf_net928;
 wire clknet_1_1__leaf_net928;
 wire clknet_0_net927;
 wire clknet_1_0__leaf_net927;
 wire clknet_1_1__leaf_net927;
 wire clknet_0_net897;
 wire clknet_1_0__leaf_net897;
 wire clknet_1_1__leaf_net897;
 wire clknet_0_net110;
 wire clknet_1_0__leaf_net110;
 wire clknet_1_1__leaf_net110;
 wire clknet_0_net96;
 wire clknet_1_0__leaf_net96;
 wire clknet_1_1__leaf_net96;
 wire clknet_0_net315;
 wire clknet_1_0__leaf_net315;
 wire clknet_1_1__leaf_net315;
 wire clknet_0_net893;
 wire clknet_1_0__leaf_net893;
 wire clknet_1_1__leaf_net893;
 wire clknet_0_net412;
 wire clknet_1_0__leaf_net412;
 wire clknet_1_1__leaf_net412;
 wire clknet_0_net193;
 wire clknet_1_0__leaf_net193;
 wire clknet_1_1__leaf_net193;
 wire clknet_0_net99;
 wire clknet_1_0__leaf_net99;
 wire clknet_1_1__leaf_net99;
 wire clknet_0_net614;
 wire clknet_1_0__leaf_net614;
 wire clknet_1_1__leaf_net614;
 wire clknet_0_net190;
 wire clknet_1_0__leaf_net190;
 wire clknet_1_1__leaf_net190;
 wire clknet_0_net196;
 wire clknet_1_0__leaf_net196;
 wire clknet_1_1__leaf_net196;
 wire clknet_0_net919;
 wire clknet_1_0__leaf_net919;
 wire clknet_1_1__leaf_net919;
 wire clknet_0_net944;
 wire clknet_1_0__leaf_net944;
 wire clknet_1_1__leaf_net944;
 wire clknet_0_net199;
 wire clknet_1_0__leaf_net199;
 wire clknet_1_1__leaf_net199;
 wire clknet_0_net200;
 wire clknet_1_0__leaf_net200;
 wire clknet_1_1__leaf_net200;
 wire clknet_0_net100;
 wire clknet_1_0__leaf_net100;
 wire clknet_1_1__leaf_net100;
 wire clknet_0_net663;
 wire clknet_1_0__leaf_net663;
 wire clknet_1_1__leaf_net663;
 wire clknet_0_net931;
 wire clknet_1_0__leaf_net931;
 wire clknet_1_1__leaf_net931;
 wire clknet_0_net924;
 wire clknet_1_0__leaf_net924;
 wire clknet_1_1__leaf_net924;
 wire clknet_0_net646;
 wire clknet_1_0__leaf_net646;
 wire clknet_1_1__leaf_net646;
 wire clknet_0_net468;
 wire clknet_1_0__leaf_net468;
 wire clknet_1_1__leaf_net468;
 wire clknet_0_net474;
 wire clknet_1_0__leaf_net474;
 wire clknet_1_1__leaf_net474;
 wire clknet_0_net467;
 wire clknet_1_0__leaf_net467;
 wire clknet_1_1__leaf_net467;
 wire clknet_0_net462;
 wire clknet_1_0__leaf_net462;
 wire clknet_1_1__leaf_net462;
 wire clknet_0_net613;
 wire clknet_1_0__leaf_net613;
 wire clknet_1_1__leaf_net613;
 wire clknet_0_net189;
 wire clknet_1_0__leaf_net189;
 wire clknet_1_1__leaf_net189;
 wire clknet_0_net169;
 wire clknet_1_0__leaf_net169;
 wire clknet_1_1__leaf_net169;
 wire clknet_0_net198;
 wire clknet_1_0__leaf_net198;
 wire clknet_1_1__leaf_net198;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;

 sky130_fd_sc_hd__mux4_2 c100 (.A0(net876),
    .A1(net799),
    .A2(net870),
    .A3(net839),
    .S0(net849),
    .S1(net865),
    .X(net0));
 sky130_fd_sc_hd__mux4_2 c101 (.A0(net869),
    .A1(net1035),
    .A2(net1029),
    .A3(net876),
    .S0(net849),
    .S1(net872),
    .X(net1));
 sky130_fd_sc_hd__mux4_2 c102 (.A0(net862),
    .A1(net866),
    .A2(net849),
    .A3(net0),
    .S0(net875),
    .S1(net873),
    .X(net2));
 sky130_fd_sc_hd__mux4_2 c103 (.A0(net799),
    .A1(net858),
    .A2(net865),
    .A3(net866),
    .S0(net0),
    .S1(net876),
    .X(net912));
 sky130_fd_sc_hd__mux4_2 c104 (.A0(net853),
    .A1(net2),
    .A2(net877),
    .A3(net875),
    .S0(net855),
    .S1(net0),
    .X(net935));
 sky130_fd_sc_hd__mux4_2 c105 (.A0(net860),
    .A1(net822),
    .A2(net870),
    .A3(net843),
    .S0(net875),
    .S1(net876),
    .X(net3));
 sky130_fd_sc_hd__mux4_2 c106 (.A0(net877),
    .A1(net3),
    .A2(net869),
    .A3(net874),
    .S0(net871),
    .S1(net0),
    .X(net4));
 sky130_fd_sc_hd__mux4_1 c107 (.A0(net870),
    .A1(net868),
    .A2(net873),
    .A3(net820),
    .S0(net4),
    .S1(net1034),
    .X(net5));
 sky130_fd_sc_hd__mux4_2 c108 (.A0(net858),
    .A1(net4),
    .A2(net5),
    .A3(net3),
    .S0(net866),
    .S1(net1005),
    .X(net6));
 sky130_fd_sc_hd__mux4_2 c109 (.A0(net5),
    .A1(net1),
    .A2(net912),
    .A3(net874),
    .S0(net3),
    .S1(net849),
    .X(net7));
 sky130_fd_sc_hd__a2111o_1 c110 (.A1(net1),
    .A2(net848),
    .B1(net0),
    .C1(net3),
    .D1(net1005),
    .X(net953));
 sky130_fd_sc_hd__a2111o_1 c111 (.A1(net849),
    .A2(net871),
    .B1(net857),
    .C1(net7),
    .D1(net1034),
    .X(net905));
 sky130_fd_sc_hd__a2111o_4 c112 (.A1(net863),
    .A2(net871),
    .B1(net1032),
    .C1(net999),
    .D1(net912),
    .X(net8));
 sky130_fd_sc_hd__a2111o_1 c113 (.A1(net0),
    .A2(net999),
    .B1(net8),
    .C1(net852),
    .D1(net953),
    .X(net9));
 sky130_fd_sc_hd__a2111o_1 c114 (.A1(net2),
    .A2(net9),
    .B1(net8),
    .C1(net1),
    .D1(net999),
    .X(net10));
 sky130_fd_sc_hd__a2111o_4 c115 (.A1(net871),
    .A2(net854),
    .B1(net1),
    .C1(net2),
    .D1(net859),
    .X(net939));
 sky130_fd_sc_hd__a2111o_1 c116 (.A1(net10),
    .A2(net871),
    .B1(net999),
    .C1(net9),
    .D1(net8),
    .X(net11));
 sky130_fd_sc_hd__a2111o_1 c117 (.A1(net830),
    .A2(net793),
    .B1(net939),
    .C1(net2),
    .D1(net953),
    .X(net12));
 sky130_fd_sc_hd__a2111o_2 c118 (.A1(net12),
    .A2(net7),
    .B1(net2),
    .C1(net939),
    .D1(net833),
    .X(net941));
 sky130_fd_sc_hd__a2111o_1 c119 (.A1(net11),
    .A2(net8),
    .B1(net953),
    .C1(net849),
    .D1(net3),
    .X(net13));
 sky130_fd_sc_hd__mux4_1 c120 (.A0(net852),
    .A1(net999),
    .A2(net12),
    .A3(net3),
    .S0(net843),
    .S1(net833),
    .X(net14));
 sky130_fd_sc_hd__a2111o_1 c121 (.A1(net13),
    .A2(net941),
    .B1(net1005),
    .C1(net12),
    .D1(net939),
    .X(net946));
 sky130_fd_sc_hd__mux4_2 c122 (.A0(net9),
    .A1(net941),
    .A2(net946),
    .A3(net830),
    .S0(net8),
    .S1(net863),
    .X(net959));
 sky130_fd_sc_hd__a2111o_1 c123 (.A1(net11),
    .A2(net848),
    .B1(net959),
    .C1(net10),
    .D1(net939),
    .X(net15));
 sky130_fd_sc_hd__a2111o_2 c124 (.A1(net857),
    .A2(net941),
    .B1(net959),
    .C1(net999),
    .D1(net8),
    .X(net16));
 sky130_fd_sc_hd__a2111o_1 c125 (.A1(net15),
    .A2(net999),
    .B1(net2),
    .C1(net16),
    .D1(net1),
    .X(net17));
 sky130_fd_sc_hd__a2111o_1 c126 (.A1(net859),
    .A2(net848),
    .B1(net14),
    .C1(net16),
    .D1(net12),
    .X(net913));
 sky130_fd_sc_hd__mux4_1 c127 (.A0(net3),
    .A1(net16),
    .A2(net17),
    .A3(net939),
    .S0(net0),
    .S1(net913),
    .X(net18));
 sky130_fd_sc_hd__mux4_1 c128 (.A0(net17),
    .A1(net939),
    .A2(net854),
    .A3(net827),
    .S0(net848),
    .S1(net946),
    .X(net881));
 sky130_fd_sc_hd__a2111o_1 c129 (.A1(net18),
    .A2(net999),
    .B1(net16),
    .C1(net11),
    .D1(net8),
    .X(net949));
 sky130_fd_sc_hd__mux4_2 c130 (.A0(net14),
    .A1(net18),
    .A2(net949),
    .A3(net16),
    .S0(net793),
    .S1(net939),
    .X(net926));
 sky130_fd_sc_hd__a2111o_1 c131 (.A1(net949),
    .A2(net941),
    .B1(net926),
    .C1(net15),
    .D1(net939),
    .X(net932));
 sky130_fd_sc_hd__a2111o_4 c132 (.A1(net801),
    .A2(net790),
    .B1(net784),
    .C1(net786),
    .D1(net1024),
    .X(net19));
 sky130_fd_sc_hd__a2111o_1 c133 (.A1(net165),
    .A2(net1035),
    .B1(net1027),
    .C1(net782),
    .D1(net19),
    .X(net20));
 sky130_fd_sc_hd__a2111o_4 c134 (.A1(net1033),
    .A2(net1074),
    .B1(net1008),
    .C1(net791),
    .D1(net1027),
    .X(net21));
 sky130_fd_sc_hd__mux4_2 c135 (.A0(net1007),
    .A1(net786),
    .A2(net790),
    .A3(net834),
    .S0(net1035),
    .S1(net1027),
    .X(net22));
 sky130_fd_sc_hd__a2111o_4 c136 (.A1(net21),
    .A2(net1074),
    .B1(net1008),
    .C1(net1003),
    .D1(net19),
    .X(net23));
 sky130_fd_sc_hd__a2111o_2 c137 (.A1(net23),
    .A2(net1031),
    .B1(net1035),
    .C1(net1007),
    .D1(net1003),
    .X(net24));
 sky130_fd_sc_hd__a2111o_1 c138 (.A1(net781),
    .A2(net786),
    .B1(net845),
    .C1(net23),
    .D1(net21),
    .X(net929));
 sky130_fd_sc_hd__a2111o_1 c139 (.A1(net790),
    .A2(net1007),
    .B1(net788),
    .C1(net19),
    .D1(net23),
    .X(net25));
 sky130_fd_sc_hd__mux4_2 c140 (.A0(net786),
    .A1(net21),
    .A2(net1008),
    .A3(net1003),
    .S0(net1031),
    .S1(net997),
    .X(net26));
 sky130_fd_sc_hd__a2111o_1 c141 (.A1(net792),
    .A2(net24),
    .B1(net790),
    .C1(net1007),
    .D1(net23),
    .X(net27));
 sky130_fd_sc_hd__a2111o_4 c142 (.A1(net1008),
    .A2(net26),
    .B1(net997),
    .C1(net24),
    .D1(net1003),
    .X(net28));
 sky130_fd_sc_hd__a2111o_4 c143 (.A1(net19),
    .A2(net25),
    .B1(net790),
    .C1(net997),
    .D1(net1007),
    .X(net29));
 sky130_fd_sc_hd__mux4_2 c144 (.A0(net29),
    .A1(net27),
    .A2(net24),
    .A3(net1027),
    .S0(net1062),
    .S1(net28),
    .X(net910));
 sky130_fd_sc_hd__a2111o_1 c145 (.A1(net27),
    .A2(net790),
    .B1(net1062),
    .C1(net29),
    .D1(net992),
    .X(net30));
 sky130_fd_sc_hd__mux4_2 c146 (.A0(net25),
    .A1(net23),
    .A2(net29),
    .A3(net27),
    .S0(net26),
    .S1(net782),
    .X(net31));
 sky130_fd_sc_hd__mux4_2 c147 (.A0(net993),
    .A1(net24),
    .A2(net31),
    .A3(net1062),
    .S0(net29),
    .S1(net783),
    .X(net32));
 sky130_fd_sc_hd__mux4_1 c148 (.A0(net801),
    .A1(net25),
    .A2(net786),
    .A3(net1024),
    .S0(net1033),
    .S1(net845),
    .X(net33));
 sky130_fd_sc_hd__mux4_2 c149 (.A0(net30),
    .A1(net29),
    .A2(net31),
    .A3(net995),
    .S0(net21),
    .S1(net993),
    .X(net34));
 sky130_fd_sc_hd__mux4_2 c150 (.A0(net34),
    .A1(net32),
    .A2(net1062),
    .A3(net790),
    .S0(net31),
    .S1(net995),
    .X(net35));
 sky130_fd_sc_hd__mux4_2 c151 (.A0(net31),
    .A1(net792),
    .A2(net25),
    .A3(net34),
    .S0(net1033),
    .S1(net30),
    .X(net36));
 sky130_fd_sc_hd__mux4_2 c152 (.A0(net36),
    .A1(net32),
    .A2(net27),
    .A3(net35),
    .S0(net34),
    .S1(net1062),
    .X(net37));
 sky130_fd_sc_hd__mux4_2 c153 (.A0(net834),
    .A1(net28),
    .A2(net36),
    .A3(net35),
    .S0(net786),
    .S1(net29),
    .X(net38));
 sky130_fd_sc_hd__a2111o_1 c154 (.A1(net465),
    .A2(net24),
    .B1(net811),
    .C1(net1031),
    .D1(net784),
    .X(net39));
 sky130_fd_sc_hd__a2111o_4 c155 (.A1(net39),
    .A2(net802),
    .B1(net19),
    .C1(net795),
    .D1(net793),
    .X(net40));
 sky130_fd_sc_hd__a2111o_4 c156 (.A1(net40),
    .A2(net805),
    .B1(net1003),
    .C1(net810),
    .D1(net1027),
    .X(net41));
 sky130_fd_sc_hd__a2111o_1 c157 (.A1(net1039),
    .A2(net809),
    .B1(net40),
    .C1(net995),
    .D1(net1038),
    .X(net42));
 sky130_fd_sc_hd__a2111o_4 c158 (.A1(net37),
    .A2(net40),
    .B1(net804),
    .C1(net813),
    .D1(net1027),
    .X(net43));
 sky130_fd_sc_hd__mux4_1 c159 (.A0(net795),
    .A1(net1034),
    .A2(net805),
    .A3(net40),
    .S0(net793),
    .S1(net990),
    .X(net44));
 sky130_fd_sc_hd__mux4_2 c160 (.A0(net806),
    .A1(net43),
    .A2(net41),
    .A3(net44),
    .S0(net811),
    .S1(net990),
    .X(net45));
 sky130_fd_sc_hd__a2111o_4 c161 (.A1(net797),
    .A2(net808),
    .B1(net800),
    .C1(net41),
    .D1(net793),
    .X(net46));
 sky130_fd_sc_hd__mux4_1 c162 (.A0(net43),
    .A1(net1039),
    .A2(net45),
    .A3(net813),
    .S0(net797),
    .S1(net990),
    .X(net47));
 sky130_fd_sc_hd__mux4_2 c163 (.A0(net45),
    .A1(net1074),
    .A2(net39),
    .A3(net40),
    .S0(net43),
    .S1(net990),
    .X(net48));
 sky130_fd_sc_hd__mux4_2 c164 (.A0(net44),
    .A1(net1034),
    .A2(net816),
    .A3(net46),
    .S0(net1063),
    .S1(net986),
    .X(net49));
 sky130_fd_sc_hd__mux4_2 c165 (.A0(net783),
    .A1(net35),
    .A2(net47),
    .A3(net46),
    .S0(net49),
    .S1(net986),
    .X(net50));
 sky130_fd_sc_hd__mux4_2 c166 (.A0(net784),
    .A1(net813),
    .A2(net986),
    .A3(net1039),
    .S0(net40),
    .S1(net49),
    .X(net51));
 sky130_fd_sc_hd__mux4_2 c167 (.A0(net32),
    .A1(net809),
    .A2(net811),
    .A3(net1034),
    .S0(net51),
    .S1(net40),
    .X(net52));
 sky130_fd_sc_hd__mux4_2 c168 (.A0(net47),
    .A1(net1027),
    .A2(net32),
    .A3(net51),
    .S0(net991),
    .S1(net50),
    .X(net53));
 sky130_fd_sc_hd__mux4_1 c169 (.A0(net49),
    .A1(net45),
    .A2(net40),
    .A3(net990),
    .S0(net806),
    .S1(net51),
    .X(net54));
 sky130_fd_sc_hd__mux4_1 c170 (.A0(net51),
    .A1(net39),
    .A2(net47),
    .A3(net796),
    .S0(net45),
    .S1(net973),
    .X(net55));
 sky130_fd_sc_hd__mux4_2 c171 (.A0(net1033),
    .A1(net49),
    .A2(net47),
    .A3(net808),
    .S0(net995),
    .S1(net50),
    .X(net56));
 sky130_fd_sc_hd__mux4_2 c172 (.A0(net800),
    .A1(net52),
    .A2(net56),
    .A3(net41),
    .S0(net804),
    .S1(net465),
    .X(net57));
 sky130_fd_sc_hd__mux4_2 c173 (.A0(net50),
    .A1(net56),
    .A2(net57),
    .A3(net52),
    .S0(net41),
    .S1(net51),
    .X(net58));
 sky130_fd_sc_hd__mux4_1 c174 (.A0(net1031),
    .A1(net50),
    .A2(net31),
    .A3(net39),
    .S0(net58),
    .S1(net56),
    .X(net59));
 sky130_fd_sc_hd__mux4_1 c175 (.A0(net59),
    .A1(net55),
    .A2(net51),
    .A3(net58),
    .S0(net43),
    .S1(net56),
    .X(net60));
 sky130_fd_sc_hd__a2111o_4 c176 (.A1(net828),
    .A2(net826),
    .B1(net813),
    .C1(net832),
    .D1(net616),
    .X(net957));
 sky130_fd_sc_hd__a2111o_1 c177 (.A1(net798),
    .A2(net1038),
    .B1(net817),
    .C1(net820),
    .D1(net31),
    .X(net61));
 sky130_fd_sc_hd__a2111o_1 c178 (.A1(net821),
    .A2(net48),
    .B1(net990),
    .C1(net837),
    .D1(net798),
    .X(net62));
 sky130_fd_sc_hd__mux4_2 c179 (.A0(net24),
    .A1(net803),
    .A2(net833),
    .A3(net839),
    .S0(net828),
    .S1(net616),
    .X(net63));
 sky130_fd_sc_hd__mux4_2 c180 (.A0(net57),
    .A1(net31),
    .A2(net820),
    .A3(net827),
    .S0(net826),
    .S1(net61),
    .X(net943));
 sky130_fd_sc_hd__mux4_2 c181 (.A0(net821),
    .A1(net810),
    .A2(net787),
    .A3(net813),
    .S0(net46),
    .S1(net616),
    .X(net64));
 sky130_fd_sc_hd__mux4_2 c182 (.A0(net803),
    .A1(net943),
    .A2(net826),
    .A3(net827),
    .S0(net990),
    .S1(net840),
    .X(net940));
 sky130_fd_sc_hd__mux4_2 c183 (.A0(net836),
    .A1(net63),
    .A2(net821),
    .A3(net64),
    .S0(net819),
    .S1(net810),
    .X(net65));
 sky130_fd_sc_hd__mux4_2 c184 (.A0(net62),
    .A1(net31),
    .A2(net839),
    .A3(net989),
    .S0(net943),
    .S1(net58),
    .X(net66));
 sky130_fd_sc_hd__mux4_1 c185 (.A0(net58),
    .A1(net940),
    .A2(net31),
    .A3(net832),
    .S0(net64),
    .S1(net616),
    .X(net67));
 sky130_fd_sc_hd__sdfbbn_2 c186 (.CLK_N(clknet_4_4_0_clk),
    .D(net1035),
    .RESET_B(net837),
    .SCD(net940),
    .SCE(net989),
    .SET_B(net656),
    .Q(net69),
    .Q_N(net68));
 sky130_fd_sc_hd__mux4_2 c187 (.A0(net64),
    .A1(net1038),
    .A2(net943),
    .A3(net838),
    .S0(net989),
    .S1(net657),
    .X(net70));
 sky130_fd_sc_hd__mux4_1 c188 (.A0(net840),
    .A1(net1063),
    .A2(net839),
    .A3(net940),
    .S0(net68),
    .S1(net943),
    .X(net71));
 sky130_fd_sc_hd__mux4_1 c189 (.A0(net1038),
    .A1(net803),
    .A2(net70),
    .A3(net989),
    .S0(net66),
    .S1(net68),
    .X(net72));
 sky130_fd_sc_hd__mux4_2 c190 (.A0(net943),
    .A1(net989),
    .A2(net68),
    .A3(net62),
    .S0(net616),
    .S1(net656),
    .X(net73));
 sky130_fd_sc_hd__mux4_2 c191 (.A0(net831),
    .A1(net989),
    .A2(net793),
    .A3(net46),
    .S0(net599),
    .S1(net657),
    .X(net74));
 sky130_fd_sc_hd__mux4_1 c192 (.A0(net63),
    .A1(net74),
    .A2(net1074),
    .A3(net827),
    .S0(net989),
    .S1(net968),
    .X(net75));
 sky130_fd_sc_hd__a2111o_1 c193 (.A1(net74),
    .A2(net70),
    .B1(net599),
    .C1(net656),
    .D1(net659),
    .X(net76));
 sky130_fd_sc_hd__mux4_1 c194 (.A0(net831),
    .A1(net74),
    .A2(net968),
    .A3(net793),
    .S0(net839),
    .S1(net1066),
    .X(net77));
 sky130_fd_sc_hd__mux4_1 c195 (.A0(net995),
    .A1(net989),
    .A2(net74),
    .A3(net68),
    .S0(net66),
    .S1(net615),
    .X(net78));
 sky130_fd_sc_hd__mux4_1 c196 (.A0(net940),
    .A1(net58),
    .A2(net74),
    .A3(net57),
    .S0(net968),
    .S1(net660),
    .X(net79));
 sky130_fd_sc_hd__mux4_1 c197 (.A0(net61),
    .A1(net70),
    .A2(net968),
    .A3(net615),
    .S0(net660),
    .S1(net661),
    .X(net80));
 sky130_fd_sc_hd__mux4_2 c198 (.A0(net851),
    .A1(net69),
    .A2(net854),
    .A3(net1074),
    .S0(net864),
    .S1(net846),
    .X(net81));
 sky130_fd_sc_hd__mux4_2 c199 (.A0(net847),
    .A1(net81),
    .A2(net63),
    .A3(net997),
    .S0(net864),
    .S1(net1070),
    .X(net82));
 sky130_fd_sc_hd__mux4_1 c200 (.A0(net81),
    .A1(net864),
    .A2(net839),
    .A3(net82),
    .S0(net985),
    .S1(net940),
    .X(net83));
 sky130_fd_sc_hd__mux4_2 c201 (.A0(net844),
    .A1(net63),
    .A2(net81),
    .A3(net787),
    .S0(net817),
    .S1(net854),
    .X(net84));
 sky130_fd_sc_hd__mux4_2 c202 (.A0(net84),
    .A1(net985),
    .A2(net817),
    .A3(net808),
    .S0(net81),
    .S1(net835),
    .X(net85));
 sky130_fd_sc_hd__mux4_2 c203 (.A0(net787),
    .A1(net817),
    .A2(net796),
    .A3(net85),
    .S0(net985),
    .S1(net81),
    .X(net86));
 sky130_fd_sc_hd__mux4_2 c204 (.A0(net86),
    .A1(net85),
    .A2(net63),
    .A3(net985),
    .S0(net864),
    .S1(net81),
    .X(net87));
 sky130_fd_sc_hd__mux4_2 c205 (.A0(net87),
    .A1(net86),
    .A2(net820),
    .A3(net85),
    .S0(net854),
    .S1(net661),
    .X(net88));
 sky130_fd_sc_hd__mux4_2 c206 (.A0(net835),
    .A1(net82),
    .A2(net88),
    .A3(net87),
    .S0(net861),
    .S1(net659),
    .X(net89));
 sky130_fd_sc_hd__mux4_1 c207 (.A0(net819),
    .A1(net854),
    .A2(net968),
    .A3(net89),
    .S0(net82),
    .S1(net1070),
    .X(net90));
 sky130_fd_sc_hd__mux4_2 c208 (.A0(net861),
    .A1(net989),
    .A2(net89),
    .A3(net841),
    .S0(net864),
    .S1(net84),
    .X(net91));
 sky130_fd_sc_hd__mux4_1 c209 (.A0(net85),
    .A1(net968),
    .A2(net864),
    .A3(net848),
    .S0(net837),
    .S1(net86),
    .X(net92));
 sky130_fd_sc_hd__mux4_1 c210 (.A0(net1074),
    .A1(net849),
    .A2(net87),
    .A3(net86),
    .S0(net88),
    .S1(net91),
    .X(net93));
 sky130_fd_sc_hd__mux4_1 c211 (.A0(net89),
    .A1(net81),
    .A2(net86),
    .A3(net88),
    .S0(clknet_1_0__leaf_net924),
    .S1(clknet_1_1__leaf_net663),
    .X(net931));
 sky130_fd_sc_hd__mux4_1 c212 (.A0(net837),
    .A1(net88),
    .A2(clknet_1_1__leaf_net931),
    .A3(net968),
    .S0(net91),
    .S1(clknet_1_0__leaf_net663),
    .X(net94));
 sky130_fd_sc_hd__mux4_1 c213 (.A0(net91),
    .A1(clknet_1_1__leaf_net931),
    .A2(net84),
    .A3(net854),
    .S0(net87),
    .S1(clknet_1_0__leaf_net663),
    .X(net95));
 sky130_fd_sc_hd__mux4_1 c214 (.A0(net850),
    .A1(net86),
    .A2(net82),
    .A3(net957),
    .S0(net598),
    .S1(clknet_1_1__leaf_net664),
    .X(net96));
 sky130_fd_sc_hd__mux4_1 c215 (.A0(net88),
    .A1(net91),
    .A2(net82),
    .A3(net854),
    .S0(clknet_1_0__leaf_net663),
    .S1(clknet_1_1__leaf_net664),
    .X(net97));
 sky130_fd_sc_hd__mux4_1 c216 (.A0(net1042),
    .A1(net84),
    .A2(net957),
    .A3(net968),
    .S0(net934),
    .S1(net630),
    .X(net98));
 sky130_fd_sc_hd__mux4_1 c217 (.A0(net826),
    .A1(net84),
    .A2(clknet_1_0__leaf_net96),
    .A3(net630),
    .S0(clknet_1_1__leaf_net663),
    .S1(net666),
    .X(net99));
 sky130_fd_sc_hd__mux4_1 c218 (.A0(net817),
    .A1(net1042),
    .A2(clknet_1_1__leaf_net99),
    .A3(net630),
    .S0(clknet_1_1__leaf_net663),
    .S1(net666),
    .X(net100));
 sky130_fd_sc_hd__mux4_1 c219 (.A0(net957),
    .A1(clknet_1_1__leaf_net99),
    .A2(clknet_1_1__leaf_net931),
    .A3(clknet_1_0__leaf_net96),
    .S0(net630),
    .S1(net666),
    .X(net101));
 sky130_fd_sc_hd__a2111o_1 c220 (.A1(net82),
    .A2(net876),
    .B1(net818),
    .C1(net865),
    .D1(net810),
    .X(net102));
 sky130_fd_sc_hd__mux4_2 c221 (.A0(net810),
    .A1(net875),
    .A2(net957),
    .A3(net874),
    .S0(net820),
    .S1(net598),
    .X(net103));
 sky130_fd_sc_hd__mux4_2 c222 (.A0(net818),
    .A1(net103),
    .A2(net846),
    .A3(net1031),
    .S0(net876),
    .S1(net865),
    .X(net895));
 sky130_fd_sc_hd__mux4_1 c223 (.A0(net103),
    .A1(net843),
    .A2(net793),
    .A3(net1001),
    .S0(net957),
    .S1(clknet_1_1__leaf_net664),
    .X(net897));
 sky130_fd_sc_hd__mux4_1 c224 (.A0(net832),
    .A1(net940),
    .A2(net846),
    .A3(net1033),
    .S0(clknet_1_0__leaf_net931),
    .S1(net1001),
    .X(net104));
 sky130_fd_sc_hd__a2111o_1 c225 (.A1(net846),
    .A2(clknet_1_0__leaf_net897),
    .B1(net973),
    .C1(net572),
    .D1(clknet_1_0__leaf_net664),
    .X(net105));
 sky130_fd_sc_hd__mux4_1 c226 (.A0(clknet_1_0__leaf_net105),
    .A1(net6),
    .A2(net103),
    .A3(net1034),
    .S0(net937),
    .S1(clknet_1_0__leaf_net924),
    .X(net952));
 sky130_fd_sc_hd__a2111o_1 c227 (.A1(net875),
    .A2(clknet_1_0__leaf_net897),
    .B1(net89),
    .C1(clknet_1_0__leaf_net952),
    .D1(net7),
    .X(net927));
 sky130_fd_sc_hd__sdfbbn_1 c228 (.CLK_N(clknet_4_0_0_clk),
    .D(net63),
    .RESET_B(net1001),
    .SCD(net1054),
    .SCE(clknet_1_0__leaf_net927),
    .SET_B(net957),
    .Q(net107),
    .Q_N(net106));
 sky130_fd_sc_hd__a2111o_1 c229 (.A1(net107),
    .A2(clknet_1_0__leaf_net897),
    .B1(net846),
    .C1(clknet_1_0__leaf_net927),
    .D1(net912),
    .X(net108));
 sky130_fd_sc_hd__a2111o_1 c230 (.A1(net107),
    .A2(clknet_1_0__leaf_net927),
    .B1(net103),
    .C1(clknet_1_0__leaf_net897),
    .D1(net82),
    .X(net109));
 sky130_fd_sc_hd__mux4_1 c231 (.A0(clknet_1_0__leaf_net99),
    .A1(clknet_1_0__leaf_net897),
    .A2(net1001),
    .A3(net855),
    .S0(net937),
    .S1(net934),
    .X(net110));
 sky130_fd_sc_hd__a2111o_1 c232 (.A1(net5),
    .A2(clknet_1_0__leaf_net105),
    .B1(net868),
    .C1(net1032),
    .D1(clknet_1_0__leaf_net897),
    .X(net111));
 sky130_fd_sc_hd__a2111o_1 c233 (.A1(net102),
    .A2(clknet_1_0__leaf_net110),
    .B1(clknet_1_1__leaf_net927),
    .C1(net106),
    .D1(net954),
    .X(net112));
 sky130_fd_sc_hd__a2111o_1 c234 (.A1(net868),
    .A2(net1054),
    .B1(clknet_1_0__leaf_net952),
    .C1(clknet_1_0__leaf_net927),
    .D1(net63),
    .X(net113));
 sky130_fd_sc_hd__a2111o_2 c235 (.A1(net873),
    .A2(net985),
    .B1(net793),
    .C1(net63),
    .D1(net598),
    .X(net936));
 sky130_fd_sc_hd__a2111o_1 c236 (.A1(net936),
    .A2(clknet_1_0__leaf_net100),
    .B1(net1005),
    .C1(clknet_1_0__leaf_net105),
    .D1(net937),
    .X(net114));
 sky130_fd_sc_hd__sdfbbp_1 c237 (.CLK(clknet_4_0_0_clk),
    .D(net866),
    .RESET_B(clknet_1_0__leaf_net927),
    .SCD(net106),
    .SCE(clknet_1_1__leaf_net952),
    .SET_B(net647),
    .Q(net116),
    .Q_N(net115));
 sky130_fd_sc_hd__a2111o_1 c238 (.A1(clknet_1_1__leaf_net114),
    .A2(net866),
    .B1(net115),
    .C1(net936),
    .D1(clknet_1_0__leaf_net664),
    .X(net117));
 sky130_fd_sc_hd__or4bb_1 c239 (.A(clknet_1_1__leaf_net952),
    .B(net106),
    .C_N(net954),
    .D_N(clknet_1_1__leaf_net924),
    .X(net928));
 sky130_fd_sc_hd__mux4_1 c240 (.A0(net115),
    .A1(clknet_1_1__leaf_net952),
    .A2(clknet_1_0__leaf_net927),
    .A3(net954),
    .S0(net647),
    .S1(clknet_1_0__leaf_net924),
    .X(net118));
 sky130_fd_sc_hd__a2111o_1 c241 (.A1(net839),
    .A2(clknet_1_0__leaf_net111),
    .B1(clknet_1_0__leaf_net952),
    .C1(net115),
    .D1(net956),
    .X(net948));
 sky130_fd_sc_hd__mux4_1 c256 (.A0(net838),
    .A1(net13),
    .A2(net107),
    .A3(net953),
    .S0(clknet_1_0__leaf_net948),
    .S1(net1034),
    .X(net119));
 sky130_fd_sc_hd__mux4_2 c257 (.A0(net89),
    .A1(net16),
    .A2(net881),
    .A3(net939),
    .S0(net905),
    .S1(net912),
    .X(net958));
 sky130_fd_sc_hd__mux4_1 c258 (.A0(net941),
    .A1(net943),
    .A2(clknet_1_0__leaf_net114),
    .A3(net958),
    .S0(net572),
    .S1(net1069),
    .X(net120));
 sky130_fd_sc_hd__mux4_1 c259 (.A0(net958),
    .A1(net999),
    .A2(net874),
    .A3(net1046),
    .S0(net843),
    .S1(net1069),
    .X(net121));
 sky130_fd_sc_hd__mux4_1 c260 (.A0(net7),
    .A1(clknet_1_0__leaf_net952),
    .A2(net926),
    .A3(net958),
    .S0(net8),
    .S1(net951),
    .X(net122));
 sky130_fd_sc_hd__mux4_1 c261 (.A0(net874),
    .A1(net872),
    .A2(net958),
    .A3(net582),
    .S0(net954),
    .X(net123));
 sky130_fd_sc_hd__a2111o_1 c262 (.A1(clknet_1_0__leaf_net114),
    .A2(net1034),
    .B1(net959),
    .D1(net960),
    .X(net124));
 sky130_fd_sc_hd__mux4_1 c263 (.A0(net8),
    .A1(net820),
    .A2(net4),
    .A3(net957),
    .S0(net955),
    .S1(net960),
    .X(net901));
 sky130_fd_sc_hd__a2111o_1 c264 (.A1(net30),
    .A2(net29),
    .B1(net36),
    .C1(net993),
    .D1(net812),
    .X(net125));
 sky130_fd_sc_hd__a2111o_2 c265 (.A1(net791),
    .A2(net996),
    .B1(net21),
    .C1(net845),
    .D1(net993),
    .X(net126));
 sky130_fd_sc_hd__a2111o_1 c266 (.A1(net38),
    .A2(net30),
    .B1(net845),
    .C1(net1033),
    .D1(net126),
    .X(net127));
 sky130_fd_sc_hd__a2111o_4 c267 (.A1(net988),
    .A2(net26),
    .B1(net1035),
    .C1(net35),
    .D1(net165),
    .X(net128));
 sky130_fd_sc_hd__a2111o_4 c268 (.A1(net782),
    .A2(net34),
    .B1(net1035),
    .C1(net128),
    .D1(net988),
    .X(net129));
 sky130_fd_sc_hd__a2111o_1 c269 (.A1(net34),
    .A2(net126),
    .B1(net988),
    .C1(net995),
    .D1(net128),
    .X(net130));
 sky130_fd_sc_hd__a2111o_1 c270 (.A1(net988),
    .A2(net128),
    .B1(net983),
    .C1(net129),
    .D1(net1074),
    .X(net131));
 sky130_fd_sc_hd__a2111o_1 c271 (.A1(net28),
    .A2(net125),
    .B1(net129),
    .C1(net988),
    .D1(net983),
    .X(net132));
 sky130_fd_sc_hd__a2111o_4 c272 (.A1(net125),
    .A2(net983),
    .B1(net812),
    .C1(net981),
    .D1(net845),
    .X(net133));
 sky130_fd_sc_hd__a2111o_1 c273 (.A1(net128),
    .A2(net981),
    .B1(net38),
    .C1(net983),
    .D1(net133),
    .X(net134));
 sky130_fd_sc_hd__mux4_2 c274 (.A0(net984),
    .A1(net791),
    .A2(net134),
    .A3(net125),
    .S0(net981),
    .S1(net1028),
    .X(net135));
 sky130_fd_sc_hd__a2111o_1 c275 (.A1(net129),
    .A2(net983),
    .B1(net135),
    .C1(net981),
    .D1(net1047),
    .X(net136));
 sky130_fd_sc_hd__mux4_2 c276 (.A0(net131),
    .A1(net26),
    .A2(net136),
    .A3(net133),
    .S0(net1065),
    .S1(net1061),
    .X(net137));
 sky130_fd_sc_hd__sdfbbn_2 c277 (.CLK_N(clknet_4_7_0_clk),
    .D(net134),
    .RESET_B(net137),
    .SCD(net1052),
    .SCE(net984),
    .SET_B(net1060),
    .Q(net139),
    .Q_N(net138));
 sky130_fd_sc_hd__mux4_2 c278 (.A0(net37),
    .A1(net133),
    .A2(net136),
    .A3(net134),
    .S0(net1061),
    .S1(net1059),
    .X(net140));
 sky130_fd_sc_hd__mux4_2 c279 (.A0(net128),
    .A1(net135),
    .A2(net134),
    .A3(net136),
    .S0(net1057),
    .S1(net138),
    .X(net141));
 sky130_fd_sc_hd__mux4_1 c280 (.A0(net139),
    .A1(net135),
    .A2(net137),
    .A3(net1047),
    .S0(net1061),
    .S1(net1033),
    .X(net142));
 sky130_fd_sc_hd__mux4_1 c281 (.A0(net136),
    .A1(net141),
    .A2(net137),
    .A3(net1058),
    .S0(net1061),
    .S1(net573),
    .X(net143));
 sky130_fd_sc_hd__mux4_1 c282 (.A0(net137),
    .A1(net1047),
    .A2(net131),
    .A3(net129),
    .S0(net981),
    .S1(net1061),
    .X(net144));
 sky130_fd_sc_hd__sdfbbn_2 c283 (.CLK_N(clknet_4_7_0_clk),
    .D(net140),
    .RESET_B(net133),
    .SCD(net128),
    .SCE(net573),
    .SET_B(net1022),
    .Q(net146),
    .Q_N(net145));
 sky130_fd_sc_hd__mux4_2 c284 (.A0(net133),
    .A1(net139),
    .A2(net28),
    .A3(net129),
    .S0(net146),
    .S1(net573),
    .X(net147));
 sky130_fd_sc_hd__mux4_2 c285 (.A0(net126),
    .A1(net146),
    .A2(net38),
    .A3(net125),
    .S0(net1047),
    .S1(net573),
    .X(net148));
 sky130_fd_sc_hd__a2111o_1 c286 (.A1(net991),
    .A2(net37),
    .B1(net811),
    .C1(net802),
    .D1(net573),
    .X(net149));
 sky130_fd_sc_hd__a2111o_1 c287 (.A1(net805),
    .A2(net986),
    .B1(net149),
    .C1(net1074),
    .D1(net573),
    .X(net150));
 sky130_fd_sc_hd__a2111o_1 c288 (.A1(net804),
    .A2(net811),
    .B1(net979),
    .C1(net1074),
    .D1(net982),
    .X(net151));
 sky130_fd_sc_hd__a2111o_1 c289 (.A1(net41),
    .A2(net129),
    .B1(net979),
    .C1(net987),
    .D1(net573),
    .X(net152));
 sky130_fd_sc_hd__mux4_2 c290 (.A0(net151),
    .A1(net149),
    .A2(net41),
    .A3(net984),
    .S0(net129),
    .S1(net1031),
    .X(net921));
 sky130_fd_sc_hd__a2111o_1 c291 (.A1(net987),
    .A2(net990),
    .B1(net54),
    .C1(net971),
    .D1(net573),
    .X(net153));
 sky130_fd_sc_hd__mux4_2 c292 (.A0(net1027),
    .A1(net811),
    .A2(net57),
    .A3(net995),
    .S0(net979),
    .S1(net41),
    .X(net154));
 sky130_fd_sc_hd__a2111o_1 c293 (.A1(net982),
    .A2(net37),
    .B1(net1031),
    .C1(net984),
    .D1(net1027),
    .X(net155));
 sky130_fd_sc_hd__a2111o_1 c294 (.A1(net155),
    .A2(net154),
    .B1(net987),
    .C1(net971),
    .D1(net979),
    .X(net156));
 sky130_fd_sc_hd__a2111o_1 c295 (.A1(net155),
    .A2(net41),
    .B1(net154),
    .C1(net802),
    .D1(net987),
    .X(net157));
 sky130_fd_sc_hd__a2111o_1 c296 (.A1(net149),
    .A2(net1078),
    .B1(net156),
    .C1(net984),
    .D1(net995),
    .X(net158));
 sky130_fd_sc_hd__mux4_2 c297 (.A0(net153),
    .A1(net129),
    .A2(net993),
    .A3(net971),
    .S0(net979),
    .S1(net987),
    .X(net159));
 sky130_fd_sc_hd__a2111o_4 c298 (.A1(net979),
    .A2(net152),
    .B1(net159),
    .C1(net154),
    .D1(net973),
    .X(net880));
 sky130_fd_sc_hd__a2111o_4 c299 (.A1(net796),
    .A2(net152),
    .B1(net987),
    .C1(net979),
    .D1(net159),
    .X(net160));
 sky130_fd_sc_hd__sdfbbp_1 c300 (.CLK(clknet_4_5_0_clk),
    .D(net54),
    .RESET_B(net153),
    .SCD(net154),
    .SCE(net966),
    .SET_B(net987),
    .Q(net162),
    .Q_N(net161));
 sky130_fd_sc_hd__mux4_1 c301 (.A0(net162),
    .A1(net966),
    .A2(net151),
    .A3(net46),
    .S0(net1078),
    .S1(net967),
    .X(net163));
 sky130_fd_sc_hd__a2111o_1 c302 (.A1(net967),
    .A2(net151),
    .B1(net808),
    .C1(net971),
    .D1(net566),
    .X(net164));
 sky130_fd_sc_hd__mux4_2 c303 (.A0(net812),
    .A1(net155),
    .A2(net966),
    .A3(net161),
    .S0(net987),
    .X(net586));
 sky130_fd_sc_hd__mux4_1 c304 (.A0(net153),
    .A1(net46),
    .A2(net966),
    .A3(net161),
    .S0(net37),
    .S1(net586),
    .X(net166));
 sky130_fd_sc_hd__mux4_1 c305 (.A0(net157),
    .A1(net41),
    .A2(net979),
    .A3(net987),
    .S0(net585),
    .S1(net668),
    .X(net167));
 sky130_fd_sc_hd__mux4_1 c306 (.A0(net966),
    .A1(net1048),
    .A2(net987),
    .A3(net1033),
    .S0(net566),
    .S1(clknet_1_1__leaf_net613),
    .X(net168));
 sky130_fd_sc_hd__mux4_2 c307 (.A0(net997),
    .A1(net566),
    .A2(net586),
    .A3(clknet_1_1__leaf_net613),
    .S0(net668),
    .S1(net669),
    .X(net169));
 sky130_fd_sc_hd__mux4_2 c308 (.A0(net990),
    .A1(net827),
    .A2(net161),
    .A3(net986),
    .S0(net662),
    .S1(net669),
    .X(net170));
 sky130_fd_sc_hd__mux4_1 c309 (.A0(net152),
    .A1(net1042),
    .A2(net66),
    .A3(net1073),
    .S0(net1068),
    .S1(net669),
    .X(net171));
 sky130_fd_sc_hd__mux4_1 c310 (.A0(net46),
    .A1(net159),
    .A2(net138),
    .A3(net986),
    .S0(net661),
    .S1(net662),
    .X(net172));
 sky130_fd_sc_hd__mux4_1 c311 (.A0(net810),
    .A1(net162),
    .A2(net993),
    .A3(net660),
    .S0(net661),
    .S1(net662),
    .X(net173));
 sky130_fd_sc_hd__mux4_1 c312 (.A0(net129),
    .A1(net1029),
    .A2(net829),
    .A3(net986),
    .S0(net947),
    .S1(net669),
    .X(net174));
 sky130_fd_sc_hd__mux4_1 c313 (.A0(net159),
    .A1(net174),
    .A2(net978),
    .A3(net967),
    .S0(net986),
    .S1(net660),
    .X(net175));
 sky130_fd_sc_hd__mux4_1 c314 (.A0(net814),
    .A1(net810),
    .A2(net66),
    .A3(net660),
    .S0(net898),
    .S1(net1020),
    .X(net176));
 sky130_fd_sc_hd__mux4_1 c315 (.A0(net156),
    .A1(net829),
    .A2(net989),
    .A3(net947),
    .S0(net1020),
    .S1(net671),
    .X(net177));
 sky130_fd_sc_hd__mux4_1 c316 (.A0(net814),
    .A1(net70),
    .A2(net973),
    .A3(net662),
    .S0(net669),
    .S1(net672),
    .X(net178));
 sky130_fd_sc_hd__mux4_2 c317 (.A0(net174),
    .A1(net46),
    .A2(net669),
    .A3(net1020),
    .S0(net1019),
    .S1(net1017),
    .X(net179));
 sky130_fd_sc_hd__mux4_1 c318 (.A0(net156),
    .A1(net1029),
    .A2(net1064),
    .A3(net599),
    .S0(net1020),
    .S1(net671),
    .X(net180));
 sky130_fd_sc_hd__mux4_1 c319 (.A0(net66),
    .A1(net173),
    .A2(net978),
    .A3(net1035),
    .S0(net662),
    .S1(net672),
    .X(net181));
 sky130_fd_sc_hd__mux4_2 c320 (.A0(net173),
    .A1(net174),
    .A2(net990),
    .A3(net1020),
    .S0(net672),
    .S1(net1017),
    .X(net182));
 sky130_fd_sc_hd__mux4_1 c321 (.A0(net70),
    .A1(net46),
    .A2(clknet_1_0__leaf_net613),
    .A3(clknet_1_0__leaf_net614),
    .S0(net1019),
    .S1(net1017),
    .X(net183));
 sky130_fd_sc_hd__mux4_1 c322 (.A0(net70),
    .A1(net829),
    .A2(net573),
    .A3(net671),
    .S0(net1019),
    .S1(net1017),
    .X(net184));
 sky130_fd_sc_hd__mux4_1 c323 (.A0(net172),
    .A1(net956),
    .A2(clknet_1_0__leaf_net614),
    .A3(net1020),
    .S0(net671),
    .S1(net672),
    .X(net185));
 sky130_fd_sc_hd__mux4_2 c324 (.A0(net182),
    .A1(net1029),
    .A2(net630),
    .A3(net650),
    .S0(net671),
    .S1(net1017),
    .X(net186));
 sky130_fd_sc_hd__mux4_2 c325 (.A0(net179),
    .A1(net956),
    .A2(net947),
    .A3(net671),
    .S0(net1019),
    .S1(net1017),
    .X(net187));
 sky130_fd_sc_hd__mux4_1 c326 (.A0(net69),
    .A1(net186),
    .A2(net172),
    .A3(net829),
    .S0(net630),
    .S1(net650),
    .X(net188));
 sky130_fd_sc_hd__mux4_1 c327 (.A0(net187),
    .A1(net186),
    .A2(clknet_1_0__leaf_net169),
    .A3(net179),
    .S0(clknet_1_0__leaf_net613),
    .S1(clknet_1_0__leaf_net614),
    .X(net944));
 sky130_fd_sc_hd__a2111o_1 c328 (.A1(net179),
    .A2(clknet_1_0__leaf_net613),
    .B1(net947),
    .C1(net650),
    .D1(net1017),
    .X(net189));
 sky130_fd_sc_hd__mux4_1 c329 (.A0(net187),
    .A1(net186),
    .A2(clknet_1_0__leaf_net189),
    .A3(clknet_1_1__leaf_net613),
    .S0(clknet_1_0__leaf_net614),
    .S1(net1019),
    .X(net190));
 sky130_fd_sc_hd__mux4_1 c330 (.A0(clknet_1_1__leaf_net99),
    .A1(clknet_1_0__leaf_net169),
    .A2(net1054),
    .A3(net968),
    .S0(net661),
    .S1(net665),
    .X(net191));
 sky130_fd_sc_hd__mux4_2 c331 (.A0(net985),
    .A1(net972),
    .A2(net1034),
    .A3(net572),
    .S0(net658),
    .S1(net666),
    .X(net192));
 sky130_fd_sc_hd__mux4_1 c332 (.A0(net186),
    .A1(clknet_1_0__leaf_net96),
    .A2(net192),
    .A3(net827),
    .S0(net138),
    .S1(net84),
    .X(net193));
 sky130_fd_sc_hd__mux4_1 c333 (.A0(net968),
    .A1(clknet_1_1__leaf_net190),
    .A2(net65),
    .A3(net855),
    .S0(net842),
    .S1(net1064),
    .X(net194));
 sky130_fd_sc_hd__mux4_1 c334 (.A0(net842),
    .A1(net192),
    .A2(clknet_1_1__leaf_net944),
    .A3(net967),
    .S0(clknet_1_1__leaf_net924),
    .S1(net1022),
    .X(net195));
 sky130_fd_sc_hd__mux4_1 c335 (.A0(clknet_1_0__leaf_net190),
    .A1(net973),
    .A2(net572),
    .A3(net650),
    .S0(net669),
    .S1(net1020),
    .X(net196));
 sky130_fd_sc_hd__mux4_1 c336 (.A0(clknet_1_0__leaf_net99),
    .A1(clknet_1_1__leaf_net931),
    .A2(net848),
    .A3(net73),
    .S0(clknet_1_0__leaf_net196),
    .S1(net675),
    .X(net197));
 sky130_fd_sc_hd__mux4_2 c337 (.A0(clknet_1_0__leaf_net169),
    .A1(net972),
    .A2(net661),
    .A3(net671),
    .S0(net1017),
    .S1(net676),
    .X(net198));
 sky130_fd_sc_hd__mux4_1 c338 (.A0(net139),
    .A1(clknet_1_1__leaf_net99),
    .A2(net192),
    .A3(net130),
    .S0(clknet_1_0__leaf_net198),
    .S1(net572),
    .X(net199));
 sky130_fd_sc_hd__mux4_1 c339 (.A0(net973),
    .A1(clknet_1_1__leaf_net199),
    .A2(net1074),
    .A3(net992),
    .S0(net57),
    .S1(net650),
    .X(net200));
 sky130_fd_sc_hd__mux4_1 c340 (.A0(clknet_1_1__leaf_net196),
    .A1(clknet_1_1__leaf_net199),
    .A2(clknet_1_1__leaf_net99),
    .A3(net985),
    .S0(net665),
    .S1(net677),
    .X(net919));
 sky130_fd_sc_hd__mux4_1 c341 (.A0(clknet_1_1__leaf_net193),
    .A1(clknet_1_0__leaf_net199),
    .A2(clknet_1_1__leaf_net919),
    .A3(net1020),
    .S0(net671),
    .S1(net676),
    .X(net201));
 sky130_fd_sc_hd__mux4_1 c342 (.A0(net130),
    .A1(clknet_1_1__leaf_net200),
    .A2(clknet_1_1__leaf_net99),
    .A3(net186),
    .S0(net665),
    .S1(net677),
    .X(net202));
 sky130_fd_sc_hd__mux4_1 c343 (.A0(clknet_1_0__leaf_net199),
    .A1(clknet_1_0__leaf_net193),
    .A2(net84),
    .A3(clknet_1_0__leaf_net200),
    .S0(net669),
    .S1(net1017),
    .X(net203));
 sky130_fd_sc_hd__mux4_1 c344 (.A0(clknet_1_0__leaf_net200),
    .A1(net73),
    .A2(clknet_1_0__leaf_net199),
    .A3(clknet_1_1__leaf_net919),
    .S0(clknet_1_0__leaf_net196),
    .S1(net916),
    .X(net204));
 sky130_fd_sc_hd__mux4_1 c345 (.A0(net84),
    .A1(clknet_1_1__leaf_net200),
    .A2(net1064),
    .A3(net173),
    .S0(net678),
    .S1(net679),
    .X(net205));
 sky130_fd_sc_hd__mux4_1 c346 (.A0(clknet_1_0__leaf_net169),
    .A1(net864),
    .A2(clknet_1_1__leaf_net96),
    .A3(clknet_1_1__leaf_net919),
    .S0(net650),
    .S1(clknet_1_1__leaf_net680),
    .X(net206));
 sky130_fd_sc_hd__mux4_1 c347 (.A0(clknet_1_1__leaf_net919),
    .A1(clknet_1_1__leaf_net199),
    .A2(clknet_1_0__leaf_net96),
    .A3(net186),
    .S0(clknet_1_0__leaf_net933),
    .S1(net679),
    .X(net207));
 sky130_fd_sc_hd__mux4_1 c348 (.A0(net65),
    .A1(clknet_1_0__leaf_net199),
    .A2(net650),
    .A3(net658),
    .S0(net916),
    .S1(clknet_1_0__leaf_net680),
    .X(net938));
 sky130_fd_sc_hd__mux4_1 c349 (.A0(net934),
    .A1(clknet_1_0__leaf_net933),
    .A2(net669),
    .A3(net676),
    .S0(net678),
    .S1(net679),
    .X(net208));
 sky130_fd_sc_hd__mux4_1 c350 (.A0(clknet_1_1__leaf_net208),
    .A1(clknet_1_1__leaf_net938),
    .A2(net934),
    .A3(net650),
    .S0(clknet_1_1__leaf_net924),
    .S1(net678),
    .X(net209));
 sky130_fd_sc_hd__mux4_1 c351 (.A0(net864),
    .A1(clknet_1_0__leaf_net198),
    .A2(net978),
    .A3(net186),
    .S0(clknet_1_0__leaf_net614),
    .S1(clknet_1_1__leaf_net680),
    .X(net907));
 sky130_fd_sc_hd__mux4_1 c352 (.A0(net6),
    .A1(clknet_1_0__leaf_net927),
    .A2(clknet_1_0__leaf_net919),
    .A3(net115),
    .S0(net898),
    .S1(clknet_1_0__leaf_net680),
    .X(net210));
 sky130_fd_sc_hd__mux4_1 c353 (.A0(clknet_1_0__leaf_net105),
    .A1(net825),
    .A2(net7),
    .A3(clknet_1_0__leaf_net100),
    .S0(clknet_1_0__leaf_net931),
    .S1(net648),
    .X(net211));
 sky130_fd_sc_hd__mux4_1 c354 (.A0(clknet_1_0__leaf_net208),
    .A1(net940),
    .A2(net7),
    .A3(net179),
    .S0(net843),
    .S1(net648),
    .X(net212));
 sky130_fd_sc_hd__mux4_1 c355 (.A0(net810),
    .A1(clknet_1_1__leaf_net919),
    .A2(clknet_1_0__leaf_net897),
    .A3(net843),
    .S0(net956),
    .S1(clknet_1_0__leaf_net680),
    .X(net213));
 sky130_fd_sc_hd__mux4_1 c356 (.A0(net814),
    .A1(net872),
    .A2(net1032),
    .A3(net985),
    .S0(clknet_1_0__leaf_net902),
    .S1(clknet_1_0__leaf_net914),
    .X(net214));
 sky130_fd_sc_hd__mux4_1 c357 (.A0(net139),
    .A1(clknet_1_0__leaf_net944),
    .A2(net1035),
    .A3(clknet_1_1__leaf_net897),
    .S0(clknet_1_0__leaf_net214),
    .S1(net647),
    .X(net215));
 sky130_fd_sc_hd__mux4_1 c358 (.A0(clknet_1_0__leaf_net214),
    .A1(net1034),
    .A2(net1001),
    .A3(clknet_1_0__leaf_net111),
    .S0(net912),
    .S1(clknet_1_0__leaf_net914),
    .X(net216));
 sky130_fd_sc_hd__mux4_1 c359 (.A0(net943),
    .A1(clknet_1_0__leaf_net208),
    .A2(clknet_1_0__leaf_net105),
    .A3(net992),
    .S0(net934),
    .S1(clknet_1_0__leaf_net924),
    .X(net217));
 sky130_fd_sc_hd__mux4_1 c360 (.A0(net865),
    .A1(net139),
    .A2(net971),
    .A3(net843),
    .S0(clknet_1_0__leaf_net105),
    .S1(net630),
    .X(net218));
 sky130_fd_sc_hd__mux4_1 c361 (.A0(clknet_1_1__leaf_net111),
    .A1(clknet_1_0__leaf_net218),
    .A2(net992),
    .A3(clknet_1_1__leaf_net105),
    .S0(net641),
    .S1(clknet_1_1__leaf_net924),
    .X(net219));
 sky130_fd_sc_hd__mux4_1 c362 (.A0(net138),
    .A1(net971),
    .A2(clknet_1_0__leaf_net214),
    .A3(clknet_1_0__leaf_net933),
    .S0(net647),
    .S1(clknet_1_1__leaf_net924),
    .X(net220));
 sky130_fd_sc_hd__mux4_1 c363 (.A0(net215),
    .A1(clknet_1_1__leaf_net220),
    .A2(clknet_1_0__leaf_net214),
    .A3(net986),
    .S0(net936),
    .S1(clknet_1_0__leaf_net680),
    .X(net221));
 sky130_fd_sc_hd__mux4_1 c364 (.A0(clknet_1_0__leaf_net220),
    .A1(clknet_1_0__leaf_net214),
    .A2(clknet_1_0__leaf_net99),
    .A3(net1001),
    .S0(clknet_1_0__leaf_net218),
    .S1(net937),
    .X(net222));
 sky130_fd_sc_hd__mux4_1 c365 (.A0(clknet_1_0__leaf_net110),
    .A1(net6),
    .A2(clknet_1_0__leaf_net222),
    .A3(net7),
    .S0(clknet_1_0__leaf_net216),
    .S1(net648),
    .X(net223));
 sky130_fd_sc_hd__mux4_1 c366 (.A0(net221),
    .A1(net855),
    .A2(clknet_1_1__leaf_net220),
    .A3(net967),
    .S0(net1064),
    .S1(net116),
    .X(net224));
 sky130_fd_sc_hd__mux4_1 c367 (.A0(clknet_1_0__leaf_net928),
    .A1(clknet_1_0__leaf_net931),
    .A2(clknet_1_0__leaf_net222),
    .A3(net6),
    .S0(net648),
    .S1(net682),
    .X(net225));
 sky130_fd_sc_hd__mux4_1 c368 (.A0(clknet_1_1__leaf_net218),
    .A1(net985),
    .A2(clknet_1_1__leaf_net220),
    .A3(net950),
    .S0(net681),
    .S1(net683),
    .X(net226));
 sky130_fd_sc_hd__mux4_1 c369 (.A0(net102),
    .A1(clknet_1_0__leaf_net220),
    .A2(clknet_1_1__leaf_net218),
    .A3(net950),
    .S0(clknet_1_0__leaf_net914),
    .S1(net681),
    .X(net942));
 sky130_fd_sc_hd__mux4_1 c370 (.A0(net219),
    .A1(clknet_1_1__leaf_net222),
    .A2(clknet_1_1__leaf_net942),
    .A3(net872),
    .S0(net950),
    .S1(clknet_1_0__leaf_net902),
    .X(net227));
 sky130_fd_sc_hd__mux4_1 c371 (.A0(net217),
    .A1(clknet_1_1__leaf_net216),
    .A2(clknet_1_1__leaf_net942),
    .A3(net6),
    .S0(clknet_1_0__leaf_net931),
    .S1(net685),
    .X(net228));
 sky130_fd_sc_hd__mux4_1 c372 (.A0(net985),
    .A1(clknet_1_0__leaf_net226),
    .A2(clknet_1_1__leaf_net948),
    .A3(net7),
    .S0(net685),
    .S1(net687),
    .X(net229));
 sky130_fd_sc_hd__mux4_1 c373 (.A0(clknet_1_0__leaf_net222),
    .A1(clknet_1_1__leaf_net110),
    .A2(clknet_1_0__leaf_net942),
    .A3(net630),
    .S0(clknet_1_0__leaf_net914),
    .S1(net687),
    .X(net230));
 sky130_fd_sc_hd__a2111o_1 c396 (.A1(net127),
    .A2(net141),
    .B1(net148),
    .C1(net1076),
    .D1(net38),
    .X(net231));
 sky130_fd_sc_hd__a2111o_1 c397 (.A1(net982),
    .A2(net131),
    .B1(net845),
    .C1(net127),
    .D1(net145),
    .X(net232));
 sky130_fd_sc_hd__a2111o_1 c398 (.A1(net136),
    .A2(net975),
    .B1(net1054),
    .C1(net165),
    .D1(net1022),
    .X(net233));
 sky130_fd_sc_hd__sdfbbn_1 c399 (.CLK_N(clknet_4_7_0_clk),
    .D(net131),
    .RESET_B(net1033),
    .SCD(net964),
    .SCE(net975),
    .SET_B(net1048),
    .Q(net235),
    .Q_N(net234));
 sky130_fd_sc_hd__a2111o_1 c400 (.A1(net134),
    .A2(net235),
    .B1(net995),
    .C1(net975),
    .D1(net993),
    .X(net236));
 sky130_fd_sc_hd__mux4_1 c401 (.A0(net140),
    .A1(net235),
    .A2(net964),
    .A3(net132),
    .S0(net969),
    .S1(net608),
    .X(net237));
 sky130_fd_sc_hd__mux4_1 c402 (.A0(net235),
    .A1(net126),
    .A2(net972),
    .A3(net975),
    .S0(net964),
    .S1(net1015),
    .X(net238));
 sky130_fd_sc_hd__mux4_1 c403 (.A0(net975),
    .A1(net234),
    .A2(net969),
    .A3(net964),
    .S0(net608),
    .S1(net1015),
    .X(net239));
 sky130_fd_sc_hd__mux4_2 c404 (.A0(net38),
    .A1(net141),
    .A2(net29),
    .A3(net969),
    .S0(net608),
    .S1(net1015),
    .X(net240));
 sky130_fd_sc_hd__a2111o_1 c405 (.A1(net235),
    .A2(net969),
    .B1(net975),
    .C1(net638),
    .D1(net1015),
    .X(net241));
 sky130_fd_sc_hd__a2111o_1 c406 (.A1(net235),
    .A2(net146),
    .B1(net969),
    .C1(net975),
    .D1(net1015),
    .X(net242));
 sky130_fd_sc_hd__mux4_2 c407 (.A0(net135),
    .A1(net235),
    .A2(net845),
    .A3(net132),
    .S0(net969),
    .S1(net1015),
    .X(net243));
 sky130_fd_sc_hd__mux4_1 c408 (.A0(net35),
    .A1(net1028),
    .A2(net242),
    .A3(net234),
    .S0(net975),
    .S1(net608),
    .X(net244));
 sky130_fd_sc_hd__mux4_1 c409 (.A0(net244),
    .A1(net241),
    .A2(net964),
    .A3(net234),
    .S0(net969),
    .S1(net1015),
    .X(net245));
 sky130_fd_sc_hd__mux4_1 c410 (.A0(net964),
    .A1(net241),
    .A2(net234),
    .A3(net29),
    .S0(net976),
    .S1(net1015),
    .X(net246));
 sky130_fd_sc_hd__mux4_1 c411 (.A0(net242),
    .A1(net140),
    .A2(net244),
    .A3(net969),
    .S0(net640),
    .S1(net690),
    .X(net247));
 sky130_fd_sc_hd__mux4_2 c412 (.A0(net243),
    .A1(net234),
    .A2(net969),
    .A3(net975),
    .S0(net640),
    .S1(net1014),
    .X(net248));
 sky130_fd_sc_hd__mux4_1 c413 (.A0(net244),
    .A1(net148),
    .A2(net963),
    .A3(net638),
    .S0(net639),
    .S1(net1014),
    .X(net249));
 sky130_fd_sc_hd__mux4_1 c414 (.A0(net963),
    .A1(net242),
    .A2(net605),
    .A3(net1015),
    .S0(net690),
    .S1(net1014),
    .X(net250));
 sky130_fd_sc_hd__mux4_1 c415 (.A0(net963),
    .A1(net608),
    .A2(net638),
    .A3(net639),
    .S0(net1015),
    .S1(net1014),
    .X(net251));
 sky130_fd_sc_hd__mux4_1 c416 (.A0(net845),
    .A1(net963),
    .A2(net1047),
    .A3(net145),
    .S0(net915),
    .S1(net1014),
    .X(net252));
 sky130_fd_sc_hd__mux4_1 c417 (.A0(net126),
    .A1(net972),
    .A2(net146),
    .A3(net963),
    .S0(net969),
    .S1(net605),
    .X(net253));
 sky130_fd_sc_hd__mux4_2 c418 (.A0(net995),
    .A1(net154),
    .A2(net982),
    .A3(net802),
    .S0(net1027),
    .S1(net585),
    .X(net254));
 sky130_fd_sc_hd__mux4_1 c419 (.A0(net811),
    .A1(net964),
    .A2(net802),
    .A3(clknet_1_0__leaf_net169),
    .S0(net585),
    .S1(net692),
    .X(net255));
 sky130_fd_sc_hd__sdfbbn_1 c420 (.CLK_N(clknet_4_7_0_clk),
    .D(net254),
    .RESET_B(net966),
    .SCD(net1031),
    .SCE(net1023),
    .SET_B(net694),
    .Q(net257),
    .Q_N(net256));
 sky130_fd_sc_hd__mux4_1 c421 (.A0(net157),
    .A1(net154),
    .A2(net1035),
    .A3(net256),
    .S0(net915),
    .S1(net1016),
    .X(net258));
 sky130_fd_sc_hd__a2111o_1 c422 (.A1(net256),
    .A2(net1004),
    .B1(net1026),
    .C1(net566),
    .D1(net695),
    .X(net259));
 sky130_fd_sc_hd__mux4_1 c423 (.A0(net257),
    .A1(net972),
    .A2(net1053),
    .A3(net154),
    .S0(net1000),
    .S1(net695),
    .X(net260));
 sky130_fd_sc_hd__mux4_1 c424 (.A0(net257),
    .A1(net157),
    .A2(net961),
    .A3(net161),
    .S0(net695),
    .S1(net696),
    .X(net261));
 sky130_fd_sc_hd__mux4_1 c425 (.A0(clknet_1_0__leaf_net169),
    .A1(net962),
    .A2(net607),
    .A3(net915),
    .S0(net1016),
    .S1(net696),
    .X(net262));
 sky130_fd_sc_hd__mux4_1 c426 (.A0(net241),
    .A1(net1048),
    .A2(net961),
    .A3(net1000),
    .S0(net808),
    .S1(net1016),
    .X(net263));
 sky130_fd_sc_hd__mux4_1 c427 (.A0(net794),
    .A1(net993),
    .A2(net257),
    .A3(net1000),
    .S0(net962),
    .S1(net966),
    .X(net264));
 sky130_fd_sc_hd__mux4_1 c428 (.A0(net1050),
    .A1(net162),
    .A2(net1037),
    .A3(net962),
    .S0(net694),
    .S1(net697),
    .X(net265));
 sky130_fd_sc_hd__mux4_1 c429 (.A0(net962),
    .A1(net807),
    .A2(net1048),
    .A3(net637),
    .S0(net694),
    .S1(net697),
    .X(net266));
 sky130_fd_sc_hd__mux4_1 c430 (.A0(net794),
    .A1(net967),
    .A2(net1036),
    .A3(net608),
    .S0(net696),
    .S1(net1013),
    .X(net267));
 sky130_fd_sc_hd__mux4_1 c431 (.A0(net809),
    .A1(net1000),
    .A2(net962),
    .A3(net637),
    .S0(net1013),
    .S1(clknet_1_0__leaf_net699),
    .X(net268));
 sky130_fd_sc_hd__mux4_1 c432 (.A0(net56),
    .A1(clknet_1_1__leaf_net169),
    .A2(net147),
    .A3(net574),
    .S0(net1016),
    .S1(clknet_1_1__leaf_net699),
    .X(net269));
 sky130_fd_sc_hd__mux4_1 c433 (.A0(net154),
    .A1(net961),
    .A2(clknet_1_0__leaf_net269),
    .A3(net566),
    .S0(net1013),
    .S1(clknet_1_0__leaf_net699),
    .X(net270));
 sky130_fd_sc_hd__mux4_2 c434 (.A0(net979),
    .A1(clknet_1_0__leaf_net269),
    .A2(net56),
    .A3(net1000),
    .S0(clknet_1_1__leaf_net933),
    .S1(clknet_1_0__leaf_net700),
    .X(net271));
 sky130_fd_sc_hd__mux4_1 c435 (.A0(net967),
    .A1(clknet_1_0__leaf_net269),
    .A2(net1048),
    .A3(clknet_1_1__leaf_net271),
    .S0(clknet_1_0__leaf_net699),
    .S1(clknet_1_0__leaf_net700),
    .X(net272));
 sky130_fd_sc_hd__mux4_1 c436 (.A0(clknet_1_1__leaf_net271),
    .A1(net961),
    .A2(net802),
    .A3(net574),
    .S0(net1013),
    .S1(clknet_1_1__leaf_net699),
    .X(net273));
 sky130_fd_sc_hd__mux4_1 c437 (.A0(clknet_1_1__leaf_net269),
    .A1(clknet_1_1__leaf_net271),
    .A2(net961),
    .A3(clknet_1_1__leaf_net699),
    .S0(clknet_1_1__leaf_net700),
    .S1(net703),
    .X(net274));
 sky130_fd_sc_hd__mux4_1 c438 (.A0(clknet_1_1__leaf_net269),
    .A1(clknet_1_1__leaf_net271),
    .A2(net637),
    .A3(net915),
    .S0(net1013),
    .S1(clknet_1_1__leaf_net700),
    .X(net275));
 sky130_fd_sc_hd__mux4_1 c439 (.A0(clknet_1_0__leaf_net275),
    .A1(clknet_1_1__leaf_net271),
    .A2(clknet_1_1__leaf_net269),
    .A3(net566),
    .S0(clknet_1_1__leaf_net700),
    .S1(net702),
    .X(net276));
 sky130_fd_sc_hd__mux4_1 c440 (.A0(net187),
    .A1(clknet_1_1__leaf_net271),
    .A2(net161),
    .A3(net1004),
    .S0(net1018),
    .S1(net693),
    .X(net277));
 sky130_fd_sc_hd__a2111o_1 c441 (.A1(net813),
    .A2(net187),
    .B1(net162),
    .C1(net636),
    .D1(net693),
    .X(net278));
 sky130_fd_sc_hd__mux4_1 c442 (.A0(net162),
    .A1(net68),
    .A2(net977),
    .A3(net961),
    .S0(net615),
    .S1(net1020),
    .X(net279));
 sky130_fd_sc_hd__mux4_1 c443 (.A0(net977),
    .A1(clknet_1_1__leaf_net277),
    .A2(net187),
    .A3(clknet_1_0__leaf_net169),
    .S0(net643),
    .S1(clknet_1_1__leaf_net933),
    .X(net280));
 sky130_fd_sc_hd__mux4_1 c444 (.A0(net808),
    .A1(net961),
    .A2(net643),
    .A3(net650),
    .S0(net693),
    .S1(net705),
    .X(net281));
 sky130_fd_sc_hd__mux4_1 c445 (.A0(clknet_1_0__leaf_net189),
    .A1(net961),
    .A2(net978),
    .A3(clknet_1_1__leaf_net277),
    .S0(net973),
    .S1(net704),
    .X(net282));
 sky130_fd_sc_hd__mux4_1 c446 (.A0(clknet_1_0__leaf_net271),
    .A1(net187),
    .A2(net607),
    .A3(net658),
    .S0(net704),
    .S1(net707),
    .X(net283));
 sky130_fd_sc_hd__mux4_1 c447 (.A0(net52),
    .A1(net973),
    .A2(net607),
    .A3(net1018),
    .S0(net705),
    .S1(net706),
    .X(net284));
 sky130_fd_sc_hd__mux4_1 c448 (.A0(net1029),
    .A1(clknet_1_0__leaf_net271),
    .A2(net978),
    .A3(clknet_1_0__leaf_net283),
    .S0(net607),
    .S1(net708),
    .X(net285));
 sky130_fd_sc_hd__mux4_1 c449 (.A0(clknet_1_1__leaf_net189),
    .A1(net278),
    .A2(net967),
    .A3(net624),
    .S0(net636),
    .S1(net706),
    .X(net286));
 sky130_fd_sc_hd__mux4_2 c450 (.A0(net284),
    .A1(net162),
    .A2(net970),
    .A3(net615),
    .S0(net705),
    .S1(net707),
    .X(net287));
 sky130_fd_sc_hd__mux4_1 c451 (.A0(net278),
    .A1(net970),
    .A2(net1032),
    .A3(net624),
    .S0(clknet_1_1__leaf_net933),
    .S1(net707),
    .X(net288));
 sky130_fd_sc_hd__mux4_1 c452 (.A0(clknet_1_0__leaf_net288),
    .A1(net961),
    .A2(net650),
    .A3(net704),
    .S0(net706),
    .S1(net708),
    .X(net289));
 sky130_fd_sc_hd__mux4_1 c453 (.A0(net287),
    .A1(clknet_1_1__leaf_net288),
    .A2(net972),
    .A3(clknet_1_0__leaf_net271),
    .S0(net284),
    .S1(clknet_1_1__leaf_net933),
    .X(net917));
 sky130_fd_sc_hd__mux4_1 c454 (.A0(net287),
    .A1(clknet_1_1__leaf_net288),
    .A2(clknet_1_0__leaf_net917),
    .A3(net52),
    .S0(net915),
    .S1(net707),
    .X(net290));
 sky130_fd_sc_hd__mux4_1 c455 (.A0(clknet_1_1__leaf_net288),
    .A1(net609),
    .A2(net915),
    .A3(net643),
    .S0(net692),
    .S1(net708),
    .X(net291));
 sky130_fd_sc_hd__mux4_1 c456 (.A0(clknet_1_1__leaf_net291),
    .A1(net287),
    .A2(clknet_1_1__leaf_net189),
    .A3(net1051),
    .S0(net609),
    .S1(net708),
    .X(net292));
 sky130_fd_sc_hd__mux4_1 c457 (.A0(net972),
    .A1(net287),
    .A2(clknet_1_1__leaf_net291),
    .A3(net615),
    .S0(net658),
    .S1(net705),
    .X(net293));
 sky130_fd_sc_hd__mux4_1 c458 (.A0(clknet_1_1__leaf_net283),
    .A1(clknet_1_1__leaf_net291),
    .A2(net287),
    .A3(clknet_1_0__leaf_net917),
    .S0(net709),
    .S1(net1012),
    .X(net294));
 sky130_fd_sc_hd__mux4_1 c459 (.A0(clknet_1_0__leaf_net288),
    .A1(clknet_1_0__leaf_net291),
    .A2(net287),
    .A3(net961),
    .S0(net709),
    .S1(net1012),
    .X(net295));
 sky130_fd_sc_hd__mux4_1 c460 (.A0(clknet_1_0__leaf_net291),
    .A1(clknet_1_0__leaf_net288),
    .A2(net607),
    .A3(net643),
    .S0(net1020),
    .S1(net711),
    .X(net296));
 sky130_fd_sc_hd__mux4_1 c461 (.A0(net287),
    .A1(clknet_1_0__leaf_net288),
    .A2(clknet_1_0__leaf_net291),
    .A3(net947),
    .S0(net624),
    .S1(net711),
    .X(net297));
 sky130_fd_sc_hd__a2111o_2 c462 (.A1(net978),
    .A2(net974),
    .B1(net992),
    .C1(net597),
    .D1(net1012),
    .X(net298));
 sky130_fd_sc_hd__mux4_1 c463 (.A0(clknet_1_1__leaf_net96),
    .A1(clknet_1_0__leaf_net271),
    .A2(net973),
    .A3(net841),
    .S0(net1029),
    .S1(net692),
    .X(net299));
 sky130_fd_sc_hd__mux4_1 c464 (.A0(clknet_1_0__leaf_net907),
    .A1(net972),
    .A2(net978),
    .A3(net629),
    .S0(net1017),
    .S1(net692),
    .X(net911));
 sky130_fd_sc_hd__mux4_1 c465 (.A0(clknet_1_0__leaf_net277),
    .A1(net947),
    .A2(clknet_1_1__leaf_net924),
    .A3(net670),
    .S0(clknet_1_0__leaf_net701),
    .S1(net1012),
    .X(net300));
 sky130_fd_sc_hd__mux4_1 c466 (.A0(net848),
    .A1(net298),
    .A2(net1023),
    .A3(net670),
    .S0(net677),
    .S1(clknet_1_0__leaf_net701),
    .X(net301));
 sky130_fd_sc_hd__sdfbbp_1 c467 (.CLK(clknet_4_3_0_clk),
    .D(net808),
    .RESET_B(clknet_1_1__leaf_net911),
    .SCD(net965),
    .SCE(clknet_1_1__leaf_net614),
    .SET_B(net679),
    .Q(net303),
    .Q_N(net302));
 sky130_fd_sc_hd__mux4_1 c468 (.A0(clknet_1_0__leaf_net277),
    .A1(clknet_1_0__leaf_net301),
    .A2(net977),
    .A3(net1042),
    .S0(net829),
    .S1(net711),
    .X(net304));
 sky130_fd_sc_hd__mux4_1 c469 (.A0(clknet_1_0__leaf_net271),
    .A1(net1029),
    .A2(net302),
    .A3(clknet_1_0__leaf_net169),
    .S0(net636),
    .S1(net1012),
    .X(net305));
 sky130_fd_sc_hd__mux4_2 c470 (.A0(clknet_1_0__leaf_net198),
    .A1(net849),
    .A2(clknet_1_1__leaf_net96),
    .A3(net855),
    .S0(net298),
    .S1(net629),
    .X(net893));
 sky130_fd_sc_hd__mux4_1 c471 (.A0(clknet_1_1__leaf_net893),
    .A1(clknet_1_0__leaf_net299),
    .A2(clknet_1_1__leaf_net911),
    .A3(net641),
    .S0(net679),
    .S1(clknet_1_1__leaf_net680),
    .X(net306));
 sky130_fd_sc_hd__mux4_1 c472 (.A0(net841),
    .A1(net848),
    .A2(clknet_1_1__leaf_net893),
    .A3(clknet_1_0__leaf_net919),
    .S0(net1054),
    .S1(net896),
    .X(net307));
 sky130_fd_sc_hd__mux4_1 c473 (.A0(clknet_1_1__leaf_net911),
    .A1(clknet_1_1__leaf_net305),
    .A2(net303),
    .A3(clknet_1_1__leaf_net893),
    .S0(net1064),
    .S1(net597),
    .X(net308));
 sky130_fd_sc_hd__mux4_1 c474 (.A0(net972),
    .A1(clknet_1_0__leaf_net305),
    .A2(net978),
    .A3(net1026),
    .S0(net629),
    .S1(net896),
    .X(net309));
 sky130_fd_sc_hd__mux4_1 c475 (.A0(clknet_1_1__leaf_net305),
    .A1(net298),
    .A2(net302),
    .A3(net781),
    .S0(clknet_1_1__leaf_net614),
    .S1(net890),
    .X(net310));
 sky130_fd_sc_hd__mux4_2 c476 (.A0(net972),
    .A1(net192),
    .A2(net781),
    .A3(net607),
    .S0(net896),
    .S1(net658),
    .X(net311));
 sky130_fd_sc_hd__mux4_1 c477 (.A0(net311),
    .A1(net192),
    .A2(clknet_1_0__leaf_net305),
    .A3(clknet_1_1__leaf_net893),
    .S0(net890),
    .S1(net702),
    .X(net312));
 sky130_fd_sc_hd__mux4_1 c478 (.A0(clknet_1_0__leaf_net305),
    .A1(net1029),
    .A2(clknet_1_1__leaf_net198),
    .A3(clknet_1_0__leaf_net612),
    .S0(net896),
    .S1(net712),
    .X(net313));
 sky130_fd_sc_hd__mux4_1 c479 (.A0(clknet_1_1__leaf_net301),
    .A1(clknet_1_1__leaf_net305),
    .A2(clknet_1_1__leaf_net198),
    .A3(net192),
    .S0(net644),
    .S1(net693),
    .X(net314));
 sky130_fd_sc_hd__mux4_1 c480 (.A0(net311),
    .A1(clknet_1_1__leaf_net96),
    .A2(net678),
    .A3(net708),
    .S0(net1011),
    .S1(net712),
    .X(net315));
 sky130_fd_sc_hd__mux4_1 c481 (.A0(net311),
    .A1(clknet_1_1__leaf_net96),
    .A2(clknet_1_0__leaf_net315),
    .A3(net302),
    .S0(clknet_1_1__leaf_net680),
    .S1(net714),
    .X(net316));
 sky130_fd_sc_hd__mux4_1 c482 (.A0(clknet_1_1__leaf_net315),
    .A1(net311),
    .A2(clknet_1_0__leaf_net612),
    .A3(net891),
    .S0(net678),
    .S1(net713),
    .X(net317));
 sky130_fd_sc_hd__mux4_1 c483 (.A0(net311),
    .A1(net891),
    .A2(net920),
    .A3(clknet_1_0__leaf_net701),
    .S0(net1011),
    .S1(net712),
    .X(net925));
 sky130_fd_sc_hd__mux4_1 c484 (.A0(clknet_1_0__leaf_net911),
    .A1(net1005),
    .A2(net998),
    .A3(net641),
    .S0(net684),
    .S1(net1011),
    .X(net318));
 sky130_fd_sc_hd__mux4_1 c485 (.A0(net298),
    .A1(clknet_1_1__leaf_net911),
    .A2(clknet_1_1__leaf_net222),
    .A3(net865),
    .S0(net1023),
    .S1(net686),
    .X(net319));
 sky130_fd_sc_hd__mux4_1 c486 (.A0(clknet_1_0__leaf_net100),
    .A1(net912),
    .A2(net876),
    .A3(net629),
    .S0(clknet_1_1__leaf_net914),
    .S1(net685),
    .X(net320));
 sky130_fd_sc_hd__mux4_1 c487 (.A0(net192),
    .A1(net865),
    .A2(clknet_1_0__leaf_net911),
    .A3(net683),
    .S0(net687),
    .S1(net1011),
    .X(net321));
 sky130_fd_sc_hd__mux4_1 c488 (.A0(net971),
    .A1(clknet_1_1__leaf_net927),
    .A2(net1045),
    .A3(net684),
    .S0(net703),
    .S1(net715),
    .X(net322));
 sky130_fd_sc_hd__mux4_1 c489 (.A0(clknet_1_1__leaf_net214),
    .A1(net1005),
    .A2(net298),
    .A3(net644),
    .S0(clknet_1_0__leaf_net902),
    .S1(net687),
    .X(net918));
 sky130_fd_sc_hd__mux4_1 c490 (.A0(net303),
    .A1(net865),
    .A2(net642),
    .A3(net644),
    .S0(net681),
    .S1(net687),
    .X(net323));
 sky130_fd_sc_hd__mux4_1 c491 (.A0(clknet_1_1__leaf_net320),
    .A1(net4),
    .A2(net855),
    .A3(net916),
    .S0(net1011),
    .S1(net923),
    .X(net324));
 sky130_fd_sc_hd__a2111o_1 c492 (.A1(clknet_1_1__leaf_net105),
    .A2(net1005),
    .B1(net644),
    .C1(net920),
    .D1(net702),
    .X(net325));
 sky130_fd_sc_hd__mux4_1 c493 (.A0(clknet_1_0__leaf_net99),
    .A1(clknet_1_0__leaf_net925),
    .A2(net1001),
    .A3(clknet_1_0__leaf_net911),
    .S0(clknet_1_0__leaf_net320),
    .S1(net688),
    .X(net326));
 sky130_fd_sc_hd__mux4_1 c494 (.A0(net303),
    .A1(clknet_1_1__leaf_net928),
    .A2(net848),
    .A3(clknet_1_1__leaf_net325),
    .S0(clknet_1_1__leaf_net680),
    .S1(net716),
    .X(net327));
 sky130_fd_sc_hd__mux4_1 c495 (.A0(clknet_1_1__leaf_net105),
    .A1(net1022),
    .A2(clknet_1_1__leaf_net914),
    .A3(net682),
    .S0(net683),
    .S1(net687),
    .X(net328));
 sky130_fd_sc_hd__mux4_1 c496 (.A0(clknet_1_0__leaf_net325),
    .A1(clknet_1_1__leaf_net927),
    .A2(clknet_1_0__leaf_net328),
    .A3(clknet_1_1__leaf_net214),
    .S0(net682),
    .S1(net923),
    .X(net329));
 sky130_fd_sc_hd__mux4_1 c497 (.A0(net865),
    .A1(net912),
    .A2(clknet_1_1__leaf_net214),
    .A3(clknet_1_0__leaf_net99),
    .S0(net916),
    .S1(net715),
    .X(net330));
 sky130_fd_sc_hd__mux4_1 c498 (.A0(clknet_1_0__leaf_net330),
    .A1(net618),
    .A2(net629),
    .A3(net641),
    .S0(net920),
    .S1(net687),
    .X(net331));
 sky130_fd_sc_hd__mux4_1 c499 (.A0(clknet_1_1__leaf_net331),
    .A1(net298),
    .A2(clknet_1_1__leaf_net214),
    .A3(net618),
    .S0(net688),
    .S1(net716),
    .X(net332));
 sky130_fd_sc_hd__mux4_1 c500 (.A0(clknet_1_0__leaf_net330),
    .A1(clknet_1_0__leaf_net325),
    .A2(clknet_1_0__leaf_net919),
    .A3(net1023),
    .S0(net688),
    .S1(net716),
    .X(net333));
 sky130_fd_sc_hd__mux4_1 c501 (.A0(net323),
    .A1(clknet_1_1__leaf_net325),
    .A2(clknet_1_1__leaf_net214),
    .A3(clknet_1_1__leaf_net918),
    .S0(net920),
    .S1(net716),
    .X(net922));
 sky130_fd_sc_hd__mux4_1 c502 (.A0(net1044),
    .A1(clknet_1_1__leaf_net222),
    .A2(clknet_1_0__leaf_net928),
    .A3(net629),
    .S0(net916),
    .S1(net687),
    .X(net334));
 sky130_fd_sc_hd__mux4_1 c503 (.A0(clknet_1_0__leaf_net331),
    .A1(net641),
    .A2(net920),
    .A3(net916),
    .S0(net687),
    .S1(net717),
    .X(net335));
 sky130_fd_sc_hd__mux4_1 c504 (.A0(net4),
    .A1(net865),
    .A2(net915),
    .A3(net1011),
    .S0(net716),
    .S1(net718),
    .X(net930));
 sky130_fd_sc_hd__mux4_1 c505 (.A0(clknet_1_1__leaf_net922),
    .A1(clknet_1_1__leaf_net330),
    .A2(clknet_1_1__leaf_net914),
    .A3(net684),
    .S0(net717),
    .S1(net718),
    .X(net336));
 sky130_fd_sc_hd__sdfbbn_1 c528 (.CLK_N(clknet_4_13_0_clk),
    .D(net975),
    .RESET_B(net1036),
    .SCD(net141),
    .SCE(net963),
    .SET_B(net690),
    .Q(net338),
    .Q_N(net337));
 sky130_fd_sc_hd__sdfbbn_1 c529 (.CLK_N(clknet_4_13_0_clk),
    .D(net141),
    .RESET_B(net1072),
    .SCD(net148),
    .SCE(net165),
    .SET_B(net1071),
    .Q(net340),
    .Q_N(net339));
 sky130_fd_sc_hd__sdfbbp_1 c530 (.CLK(clknet_4_13_0_clk),
    .D(net36),
    .RESET_B(net780),
    .SCD(net339),
    .SCE(net963),
    .SET_B(net1014),
    .Q(net342),
    .Q_N(net341));
 sky130_fd_sc_hd__mux4_1 c531 (.A0(net788),
    .A1(net342),
    .A2(net141),
    .A3(net339),
    .S0(net337),
    .S1(net609),
    .X(net343));
 sky130_fd_sc_hd__mux4_2 c532 (.A0(net342),
    .A1(net338),
    .A2(net788),
    .A3(net339),
    .S0(net655),
    .S1(net1022),
    .X(net344));
 sky130_fd_sc_hd__mux4_2 c533 (.A0(net340),
    .A1(net338),
    .A2(net341),
    .A3(net609),
    .S0(net655),
    .S1(net692),
    .X(net345));
 sky130_fd_sc_hd__mux4_1 c534 (.A0(net29),
    .A1(net344),
    .A2(net248),
    .A3(net341),
    .S0(net145),
    .S1(net690),
    .X(net346));
 sky130_fd_sc_hd__mux4_1 c535 (.A0(net344),
    .A1(net248),
    .A2(net337),
    .A3(net1006),
    .S0(net640),
    .S1(net692),
    .X(net347));
 sky130_fd_sc_hd__mux4_1 c536 (.A0(net342),
    .A1(net963),
    .A2(net1006),
    .A3(net339),
    .S0(net563),
    .S1(clknet_1_1__leaf_net720),
    .X(net348));
 sky130_fd_sc_hd__mux4_1 c537 (.A0(net963),
    .A1(net243),
    .A2(net1006),
    .A3(net563),
    .S0(clknet_1_1__leaf_net720),
    .S1(clknet_1_1__leaf_net721),
    .X(net349));
 sky130_fd_sc_hd__mux4_1 c538 (.A0(net344),
    .A1(net36),
    .A2(net963),
    .A3(clknet_1_1__leaf_net720),
    .S0(clknet_1_0__leaf_net721),
    .S1(net723),
    .X(net350));
 sky130_fd_sc_hd__mux4_1 c539 (.A0(net243),
    .A1(net341),
    .A2(net1006),
    .A3(net691),
    .S0(clknet_1_1__leaf_net720),
    .S1(net722),
    .X(net351));
 sky130_fd_sc_hd__mux4_1 c540 (.A0(net341),
    .A1(net248),
    .A2(net609),
    .A3(clknet_1_1__leaf_net720),
    .S0(clknet_1_1__leaf_net721),
    .S1(net723),
    .X(net352));
 sky130_fd_sc_hd__mux4_1 c541 (.A0(net344),
    .A1(clknet_1_1__leaf_net351),
    .A2(net337),
    .A3(net562),
    .S0(clknet_1_1__leaf_net721),
    .S1(net724),
    .X(net353));
 sky130_fd_sc_hd__mux4_1 c542 (.A0(net1028),
    .A1(net655),
    .A2(net1016),
    .A3(clknet_1_0__leaf_net720),
    .S0(net725),
    .S1(net726),
    .X(net354));
 sky130_fd_sc_hd__mux4_1 c543 (.A0(net1006),
    .A1(clknet_1_1__leaf_net354),
    .A2(net655),
    .A3(clknet_1_0__leaf_net720),
    .S0(clknet_1_0__leaf_net721),
    .S1(net724),
    .X(net355));
 sky130_fd_sc_hd__mux4_1 c544 (.A0(clknet_1_1__leaf_net354),
    .A1(clknet_1_0__leaf_net351),
    .A2(clknet_1_0__leaf_net355),
    .A3(clknet_1_0__leaf_net720),
    .S0(net724),
    .S1(net726),
    .X(net356));
 sky130_fd_sc_hd__mux4_1 c545 (.A0(clknet_1_0__leaf_net351),
    .A1(clknet_1_1__leaf_net354),
    .A2(net145),
    .A3(net341),
    .S0(clknet_1_1__leaf_net645),
    .S1(net1016),
    .X(net357));
 sky130_fd_sc_hd__mux4_1 c546 (.A0(net342),
    .A1(clknet_1_1__leaf_net354),
    .A2(net345),
    .A3(net562),
    .S0(clknet_1_1__leaf_net645),
    .S1(net727),
    .X(net358));
 sky130_fd_sc_hd__mux4_1 c547 (.A0(clknet_1_1__leaf_net351),
    .A1(clknet_1_0__leaf_net358),
    .A2(clknet_1_1__leaf_net354),
    .A3(clknet_1_0__leaf_net720),
    .S0(net725),
    .S1(net728),
    .X(net359));
 sky130_fd_sc_hd__mux4_1 c548 (.A0(clknet_1_1__leaf_net355),
    .A1(clknet_1_0__leaf_net358),
    .A2(net342),
    .A3(net562),
    .S0(clknet_1_1__leaf_net645),
    .S1(net690),
    .X(net360));
 sky130_fd_sc_hd__mux4_1 c549 (.A0(clknet_1_0__leaf_net355),
    .A1(net360),
    .A2(clknet_1_0__leaf_net720),
    .A3(net722),
    .S0(net728),
    .S1(net904),
    .X(net361));
 sky130_fd_sc_hd__mux4_1 c550 (.A0(net340),
    .A1(net996),
    .A2(net998),
    .A3(net976),
    .S0(net574),
    .S1(net1023),
    .X(net362));
 sky130_fd_sc_hd__mux4_1 c551 (.A0(net56),
    .A1(net1000),
    .A2(net362),
    .A3(net966),
    .S0(clknet_1_1__leaf_net275),
    .S1(net728),
    .X(net363));
 sky130_fd_sc_hd__a2111o_1 c552 (.A1(net1040),
    .A2(net966),
    .B1(net808),
    .C1(net574),
    .D1(net1022),
    .X(net364));
 sky130_fd_sc_hd__a2111o_1 c553 (.A1(net816),
    .A2(net976),
    .B1(net340),
    .C1(clknet_1_1__leaf_net361),
    .D1(net1000),
    .X(net365));
 sky130_fd_sc_hd__a2111o_1 c554 (.A1(net1026),
    .A2(net604),
    .B1(clknet_1_1__leaf_net645),
    .C1(net1023),
    .D1(net697),
    .X(net366));
 sky130_fd_sc_hd__mux4_1 c555 (.A0(net813),
    .A1(net979),
    .A2(net52),
    .A3(net604),
    .S0(net1013),
    .S1(net729),
    .X(net367));
 sky130_fd_sc_hd__mux4_1 c556 (.A0(net367),
    .A1(clknet_1_1__leaf_net366),
    .A2(net340),
    .A3(net980),
    .S0(net728),
    .S1(net904),
    .X(net368));
 sky130_fd_sc_hd__a2111o_1 c557 (.A1(net362),
    .A2(clknet_1_1__leaf_net368),
    .B1(net1022),
    .C1(net904),
    .D1(net729),
    .X(net369));
 sky130_fd_sc_hd__mux4_1 c558 (.A0(net367),
    .A1(clknet_1_0__leaf_net369),
    .A2(net976),
    .A3(clknet_1_1__leaf_net169),
    .S0(clknet_1_1__leaf_net368),
    .S1(net697),
    .X(net370));
 sky130_fd_sc_hd__a2111o_1 c559 (.A1(net362),
    .A2(net52),
    .B1(clknet_1_1__leaf_net369),
    .C1(clknet_1_1__leaf_net365),
    .D1(clknet_1_0__leaf_net645),
    .X(net371));
 sky130_fd_sc_hd__sdfbbn_1 c560 (.CLK_N(clknet_4_14_0_clk),
    .D(clknet_1_1__leaf_net369),
    .RESET_B(net998),
    .SCD(net996),
    .SCE(net563),
    .SET_B(net1013),
    .Q(net373),
    .Q_N(net372));
 sky130_fd_sc_hd__mux4_1 c561 (.A0(net57),
    .A1(net980),
    .A2(clknet_1_1__leaf_net366),
    .A3(net372),
    .S0(net654),
    .S1(net1013),
    .X(net909));
 sky130_fd_sc_hd__mux4_1 c562 (.A0(net56),
    .A1(clknet_1_0__leaf_net369),
    .A2(net372),
    .A3(clknet_1_0__leaf_net909),
    .S0(net654),
    .S1(net729),
    .X(net374));
 sky130_fd_sc_hd__mux4_1 c563 (.A0(net802),
    .A1(net1040),
    .A2(net980),
    .A3(clknet_1_0__leaf_net645),
    .S0(net1013),
    .S1(net730),
    .X(net375));
 sky130_fd_sc_hd__mux4_1 c564 (.A0(clknet_1_0__leaf_net375),
    .A1(clknet_1_0__leaf_net368),
    .A2(clknet_1_0__leaf_net909),
    .A3(clknet_1_1__leaf_net366),
    .S0(clknet_1_0__leaf_net645),
    .S1(net730),
    .X(net376));
 sky130_fd_sc_hd__mux4_1 c565 (.A0(net372),
    .A1(net254),
    .A2(clknet_1_0__leaf_net369),
    .A3(clknet_1_0__leaf_net376),
    .S0(net605),
    .S1(net730),
    .X(net377));
 sky130_fd_sc_hd__mux4_1 c566 (.A0(net980),
    .A1(clknet_1_0__leaf_net375),
    .A2(clknet_1_1__leaf_net361),
    .A3(clknet_1_1__leaf_net369),
    .S0(net635),
    .S1(net730),
    .X(net378));
 sky130_fd_sc_hd__mux4_1 c567 (.A0(clknet_1_0__leaf_net368),
    .A1(clknet_1_0__leaf_net909),
    .A2(net991),
    .A3(net980),
    .S0(net635),
    .S1(net1010),
    .X(net379));
 sky130_fd_sc_hd__mux4_1 c568 (.A0(clknet_1_0__leaf_net379),
    .A1(net1000),
    .A2(clknet_1_1__leaf_net376),
    .A3(net635),
    .S0(net730),
    .S1(net1010),
    .X(net380));
 sky130_fd_sc_hd__mux4_1 c569 (.A0(clknet_1_1__leaf_net379),
    .A1(net373),
    .A2(clknet_1_1__leaf_net376),
    .A3(net730),
    .S0(net1010),
    .S1(net733),
    .X(net381));
 sky130_fd_sc_hd__mux4_1 c570 (.A0(clknet_1_0__leaf_net376),
    .A1(net373),
    .A2(net259),
    .A3(clknet_1_0__leaf_net366),
    .S0(net696),
    .S1(net733),
    .X(net382));
 sky130_fd_sc_hd__mux4_1 c571 (.A0(clknet_1_1__leaf_net369),
    .A1(net1050),
    .A2(net373),
    .A3(clknet_1_1__leaf_net365),
    .S0(net654),
    .S1(net734),
    .X(net383));
 sky130_fd_sc_hd__mux4_1 c572 (.A0(net182),
    .A1(net825),
    .A2(net1029),
    .A3(net906),
    .S0(net729),
    .S1(net734),
    .X(net384));
 sky130_fd_sc_hd__mux4_1 c573 (.A0(net978),
    .A1(net384),
    .A2(net1029),
    .A3(net808),
    .S0(clknet_1_0__leaf_net701),
    .S1(net709),
    .X(net385));
 sky130_fd_sc_hd__mux4_1 c574 (.A0(net384),
    .A1(net813),
    .A2(clknet_1_0__leaf_net354),
    .A3(net658),
    .S0(net693),
    .S1(net702),
    .X(net386));
 sky130_fd_sc_hd__mux4_1 c575 (.A0(clknet_1_0__leaf_net375),
    .A1(net182),
    .A2(clknet_1_1__leaf_net169),
    .A3(clknet_1_1__leaf_net701),
    .S0(net709),
    .S1(net1012),
    .X(net387));
 sky130_fd_sc_hd__mux4_1 c576 (.A0(clknet_1_0__leaf_net366),
    .A1(net182),
    .A2(clknet_1_1__leaf_net385),
    .A3(net702),
    .S0(net710),
    .S1(net729),
    .X(net388));
 sky130_fd_sc_hd__mux4_1 c577 (.A0(clknet_1_0__leaf_net385),
    .A1(clknet_1_0__leaf_net386),
    .A2(clknet_1_0__leaf_net387),
    .A3(net692),
    .S0(net709),
    .S1(net732),
    .X(net389));
 sky130_fd_sc_hd__mux4_1 c578 (.A0(clknet_1_0__leaf_net389),
    .A1(net170),
    .A2(net1006),
    .A3(clknet_1_0__leaf_net387),
    .S0(net1026),
    .S1(net702),
    .X(net390));
 sky130_fd_sc_hd__mux4_1 c579 (.A0(net1033),
    .A1(net170),
    .A2(net977),
    .A3(clknet_1_0__leaf_net645),
    .S0(net1012),
    .S1(net888),
    .X(net391));
 sky130_fd_sc_hd__mux4_1 c580 (.A0(clknet_1_0__leaf_net354),
    .A1(net182),
    .A2(net654),
    .A3(clknet_1_1__leaf_net701),
    .S0(net1010),
    .S1(net888),
    .X(net392));
 sky130_fd_sc_hd__mux4_1 c581 (.A0(clknet_1_0__leaf_net387),
    .A1(clknet_1_0__leaf_net917),
    .A2(net182),
    .A3(clknet_1_0__leaf_net388),
    .S0(net1018),
    .S1(net888),
    .X(net393));
 sky130_fd_sc_hd__mux4_1 c582 (.A0(clknet_1_1__leaf_net361),
    .A1(net182),
    .A2(net998),
    .A3(clknet_1_0__leaf_net387),
    .S0(net729),
    .S1(net737),
    .X(net394));
 sky130_fd_sc_hd__mux4_1 c583 (.A0(clknet_1_0__leaf_net394),
    .A1(clknet_1_0__leaf_net388),
    .A2(net52),
    .A3(clknet_1_0__leaf_net387),
    .S0(clknet_1_1__leaf_net389),
    .S1(net737),
    .X(net395));
 sky130_fd_sc_hd__mux4_1 c584 (.A0(clknet_1_0__leaf_net366),
    .A1(clknet_1_1__leaf_net392),
    .A2(clknet_1_0__leaf_net394),
    .A3(net560),
    .S0(net906),
    .S1(net888),
    .X(net396));
 sky130_fd_sc_hd__mux4_1 c585 (.A0(clknet_1_1__leaf_net386),
    .A1(clknet_1_0__leaf_net361),
    .A2(clknet_1_1__leaf_net394),
    .A3(net52),
    .S0(net1012),
    .S1(clknet_1_1__leaf_net738),
    .X(net397));
 sky130_fd_sc_hd__mux4_1 c586 (.A0(clknet_1_0__leaf_net354),
    .A1(clknet_1_1__leaf_net387),
    .A2(clknet_1_1__leaf_net394),
    .A3(net736),
    .S0(net737),
    .S1(clknet_1_1__leaf_net739),
    .X(net398));
 sky130_fd_sc_hd__mux4_1 c587 (.A0(clknet_1_0__leaf_net392),
    .A1(net994),
    .A2(net1006),
    .A3(net732),
    .S0(clknet_1_0__leaf_net739),
    .S1(clknet_1_0__leaf_net740),
    .X(net399));
 sky130_fd_sc_hd__mux4_1 c588 (.A0(clknet_1_1__leaf_net388),
    .A1(clknet_1_0__leaf_net392),
    .A2(clknet_1_1__leaf_net399),
    .A3(net709),
    .S0(clknet_1_1__leaf_net738),
    .S1(clknet_1_0__leaf_net739),
    .X(net400));
 sky130_fd_sc_hd__mux4_1 c589 (.A0(net373),
    .A1(clknet_1_1__leaf_net387),
    .A2(clknet_1_1__leaf_net399),
    .A3(clknet_1_1__leaf_net400),
    .S0(clknet_1_0__leaf_net739),
    .S1(clknet_1_0__leaf_net740),
    .X(net401));
 sky130_fd_sc_hd__mux4_1 c590 (.A0(clknet_1_1__leaf_net391),
    .A1(clknet_1_0__leaf_net354),
    .A2(net560),
    .A3(net709),
    .S0(net1010),
    .S1(clknet_1_1__leaf_net739),
    .X(net402));
 sky130_fd_sc_hd__mux4_1 c591 (.A0(clknet_1_0__leaf_net400),
    .A1(clknet_1_1__leaf_net402),
    .A2(net559),
    .A3(net693),
    .S0(net737),
    .S1(clknet_1_0__leaf_net738),
    .X(net403));
 sky130_fd_sc_hd__mux4_1 c592 (.A0(clknet_1_1__leaf_net392),
    .A1(net559),
    .A2(net709),
    .A3(clknet_1_0__leaf_net738),
    .S0(clknet_1_0__leaf_net739),
    .S1(net741),
    .X(net404));
 sky130_fd_sc_hd__mux4_1 c593 (.A0(clknet_1_0__leaf_net391),
    .A1(clknet_1_1__leaf_net402),
    .A2(net991),
    .A3(net709),
    .S0(net1012),
    .S1(clknet_1_1__leaf_net739),
    .X(net405));
 sky130_fd_sc_hd__mux4_1 c594 (.A0(net848),
    .A1(clknet_1_0__leaf_net299),
    .A2(clknet_1_1__leaf_net100),
    .A3(net674),
    .S0(clknet_1_0__leaf_net701),
    .S1(net710),
    .X(net406));
 sky130_fd_sc_hd__mux4_1 c595 (.A0(net1030),
    .A1(clknet_1_1__leaf_net893),
    .A2(net659),
    .A3(net693),
    .S0(net712),
    .S1(net714),
    .X(net407));
 sky130_fd_sc_hd__mux4_1 c596 (.A0(clknet_1_1__leaf_net404),
    .A1(net560),
    .A2(net702),
    .A3(net710),
    .S0(net904),
    .S1(net733),
    .X(net908));
 sky130_fd_sc_hd__mux4_1 c597 (.A0(clknet_1_1__leaf_net405),
    .A1(clknet_1_0__leaf_net893),
    .A2(clknet_1_0__leaf_net908),
    .A3(clknet_1_1__leaf_net399),
    .S0(net659),
    .S1(net678),
    .X(net408));
 sky130_fd_sc_hd__mux4_1 c598 (.A0(clknet_1_1__leaf_net299),
    .A1(clknet_1_1__leaf_net893),
    .A2(clknet_1_0__leaf_net908),
    .A3(net1012),
    .S0(net732),
    .S1(net735),
    .X(net409));
 sky130_fd_sc_hd__mux4_1 c599 (.A0(clknet_1_1__leaf_net299),
    .A1(net965),
    .A2(net170),
    .A3(net659),
    .S0(net904),
    .S1(net741),
    .X(net410));
 sky130_fd_sc_hd__mux4_1 c600 (.A0(net808),
    .A1(clknet_1_0__leaf_net365),
    .A2(clknet_1_0__leaf_net299),
    .A3(net978),
    .S0(net68),
    .S1(net659),
    .X(net411));
 sky130_fd_sc_hd__mux4_1 c601 (.A0(net1055),
    .A1(clknet_1_0__leaf_net893),
    .A2(net1041),
    .A3(net735),
    .S0(net741),
    .S1(net745),
    .X(net412));
 sky130_fd_sc_hd__mux4_1 c602 (.A0(clknet_1_0__leaf_net361),
    .A1(net170),
    .A2(clknet_1_0__leaf_net907),
    .A3(net920),
    .S0(net659),
    .S1(net734),
    .X(net413));
 sky130_fd_sc_hd__mux4_1 c603 (.A0(clknet_1_1__leaf_net169),
    .A1(net1053),
    .A2(clknet_1_0__leaf_net405),
    .A3(clknet_1_0__leaf_net361),
    .S0(clknet_1_0__leaf_net412),
    .S1(clknet_1_1__leaf_net299),
    .X(net414));
 sky130_fd_sc_hd__mux4_1 c604 (.A0(net413),
    .A1(clknet_1_0__leaf_net361),
    .A2(net855),
    .A3(net967),
    .S0(net674),
    .S1(net735),
    .X(net415));
 sky130_fd_sc_hd__mux4_1 c605 (.A0(clknet_1_1__leaf_net299),
    .A1(net631),
    .A2(net693),
    .A3(net703),
    .S0(net733),
    .S1(net743),
    .X(net416));
 sky130_fd_sc_hd__mux4_2 c606 (.A0(net974),
    .A1(net678),
    .A2(net904),
    .A3(net732),
    .S0(net745),
    .S1(net747),
    .X(net417));
 sky130_fd_sc_hd__mux4_1 c607 (.A0(net977),
    .A1(clknet_1_0__leaf_net365),
    .A2(net417),
    .A3(clknet_1_0__leaf_net908),
    .S0(net631),
    .S1(net744),
    .X(net892));
 sky130_fd_sc_hd__mux4_1 c608 (.A0(net407),
    .A1(clknet_1_1__leaf_net892),
    .A2(net417),
    .A3(net744),
    .S0(net746),
    .S1(net747),
    .X(net418));
 sky130_fd_sc_hd__mux4_1 c609 (.A0(net977),
    .A1(clknet_1_1__leaf_net892),
    .A2(net631),
    .A3(net1018),
    .S0(net742),
    .S1(net747),
    .X(net419));
 sky130_fd_sc_hd__mux4_1 c610 (.A0(net417),
    .A1(clknet_1_1__leaf_net399),
    .A2(net653),
    .A3(net712),
    .S0(net903),
    .S1(net747),
    .X(net420));
 sky130_fd_sc_hd__mux4_1 c611 (.A0(net417),
    .A1(clknet_1_0__leaf_net420),
    .A2(clknet_1_0__leaf_net405),
    .A3(net974),
    .S0(net653),
    .S1(net746),
    .X(net421));
 sky130_fd_sc_hd__mux4_1 c612 (.A0(clknet_1_0__leaf_net421),
    .A1(clknet_1_1__leaf_net420),
    .A2(clknet_1_0__leaf_net365),
    .A3(net745),
    .S0(net746),
    .S1(net748),
    .X(net422));
 sky130_fd_sc_hd__mux4_1 c613 (.A0(clknet_1_0__leaf_net420),
    .A1(net965),
    .A2(net1036),
    .A3(clknet_1_1__leaf_net169),
    .S0(clknet_1_0__leaf_net421),
    .S1(net653),
    .X(net423));
 sky130_fd_sc_hd__mux4_1 c614 (.A0(clknet_1_1__leaf_net420),
    .A1(net894),
    .A2(net904),
    .A3(net903),
    .S0(net746),
    .S1(net748),
    .X(net424));
 sky130_fd_sc_hd__mux4_1 c615 (.A0(net424),
    .A1(clknet_1_0__leaf_net908),
    .A2(clknet_1_1__leaf_net421),
    .A3(net625),
    .S0(net653),
    .S1(net675),
    .X(net425));
 sky130_fd_sc_hd__mux4_1 c616 (.A0(net116),
    .A1(clknet_1_0__leaf_net100),
    .A2(net1001),
    .A3(clknet_1_0__leaf_net402),
    .S0(net686),
    .S1(net742),
    .X(net426));
 sky130_fd_sc_hd__mux4_1 c617 (.A0(clknet_1_0__leaf_net402),
    .A1(net971),
    .A2(clknet_1_0__leaf_net331),
    .A3(net1005),
    .S0(clknet_1_0__leaf_net100),
    .S1(net1030),
    .X(net427));
 sky130_fd_sc_hd__mux4_1 c618 (.A0(clknet_1_0__leaf_net328),
    .A1(net1001),
    .A2(clknet_1_0__leaf_net365),
    .A3(clknet_1_0__leaf_net399),
    .S0(clknet_1_1__leaf_net902),
    .S1(net686),
    .X(net428));
 sky130_fd_sc_hd__mux4_1 c619 (.A0(clknet_1_0__leaf_net100),
    .A1(net856),
    .A2(clknet_1_0__leaf_net917),
    .A3(net967),
    .S0(clknet_1_0__leaf_net328),
    .S1(net688),
    .X(net429));
 sky130_fd_sc_hd__mux4_1 c620 (.A0(net855),
    .A1(clknet_1_1__leaf_net328),
    .A2(net876),
    .A3(net896),
    .S0(net743),
    .S1(net886),
    .X(net430));
 sky130_fd_sc_hd__mux4_1 c621 (.A0(net895),
    .A1(net855),
    .A2(clknet_1_0__leaf_net907),
    .A3(net641),
    .S0(clknet_1_0__leaf_net701),
    .S1(clknet_1_0__leaf_net719),
    .X(net431));
 sky130_fd_sc_hd__mux4_1 c622 (.A0(net1024),
    .A1(clknet_1_1__leaf_net897),
    .A2(net641),
    .A3(net642),
    .S0(net891),
    .S1(net742),
    .X(net432));
 sky130_fd_sc_hd__mux4_1 c623 (.A0(clknet_1_0__leaf_net399),
    .A1(net432),
    .A2(net1030),
    .A3(clknet_1_0__leaf_net893),
    .S0(net900),
    .S1(net886),
    .X(net899));
 sky130_fd_sc_hd__mux4_1 c624 (.A0(net426),
    .A1(net876),
    .A2(net971),
    .A3(clknet_1_1__leaf_net331),
    .S0(clknet_1_1__leaf_net902),
    .S1(net681),
    .X(net433));
 sky130_fd_sc_hd__mux4_1 c625 (.A0(clknet_1_1__leaf_net331),
    .A1(clknet_1_0__leaf_net226),
    .A2(clknet_1_0__leaf_net100),
    .A3(net116),
    .S0(net642),
    .S1(net718),
    .X(net434));
 sky130_fd_sc_hd__mux4_1 c626 (.A0(net431),
    .A1(clknet_1_1__leaf_net907),
    .A2(clknet_1_1__leaf_net328),
    .A3(net682),
    .S0(net749),
    .S1(net752),
    .X(net435));
 sky130_fd_sc_hd__mux4_1 c627 (.A0(clknet_1_0__leaf_net365),
    .A1(clknet_1_0__leaf_net399),
    .A2(clknet_1_1__leaf_net909),
    .A3(clknet_1_1__leaf_net899),
    .S0(net994),
    .S1(net903),
    .X(net436));
 sky130_fd_sc_hd__mux4_1 c628 (.A0(net116),
    .A1(clknet_1_0__leaf_net909),
    .A2(clknet_1_1__leaf_net899),
    .A3(net668),
    .S0(net886),
    .S1(net752),
    .X(net437));
 sky130_fd_sc_hd__a2111o_1 c629 (.A1(net1005),
    .A2(clknet_1_1__leaf_net899),
    .B1(clknet_1_0__leaf_net893),
    .C1(net642),
    .D1(net682),
    .X(net438));
 sky130_fd_sc_hd__mux4_1 c630 (.A0(net430),
    .A1(clknet_1_0__leaf_net899),
    .A2(net596),
    .A3(net885),
    .S0(net718),
    .S1(net751),
    .X(net439));
 sky130_fd_sc_hd__mux4_1 c631 (.A0(net1006),
    .A1(clknet_1_1__leaf_net897),
    .A2(clknet_1_1__leaf_net907),
    .A3(clknet_1_1__leaf_net428),
    .S0(clknet_1_1__leaf_net100),
    .S1(net596),
    .X(net440));
 sky130_fd_sc_hd__mux4_1 c632 (.A0(net116),
    .A1(clknet_1_1__leaf_net897),
    .A2(net718),
    .A3(net743),
    .S0(net886),
    .S1(net752),
    .X(net441));
 sky130_fd_sc_hd__mux4_1 c633 (.A0(clknet_1_0__leaf_net892),
    .A1(net1056),
    .A2(net1031),
    .A3(net890),
    .S0(net642),
    .S1(net750),
    .X(net442));
 sky130_fd_sc_hd__mux4_1 c634 (.A0(clknet_1_1__leaf_net328),
    .A1(net441),
    .A2(clknet_1_0__leaf_net899),
    .A3(net688),
    .S0(net718),
    .S1(net751),
    .X(net443));
 sky130_fd_sc_hd__mux4_1 c635 (.A0(net1050),
    .A1(net856),
    .A2(clknet_1_1__leaf_net899),
    .A3(net885),
    .S0(net632),
    .S1(net686),
    .X(net444));
 sky130_fd_sc_hd__mux4_1 c636 (.A0(clknet_1_0__leaf_net428),
    .A1(net627),
    .A2(net632),
    .A3(net896),
    .S0(net641),
    .S1(net751),
    .X(net445));
 sky130_fd_sc_hd__mux4_1 c637 (.A0(net876),
    .A1(clknet_1_0__leaf_net404),
    .A2(clknet_1_0__leaf_net909),
    .A3(net627),
    .S0(net632),
    .S1(net685),
    .X(net446));
 sky130_fd_sc_hd__a2111o_1 c660 (.A1(net345),
    .A2(net1026),
    .B1(net725),
    .C1(net1014),
    .D1(net970),
    .X(net447));
 sky130_fd_sc_hd__a2111o_4 c661 (.A1(net146),
    .A2(net21),
    .B1(net780),
    .C1(net1022),
    .D1(net1014),
    .X(net448));
 sky130_fd_sc_hd__a2111o_1 c662 (.A1(net141),
    .A2(net338),
    .B1(net148),
    .C1(net1022),
    .D1(net1014),
    .X(net449));
 sky130_fd_sc_hd__a2111o_1 c663 (.A1(clknet_1_1__leaf_net358),
    .A2(net447),
    .B1(net448),
    .C1(net611),
    .D1(net726),
    .X(net450));
 sky130_fd_sc_hd__a2111o_1 c664 (.A1(net970),
    .A2(net1024),
    .B1(net447),
    .C1(net337),
    .D1(net725),
    .X(net451));
 sky130_fd_sc_hd__sdfbbn_1 c665 (.CLK_N(clknet_4_15_0_clk),
    .D(net21),
    .RESET_B(net141),
    .SCD(net965),
    .SCE(net1022),
    .SET_B(net691),
    .Q(net453),
    .Q_N(net452));
 sky130_fd_sc_hd__sdfbbp_1 c666 (.CLK(clknet_4_15_0_clk),
    .D(net453),
    .RESET_B(net1050),
    .SCD(net141),
    .SCE(net337),
    .SET_B(net724),
    .Q(net455),
    .Q_N(net454));
 sky130_fd_sc_hd__sdfbbn_2 c667 (.CLK_N(clknet_4_15_0_clk),
    .D(net451),
    .RESET_B(net455),
    .SCD(net447),
    .SCE(net452),
    .SET_B(net1067),
    .Q(net457),
    .Q_N(net456));
 sky130_fd_sc_hd__a2111o_1 c668 (.A1(net455),
    .A2(net457),
    .B1(net451),
    .C1(net21),
    .D1(net1014),
    .X(net458));
 sky130_fd_sc_hd__a2111o_1 c669 (.A1(net338),
    .A2(net456),
    .B1(net165),
    .C1(net623),
    .D1(net691),
    .X(net459));
 sky130_fd_sc_hd__a2111o_2 c670 (.A1(net453),
    .A2(net456),
    .B1(net454),
    .C1(net459),
    .D1(net727),
    .X(net460));
 sky130_fd_sc_hd__a2111o_1 c671 (.A1(net141),
    .A2(net455),
    .B1(net452),
    .C1(net1002),
    .D1(net456),
    .X(net461));
 sky130_fd_sc_hd__mux4_2 c672 (.A0(net148),
    .A1(net447),
    .A2(net452),
    .A3(net456),
    .S0(net448),
    .S1(clknet_1_1__leaf_net646),
    .X(net462));
 sky130_fd_sc_hd__mux4_1 c673 (.A0(net447),
    .A1(net452),
    .A2(net448),
    .A3(clknet_1_0__leaf_net462),
    .S0(net1002),
    .S1(net611),
    .X(net463));
 sky130_fd_sc_hd__mux4_1 c674 (.A0(net459),
    .A1(net338),
    .A2(net455),
    .A3(net457),
    .S0(net453),
    .S1(net1002),
    .X(net464));
 sky130_fd_sc_hd__mux4_2 c675 (.A0(net464),
    .A1(clknet_1_1__leaf_net462),
    .A2(net1002),
    .A3(net451),
    .S1(net691),
    .X(net646));
 sky130_fd_sc_hd__mux4_1 c676 (.A0(net464),
    .A1(clknet_1_1__leaf_net450),
    .A2(net454),
    .A3(net460),
    .S0(net448),
    .S1(net753),
    .X(net466));
 sky130_fd_sc_hd__a2111o_1 c677 (.A1(net459),
    .A2(net456),
    .B1(net640),
    .C1(net753),
    .D1(clknet_1_0__leaf_net646),
    .X(net467));
 sky130_fd_sc_hd__or4bb_4 c678 (.A(net454),
    .B(clknet_1_0__leaf_net467),
    .C_N(clknet_1_1__leaf_net646),
    .D_N(net725),
    .X(net468));
 sky130_fd_sc_hd__a2111o_1 c679 (.A1(clknet_1_0__leaf_net462),
    .A2(net453),
    .B1(clknet_1_1__leaf_net467),
    .C1(clknet_1_1__leaf_net468),
    .D1(clknet_1_1__leaf_net358),
    .X(net469));
 sky130_fd_sc_hd__a2111o_1 c680 (.A1(net454),
    .A2(clknet_1_1__leaf_net468),
    .B1(net640),
    .C1(clknet_1_0__leaf_net646),
    .D1(net753),
    .X(net470));
 sky130_fd_sc_hd__mux4_1 c681 (.A0(net470),
    .A1(net464),
    .A2(net453),
    .A3(net964),
    .S0(net457),
    .S1(net640),
    .X(net471));
 sky130_fd_sc_hd__mux4_1 c682 (.A0(net254),
    .A1(net57),
    .A2(net460),
    .A3(net1051),
    .S0(net736),
    .S1(net753),
    .X(net472));
 sky130_fd_sc_hd__mux4_1 c683 (.A0(clknet_1_1__leaf_net375),
    .A1(net1036),
    .A2(net611),
    .A3(net1013),
    .S0(net1010),
    .S1(net1009),
    .X(net473));
 sky130_fd_sc_hd__mux4_2 c684 (.A0(net448),
    .A1(clknet_1_0__leaf_net468),
    .A2(net455),
    .A3(net1032),
    .S0(net736),
    .S1(net753),
    .X(net474));
 sky130_fd_sc_hd__mux4_2 c685 (.A0(net1000),
    .A1(net1028),
    .A2(net667),
    .A3(net727),
    .S0(net1010),
    .S1(net1009),
    .X(net475));
 sky130_fd_sc_hd__mux4_1 c686 (.A0(net996),
    .A1(clknet_1_1__leaf_net473),
    .A2(net1031),
    .A3(net623),
    .S0(net736),
    .S1(net1009),
    .X(net476));
 sky130_fd_sc_hd__mux4_1 c687 (.A0(clknet_1_0__leaf_net450),
    .A1(net966),
    .A2(net57),
    .A3(net475),
    .S0(clknet_1_1__leaf_net476),
    .S1(clknet_1_0__leaf_net473),
    .X(net477));
 sky130_fd_sc_hd__mux4_1 c688 (.A0(net475),
    .A1(clknet_1_0__leaf_net468),
    .A2(clknet_1_1__leaf_net476),
    .A3(net974),
    .S0(net668),
    .S1(net727),
    .X(net478));
 sky130_fd_sc_hd__mux4_1 c689 (.A0(clknet_1_1__leaf_net473),
    .A1(net964),
    .A2(net698),
    .A3(net726),
    .S0(net731),
    .S1(net736),
    .X(net479));
 sky130_fd_sc_hd__mux4_1 c690 (.A0(net964),
    .A1(net455),
    .A2(net1036),
    .A3(clknet_1_1__leaf_net476),
    .S0(net649),
    .S1(net1009),
    .X(net480));
 sky130_fd_sc_hd__mux4_1 c691 (.A0(net457),
    .A1(net475),
    .A2(net970),
    .A3(net698),
    .S0(net1009),
    .S1(clknet_1_0__leaf_net757),
    .X(net481));
 sky130_fd_sc_hd__mux4_1 c692 (.A0(clknet_1_1__leaf_net481),
    .A1(net448),
    .A2(clknet_1_1__leaf_net476),
    .A3(net965),
    .S0(net733),
    .S1(net736),
    .X(net482));
 sky130_fd_sc_hd__mux4_1 c693 (.A0(net259),
    .A1(net345),
    .A2(net160),
    .A3(clknet_1_1__leaf_net476),
    .S0(net57),
    .S1(clknet_1_0__leaf_net757),
    .X(net483));
 sky130_fd_sc_hd__mux4_1 c694 (.A0(clknet_1_0__leaf_net474),
    .A1(net448),
    .A2(net649),
    .A3(net731),
    .S0(net755),
    .S1(clknet_1_0__leaf_net757),
    .X(net484));
 sky130_fd_sc_hd__mux4_1 c695 (.A0(clknet_1_0__leaf_net468),
    .A1(clknet_1_1__leaf_net375),
    .A2(clknet_1_1__leaf_net484),
    .A3(clknet_1_1__leaf_net481),
    .S0(clknet_1_1__leaf_net476),
    .S1(clknet_1_1__leaf_net757),
    .X(net485));
 sky130_fd_sc_hd__mux4_1 c696 (.A0(net460),
    .A1(clknet_1_0__leaf_net473),
    .A2(clknet_1_1__leaf_net361),
    .A3(net456),
    .S0(net639),
    .S1(net759),
    .X(net486));
 sky130_fd_sc_hd__mux4_2 c697 (.A0(net807),
    .A1(clknet_1_1__leaf_net474),
    .A2(net1000),
    .A3(net727),
    .S0(clknet_1_0__leaf_net757),
    .S1(clknet_1_1__leaf_net758),
    .X(net487));
 sky130_fd_sc_hd__mux4_1 c698 (.A0(clknet_1_1__leaf_net486),
    .A1(net475),
    .A2(clknet_1_1__leaf_net476),
    .A3(net1032),
    .S0(clknet_1_0__leaf_net487),
    .S1(net639),
    .X(net488));
 sky130_fd_sc_hd__mux4_2 c699 (.A0(net457),
    .A1(clknet_1_0__leaf_net487),
    .A2(clknet_1_1__leaf_net481),
    .A3(net755),
    .S0(clknet_1_1__leaf_net758),
    .S1(net761),
    .X(net489));
 sky130_fd_sc_hd__mux4_2 c700 (.A0(clknet_1_1__leaf_net484),
    .A1(net475),
    .A2(net996),
    .A3(clknet_1_0__leaf_net489),
    .S0(net1010),
    .S1(net759),
    .X(net490));
 sky130_fd_sc_hd__mux4_1 c701 (.A0(clknet_1_1__leaf_net489),
    .A1(clknet_1_1__leaf_net487),
    .A2(clknet_1_1__leaf_net476),
    .A3(net623),
    .S0(net754),
    .S1(clknet_1_1__leaf_net757),
    .X(net491));
 sky130_fd_sc_hd__mux4_1 c702 (.A0(clknet_1_0__leaf_net489),
    .A1(net460),
    .A2(clknet_1_1__leaf_net476),
    .A3(net726),
    .S0(clknet_1_1__leaf_net757),
    .S1(net760),
    .X(net492));
 sky130_fd_sc_hd__mux4_1 c703 (.A0(clknet_1_1__leaf_net487),
    .A1(clknet_1_1__leaf_net489),
    .A2(net649),
    .A3(net755),
    .S0(clknet_1_1__leaf_net756),
    .S1(net763),
    .X(net493));
 sky130_fd_sc_hd__mux4_1 c704 (.A0(net1030),
    .A1(clknet_1_1__leaf_net404),
    .A2(net649),
    .A3(net1021),
    .S0(net888),
    .S1(net1009),
    .X(net494));
 sky130_fd_sc_hd__mux4_1 c705 (.A0(net1032),
    .A1(clknet_1_1__leaf_net404),
    .A2(net1030),
    .A3(clknet_1_1__leaf_net375),
    .S0(net1010),
    .S1(net736),
    .X(net495));
 sky130_fd_sc_hd__mux4_1 c706 (.A0(clknet_1_0__leaf_net495),
    .A1(clknet_1_1__leaf_net494),
    .A2(net454),
    .A3(clknet_1_0__leaf_net476),
    .S0(clknet_1_1__leaf_net701),
    .S1(net763),
    .X(net496));
 sky130_fd_sc_hd__mux4_1 c707 (.A0(clknet_1_1__leaf_net495),
    .A1(clknet_1_0__leaf_net481),
    .A2(net1010),
    .A3(clknet_1_1__leaf_net740),
    .S0(net754),
    .S1(net755),
    .X(net497));
 sky130_fd_sc_hd__mux4_1 c708 (.A0(net52),
    .A1(clknet_1_0__leaf_net917),
    .A2(clknet_1_1__leaf_net494),
    .A3(net668),
    .S0(clknet_1_0__leaf_net740),
    .S1(net755),
    .X(net498));
 sky130_fd_sc_hd__mux4_1 c709 (.A0(clknet_1_1__leaf_net495),
    .A1(clknet_1_1__leaf_net402),
    .A2(net457),
    .A3(clknet_1_1__leaf_net497),
    .S0(net595),
    .S1(net644),
    .X(net499));
 sky130_fd_sc_hd__mux4_1 c710 (.A0(net1051),
    .A1(net456),
    .A2(net644),
    .A3(clknet_1_1__leaf_net701),
    .S0(clknet_1_1__leaf_net758),
    .S1(net760),
    .X(net500));
 sky130_fd_sc_hd__mux4_1 c711 (.A0(clknet_1_0__leaf_net494),
    .A1(net57),
    .A2(net1006),
    .A3(clknet_1_1__leaf_net917),
    .S0(net595),
    .S1(net762),
    .X(net501));
 sky130_fd_sc_hd__mux4_1 c712 (.A0(clknet_1_0__leaf_net481),
    .A1(net644),
    .A2(clknet_1_1__leaf_net740),
    .A3(net1009),
    .S0(net755),
    .S1(net760),
    .X(net502));
 sky130_fd_sc_hd__mux4_1 c713 (.A0(clknet_1_1__leaf_net502),
    .A1(clknet_1_1__leaf_net495),
    .A2(clknet_1_0__leaf_net361),
    .A3(net755),
    .S0(net765),
    .S1(net766),
    .X(net503));
 sky130_fd_sc_hd__mux4_1 c714 (.A0(net457),
    .A1(clknet_1_0__leaf_net484),
    .A2(net888),
    .A3(net759),
    .S0(net764),
    .S1(net767),
    .X(net504));
 sky130_fd_sc_hd__mux4_1 c715 (.A0(net69),
    .A1(net965),
    .A2(clknet_1_1__leaf_net502),
    .A3(net732),
    .S0(net767),
    .S1(net768),
    .X(net505));
 sky130_fd_sc_hd__mux4_1 c716 (.A0(clknet_1_0__leaf_net504),
    .A1(net973),
    .A2(net1002),
    .A3(net595),
    .S0(net610),
    .S1(net768),
    .X(net506));
 sky130_fd_sc_hd__mux4_1 c717 (.A0(net595),
    .A1(net610),
    .A2(clknet_1_1__leaf_net701),
    .A3(clknet_1_1__leaf_net740),
    .S0(net753),
    .S1(net768),
    .X(net507));
 sky130_fd_sc_hd__mux4_1 c718 (.A0(clknet_1_1__leaf_net504),
    .A1(clknet_1_1__leaf_net402),
    .A2(clknet_1_1__leaf_net494),
    .A3(net1002),
    .S0(net1009),
    .S1(net767),
    .X(net508));
 sky130_fd_sc_hd__mux4_1 c719 (.A0(clknet_1_0__leaf_net497),
    .A1(net508),
    .A2(clknet_1_1__leaf_net917),
    .A3(clknet_1_1__leaf_net506),
    .S0(net764),
    .S1(net768),
    .X(net509));
 sky130_fd_sc_hd__mux4_1 c720 (.A0(net500),
    .A1(clknet_1_0__leaf_net484),
    .A2(clknet_1_1__leaf_net502),
    .A3(net644),
    .S0(clknet_1_1__leaf_net740),
    .S1(net767),
    .X(net510));
 sky130_fd_sc_hd__mux4_1 c721 (.A0(clknet_1_0__leaf_net506),
    .A1(net69),
    .A2(clknet_1_0__leaf_net495),
    .A3(net610),
    .S0(net733),
    .S1(net770),
    .X(net511));
 sky130_fd_sc_hd__mux4_1 c722 (.A0(net507),
    .A1(clknet_1_1__leaf_net511),
    .A2(clknet_1_0__leaf_net476),
    .A3(net823),
    .S0(net768),
    .S1(net878),
    .X(net512));
 sky130_fd_sc_hd__mux4_1 c723 (.A0(net1032),
    .A1(clknet_1_0__leaf_net504),
    .A2(clknet_1_0__leaf_net511),
    .A3(net52),
    .S0(clknet_1_1__leaf_net506),
    .S1(net764),
    .X(net513));
 sky130_fd_sc_hd__mux4_1 c724 (.A0(net1051),
    .A1(clknet_1_0__leaf_net506),
    .A2(clknet_1_0__leaf_net511),
    .A3(net755),
    .S0(net767),
    .S1(net768),
    .X(net514));
 sky130_fd_sc_hd__sdfbbn_1 c725 (.CLK_N(clknet_4_11_0_clk),
    .D(net69),
    .RESET_B(clknet_1_1__leaf_net511),
    .SCD(clknet_1_0__leaf_net917),
    .SCE(net639),
    .SET_B(net769),
    .Q(net516),
    .Q_N(net515));
 sky130_fd_sc_hd__mux4_1 c726 (.A0(net408),
    .A1(net455),
    .A2(net974),
    .A3(clknet_1_0__leaf_net502),
    .S0(net1002),
    .S1(net878),
    .X(net517));
 sky130_fd_sc_hd__mux4_1 c727 (.A0(net1053),
    .A1(net69),
    .A2(net674),
    .A3(net1009),
    .S0(clknet_1_1__leaf_net756),
    .S1(net770),
    .X(net518));
 sky130_fd_sc_hd__mux4_1 c728 (.A0(clknet_1_0__leaf_net476),
    .A1(net994),
    .A2(clknet_1_1__leaf_net917),
    .A3(net703),
    .S0(net765),
    .S1(net773),
    .X(net519));
 sky130_fd_sc_hd__mux4_1 c729 (.A0(clknet_1_0__leaf_net476),
    .A1(net625),
    .A2(net675),
    .A3(clknet_1_1__leaf_net701),
    .S0(clknet_1_0__leaf_net758),
    .S1(net878),
    .X(net520));
 sky130_fd_sc_hd__mux4_1 c730 (.A0(clknet_1_1__leaf_net412),
    .A1(clknet_1_0__leaf_net402),
    .A2(clknet_1_1__leaf_net917),
    .A3(clknet_1_0__leaf_net486),
    .S0(net765),
    .S1(net774),
    .X(net521));
 sky130_fd_sc_hd__mux4_1 c731 (.A0(net516),
    .A1(net678),
    .A2(net714),
    .A3(net1009),
    .S0(net761),
    .S1(net765),
    .X(net522));
 sky130_fd_sc_hd__mux4_1 c732 (.A0(clknet_1_0__leaf_net494),
    .A1(net515),
    .A2(net625),
    .A3(net678),
    .S0(net771),
    .S1(net772),
    .X(net523));
 sky130_fd_sc_hd__mux4_1 c733 (.A0(clknet_1_1__leaf_net404),
    .A1(clknet_1_1__leaf_net100),
    .A2(net454),
    .A3(net747),
    .S0(net748),
    .S1(net766),
    .X(net884));
 sky130_fd_sc_hd__mux4_1 c734 (.A0(net974),
    .A1(net965),
    .A2(clknet_1_0__leaf_net502),
    .A3(net675),
    .S0(net732),
    .S1(clknet_1_1__leaf_net756),
    .X(net524));
 sky130_fd_sc_hd__mux4_1 c735 (.A0(net522),
    .A1(clknet_1_0__leaf_net884),
    .A2(net771),
    .A3(net772),
    .S0(net773),
    .S1(net774),
    .X(net525));
 sky130_fd_sc_hd__mux4_1 c736 (.A0(clknet_1_0__leaf_net884),
    .A1(net1002),
    .A2(net974),
    .A3(net601),
    .S0(net1021),
    .S1(net748),
    .X(net526));
 sky130_fd_sc_hd__mux4_1 c737 (.A0(net518),
    .A1(net1036),
    .A2(clknet_1_1__leaf_net612),
    .A3(net713),
    .S0(net766),
    .S1(net774),
    .X(net527));
 sky130_fd_sc_hd__mux4_1 c738 (.A0(clknet_1_1__leaf_net917),
    .A1(net601),
    .A2(net747),
    .A3(net748),
    .S0(net887),
    .S1(net769),
    .X(net528));
 sky130_fd_sc_hd__mux4_1 c739 (.A0(net523),
    .A1(clknet_1_0__leaf_net527),
    .A2(net515),
    .A3(clknet_1_1__leaf_net701),
    .S0(net762),
    .S1(clknet_1_1__leaf_net945),
    .X(net529));
 sky130_fd_sc_hd__mux4_1 c740 (.A0(net516),
    .A1(clknet_1_0__leaf_net476),
    .A2(clknet_1_1__leaf_net527),
    .A3(net713),
    .S0(net762),
    .S1(net771),
    .X(net530));
 sky130_fd_sc_hd__mux4_1 c741 (.A0(net867),
    .A1(clknet_1_1__leaf_net917),
    .A2(net651),
    .A3(net766),
    .S0(net772),
    .S1(net774),
    .X(net531));
 sky130_fd_sc_hd__a2111o_1 c742 (.A1(clknet_1_0__leaf_net502),
    .A2(clknet_1_0__leaf_net404),
    .B1(net600),
    .C1(net651),
    .D1(net769),
    .X(net532));
 sky130_fd_sc_hd__mux4_1 c743 (.A0(clknet_1_1__leaf_net100),
    .A1(clknet_1_0__leaf_net494),
    .A2(net634),
    .A3(net773),
    .S0(clknet_1_0__leaf_net945),
    .S1(clknet_1_0__leaf_net883),
    .X(net533));
 sky130_fd_sc_hd__mux4_1 c744 (.A0(clknet_1_0__leaf_net533),
    .A1(net634),
    .A2(net703),
    .A3(net765),
    .S0(net772),
    .S1(clknet_1_1__leaf_net883),
    .X(net534));
 sky130_fd_sc_hd__a2111o_1 c745 (.A1(net974),
    .A2(clknet_1_0__leaf_net533),
    .B1(net600),
    .C1(net651),
    .D1(net773),
    .X(net535));
 sky130_fd_sc_hd__a2111o_1 c746 (.A1(clknet_1_1__leaf_net533),
    .A2(net622),
    .B1(net649),
    .C1(net651),
    .D1(clknet_1_0__leaf_net758),
    .X(net536));
 sky130_fd_sc_hd__mux4_1 c747 (.A0(clknet_1_1__leaf_net533),
    .A1(net965),
    .A2(net622),
    .A3(net649),
    .S0(net651),
    .S1(net772),
    .X(net537));
 sky130_fd_sc_hd__mux4_1 c748 (.A0(net1002),
    .A1(clknet_1_0__leaf_net486),
    .A2(net998),
    .A3(net854),
    .S0(net1023),
    .S1(net749),
    .X(net538));
 sky130_fd_sc_hd__mux4_1 c749 (.A0(clknet_1_0__leaf_net917),
    .A1(clknet_1_1__leaf_net612),
    .A2(net633),
    .A3(clknet_1_0__leaf_net719),
    .S0(net888),
    .S1(net749),
    .X(net539));
 sky130_fd_sc_hd__mux4_1 c750 (.A0(net1006),
    .A1(clknet_1_0__leaf_net226),
    .A2(net633),
    .A3(net1023),
    .S0(clknet_1_1__leaf_net719),
    .S1(net888),
    .X(net540));
 sky130_fd_sc_hd__mux4_1 c751 (.A0(net417),
    .A1(clknet_1_1__leaf_net701),
    .A2(net717),
    .A3(net882),
    .S0(net886),
    .S1(net769),
    .X(net541));
 sky130_fd_sc_hd__mux4_1 c752 (.A0(clknet_1_1__leaf_net446),
    .A1(clknet_1_0__leaf_net486),
    .A2(clknet_1_1__leaf_net226),
    .A3(net623),
    .S0(net633),
    .S1(clknet_1_0__leaf_net945),
    .X(net542));
 sky130_fd_sc_hd__mux4_1 c753 (.A0(net417),
    .A1(net1032),
    .A2(clknet_1_0__leaf_net446),
    .A3(net634),
    .S0(net882),
    .S1(clknet_1_0__leaf_net756),
    .X(net543));
 sky130_fd_sc_hd__mux4_1 c754 (.A0(clknet_1_0__leaf_net404),
    .A1(clknet_1_0__leaf_net908),
    .A2(net1023),
    .A3(net717),
    .S0(net750),
    .S1(clknet_1_0__leaf_net775),
    .X(net544));
 sky130_fd_sc_hd__mux4_1 c755 (.A0(net1032),
    .A1(net1021),
    .A2(net703),
    .A3(net717),
    .S0(clknet_1_1__leaf_net719),
    .S1(net882),
    .X(net879));
 sky130_fd_sc_hd__mux4_1 c756 (.A0(net541),
    .A1(clknet_1_1__leaf_net226),
    .A2(clknet_1_0__leaf_net486),
    .A3(net815),
    .S0(net623),
    .S1(clknet_1_1__leaf_net775),
    .X(net545));
 sky130_fd_sc_hd__mux4_1 c757 (.A0(clknet_1_0__leaf_net446),
    .A1(net652),
    .A2(net703),
    .A3(clknet_1_1__leaf_net719),
    .S0(clknet_1_0__leaf_net756),
    .S1(clknet_1_0__leaf_net775),
    .X(net546));
 sky130_fd_sc_hd__mux4_1 c758 (.A0(net417),
    .A1(net815),
    .A2(net882),
    .A3(net750),
    .S0(clknet_1_0__leaf_net883),
    .S1(clknet_1_0__leaf_net775),
    .X(net547));
 sky130_fd_sc_hd__mux4_1 c759 (.A0(net544),
    .A1(clknet_1_1__leaf_net908),
    .A2(net880),
    .A3(clknet_1_1__leaf_net226),
    .S0(net652),
    .S1(net776),
    .X(net548));
 sky130_fd_sc_hd__mux4_1 c760 (.A0(net516),
    .A1(clknet_1_1__leaf_net446),
    .A2(net1026),
    .A3(net652),
    .S0(clknet_1_1__leaf_net775),
    .S1(net777),
    .X(net549));
 sky130_fd_sc_hd__mux4_1 c761 (.A0(net547),
    .A1(net1005),
    .A2(clknet_1_0__leaf_net226),
    .A3(net642),
    .S0(clknet_1_1__leaf_net775),
    .S1(net777),
    .X(net550));
 sky130_fd_sc_hd__mux4_1 c762 (.A0(clknet_1_0__leaf_net527),
    .A1(clknet_1_0__leaf_net446),
    .A2(clknet_1_1__leaf_net917),
    .A3(net649),
    .S0(net717),
    .S1(net888),
    .X(net551));
 sky130_fd_sc_hd__mux4_1 c763 (.A0(clknet_1_0__leaf_net404),
    .A1(net894),
    .A2(net652),
    .A3(net750),
    .S0(net887),
    .S1(net774),
    .X(net552));
 sky130_fd_sc_hd__mux4_1 c764 (.A0(clknet_1_1__leaf_net446),
    .A1(clknet_1_1__leaf_net917),
    .A2(clknet_1_1__leaf_net226),
    .A3(net885),
    .S0(net753),
    .S1(net887),
    .X(net553));
 sky130_fd_sc_hd__mux4_1 c765 (.A0(net552),
    .A1(net815),
    .A2(clknet_1_0__leaf_net402),
    .A3(clknet_1_1__leaf_net226),
    .S0(net622),
    .S1(net777),
    .X(net554));
 sky130_fd_sc_hd__mux4_1 c766 (.A0(net1002),
    .A1(net626),
    .A2(net649),
    .A3(net746),
    .S0(net776),
    .S1(net779),
    .X(net555));
 sky130_fd_sc_hd__mux4_1 c767 (.A0(net555),
    .A1(net642),
    .A2(net886),
    .A3(net887),
    .S0(net774),
    .S1(net778),
    .X(net889));
 sky130_fd_sc_hd__mux4_1 c768 (.A0(clknet_1_0__leaf_net476),
    .A1(net880),
    .A2(clknet_1_1__leaf_net917),
    .A3(net555),
    .S0(net766),
    .S1(net778),
    .X(net556));
 sky130_fd_sc_hd__mux4_1 c769 (.A0(net555),
    .A1(net622),
    .A2(net623),
    .A3(net626),
    .S0(net776),
    .S1(net779));
 sky130_fd_sc_hd__and2_0 merge790 (.A(net472),
    .B(net479),
    .X(net557));
 sky130_fd_sc_hd__and2_0 merge791 (.A(net371),
    .B(net381),
    .X(net558));
 sky130_fd_sc_hd__dfrbp_1 merge792 (.CLK(clknet_4_9_0_clk),
    .D(net395),
    .RESET_B(net401),
    .Q(net560),
    .Q_N(net559));
 sky130_fd_sc_hd__and2_0 merge793 (.A(net513),
    .B(net514),
    .X(net561));
 sky130_fd_sc_hd__dfrbp_1 merge794 (.CLK(clknet_4_13_0_clk),
    .D(net346),
    .RESET_B(net350),
    .Q(net563),
    .Q_N(net562));
 sky130_fd_sc_hd__and2_0 merge795 (.A(net435),
    .B(net436),
    .X(net564));
 sky130_fd_sc_hd__and2_0 merge796 (.A(net212),
    .B(net229),
    .X(net565));
 sky130_fd_sc_hd__dfrtn_1 merge797 (.CLK_N(clknet_4_5_0_clk),
    .D(net158),
    .RESET_B(net163),
    .Q(net566));
 sky130_fd_sc_hd__and2_0 merge798 (.A(net195),
    .B(net194),
    .X(net567));
 sky130_fd_sc_hd__and2_0 merge799 (.A(net322),
    .B(net324),
    .X(net568));
 sky130_fd_sc_hd__and2_0 merge800 (.A(net296),
    .B(net285),
    .X(net569));
 sky130_fd_sc_hd__and2_0 merge801 (.A(net406),
    .B(net423),
    .X(net570));
 sky130_fd_sc_hd__and2_0 merge802 (.A(net249),
    .B(net250),
    .X(net571));
 sky130_fd_sc_hd__dfrtp_4 merge803 (.CLK(clknet_4_4_0_clk),
    .D(net101),
    .RESET_B(net83),
    .Q(net572));
 sky130_fd_sc_hd__dfrtp_4 merge804 (.CLK(clknet_4_7_0_clk),
    .D(net144),
    .RESET_B(net142),
    .Q(net573));
 sky130_fd_sc_hd__dfrtp_1 merge805 (.CLK(clknet_4_12_0_clk),
    .D(net262),
    .RESET_B(net274),
    .Q(net574));
 sky130_fd_sc_hd__and2_0 merge806 (.A(net526),
    .B(net530),
    .X(net575));
 sky130_fd_sc_hd__and2_0 merge807 (.A(net300),
    .B(net304),
    .X(net576));
 sky130_fd_sc_hd__and2_0 merge808 (.A(net108),
    .B(net113),
    .X(net577));
 sky130_fd_sc_hd__and2_0 merge809 (.A(net538),
    .B(net540),
    .X(net578));
 sky130_fd_sc_hd__and2_0 merge810 (.A(net171),
    .B(net180),
    .X(net579));
 sky130_fd_sc_hd__and2_0 merge811 (.A(net466),
    .B(net469),
    .X(net580));
 sky130_fd_sc_hd__and2_0 merge812 (.A(net71),
    .B(net75),
    .X(net581));
 sky130_fd_sc_hd__dfsbp_1 merge813 (.CLK(clknet_4_0_0_clk),
    .SET_B(net121),
    .Q(net955),
    .Q_N(net124));
 sky130_fd_sc_hd__and2_0 merge814 (.A(net117),
    .B(net118),
    .X(net583));
 sky130_fd_sc_hd__and2_0 merge815 (.A(net561),
    .B(net483),
    .X(net584));
 sky130_fd_sc_hd__dfsbp_1 merge816 (.CLK(clknet_4_7_0_clk),
    .D(net164),
    .Q(net586),
    .Q_N(net585));
 sky130_fd_sc_hd__and2_0 merge817 (.A(net534),
    .B(net531),
    .X(net587));
 sky130_fd_sc_hd__dfstp_2 merge818 (.CLK(clknet_4_1_0_clk),
    .D(net76),
    .SET_B(net583),
    .Q(net956));
 sky130_fd_sc_hd__and2_0 merge819 (.A(net565),
    .B(net183),
    .X(net588));
 sky130_fd_sc_hd__and2_0 merge820 (.A(net306),
    .B(net317),
    .X(net589));
 sky130_fd_sc_hd__and2_0 merge821 (.A(net437),
    .B(net445),
    .X(net590));
 sky130_fd_sc_hd__and2_0 merge822 (.A(net438),
    .B(net556),
    .X(net591));
 sky130_fd_sc_hd__and2_0 merge823 (.A(net439),
    .B(net551),
    .X(net592));
 sky130_fd_sc_hd__and2_0 merge824 (.A(net440),
    .B(net444),
    .X(net593));
 sky130_fd_sc_hd__and2_0 merge825 (.A(net545),
    .B(net549),
    .X(net594));
 sky130_fd_sc_hd__dfstp_1 merge826 (.CLK(clknet_4_8_0_clk),
    .D(net594),
    .SET_B(net570),
    .Q(net894));
 sky130_fd_sc_hd__dfstp_1 merge827 (.CLK(clknet_4_11_0_clk),
    .D(net493),
    .SET_B(net491),
    .Q(net595));
 sky130_fd_sc_hd__dlrbn_1 merge828 (.D(net286),
    .GATE_N(clknet_4_3_0_clk),
    .RESET_B(net410),
    .Q(net597),
    .Q_N(net596));
 sky130_fd_sc_hd__dlrbn_1 merge829 (.D(net581),
    .GATE_N(clknet_4_4_0_clk),
    .RESET_B(net90),
    .Q(net599),
    .Q_N(net598));
 sky130_fd_sc_hd__dlrbp_1 merge830 (.D(net521),
    .GATE(clknet_4_10_0_clk),
    .RESET_B(net575),
    .Q(net601),
    .Q_N(net600));
 sky130_fd_sc_hd__and2_0 merge831 (.A(net316),
    .B(net313),
    .X(net602));
 sky130_fd_sc_hd__and2_0 merge832 (.A(net289),
    .B(net333),
    .X(net603));
 sky130_fd_sc_hd__dlrbp_1 merge833 (.D(net571),
    .GATE(clknet_4_13_0_clk),
    .RESET_B(net364),
    .Q(net605),
    .Q_N(net604));
 sky130_fd_sc_hd__and2_0 merge834 (.A(net185),
    .B(net294),
    .X(net606));
 sky130_fd_sc_hd__dlrtn_1 merge835 (.D(net261),
    .GATE_N(clknet_4_6_0_clk),
    .RESET_B(net276),
    .Q(net607));
 sky130_fd_sc_hd__dlrtn_2 merge836 (.D(net231),
    .GATE_N(clknet_4_7_0_clk),
    .RESET_B(net238),
    .Q(net608));
 sky130_fd_sc_hd__dlrtn_1 merge837 (.D(net104),
    .GATE_N(clknet_4_0_0_clk),
    .RESET_B(net112),
    .Q(net937));
 sky130_fd_sc_hd__dlrtp_2 merge838 (.D(net290),
    .GATE(clknet_4_12_0_clk),
    .RESET_B(net253),
    .Q(net609));
 sky130_fd_sc_hd__dlrtp_2 merge839 (.D(net207),
    .GATE(clknet_4_1_0_clk),
    .RESET_B(net94),
    .Q(net934));
 sky130_fd_sc_hd__dlrtp_1 merge840 (.D(net592),
    .GATE(clknet_4_8_0_clk),
    .RESET_B(net591),
    .Q(net885));
 sky130_fd_sc_hd__edfxbp_1 merge841 (.CLK(clknet_4_14_0_clk),
    .D(net449),
    .DE(net505),
    .Q(net611),
    .Q_N(net610));
 sky130_fd_sc_hd__edfxtp_1 merge842 (.CLK(clknet_4_0_0_clk),
    .D(net577),
    .DE(net122),
    .Q(net954));
 sky130_fd_sc_hd__sdlclkp_1 merge843 (.CLK(clknet_4_8_0_clk),
    .GATE(net519),
    .SCE(net307),
    .GCLK(net612));
 sky130_fd_sc_hd__sdlclkp_2 merge844 (.CLK(clknet_4_6_0_clk),
    .GATE(net167),
    .SCE(net188),
    .GCLK(net613));
 sky130_fd_sc_hd__sdlclkp_4 merge845 (.CLK(clknet_4_1_0_clk),
    .GATE(net202),
    .SCE(net181),
    .GCLK(net614));
 sky130_fd_sc_hd__dfrbp_2 merge846 (.CLK(clknet_4_5_0_clk),
    .D(net60),
    .RESET_B(net77),
    .Q(net616),
    .Q_N(net615));
 sky130_fd_sc_hd__and2_0 merge847 (.A(net429),
    .B(net442),
    .X(net617));
 sky130_fd_sc_hd__dfrbp_1 merge848 (.CLK(clknet_4_2_0_clk),
    .D(net329),
    .RESET_B(net327),
    .Q(net618),
    .Q_N(net900));
 sky130_fd_sc_hd__and2_0 merge849 (.A(net310),
    .B(net308),
    .X(net619));
 sky130_fd_sc_hd__and2_0 merge850 (.A(net539),
    .B(net578),
    .X(net620));
 sky130_fd_sc_hd__dfrtn_1 merge851 (.CLK_N(clknet_4_8_0_clk),
    .D(net590),
    .RESET_B(net309),
    .Q(net890));
 sky130_fd_sc_hd__and2_0 merge852 (.A(net542),
    .B(net587),
    .X(net621));
 sky130_fd_sc_hd__dfrtp_1 merge853 (.CLK(clknet_4_10_0_clk),
    .D(net535),
    .RESET_B(net553),
    .Q(net622));
 sky130_fd_sc_hd__dfrtp_4 merge854 (.CLK(clknet_4_4_0_clk),
    .D(net606),
    .RESET_B(net579),
    .Q(net947));
 sky130_fd_sc_hd__dfrtp_4 merge855 (.CLK(clknet_4_15_0_clk),
    .D(net458),
    .RESET_B(net537),
    .Q(net623));
 sky130_fd_sc_hd__dfsbp_1 merge856 (.CLK(clknet_4_3_0_clk),
    .D(net422),
    .SET_B(net569),
    .Q(net625),
    .Q_N(net624));
 sky130_fd_sc_hd__dfsbp_1 merge857 (.CLK(clknet_4_8_0_clk),
    .D(net593),
    .SET_B(net550),
    .Q(net627),
    .Q_N(net626));
 sky130_fd_sc_hd__dfstp_1 merge858 (.CLK(clknet_4_0_0_clk),
    .SET_B(net120),
    .Q(net123));
 sky130_fd_sc_hd__and2_0 merge859 (.A(net548),
    .B(net564),
    .X(net628));
 sky130_fd_sc_hd__dfstp_2 merge860 (.CLK(clknet_4_3_0_clk),
    .D(net319),
    .SET_B(net297),
    .Q(net629));
 sky130_fd_sc_hd__dfstp_2 merge861 (.CLK(clknet_4_1_0_clk),
    .D(net588),
    .SET_B(net97),
    .Q(net630));
 sky130_fd_sc_hd__dlrbn_1 merge862 (.D(net443),
    .GATE_N(clknet_4_8_0_clk),
    .RESET_B(net415),
    .Q(net632),
    .Q_N(net631));
 sky130_fd_sc_hd__dlrbn_1 merge863 (.D(net532),
    .GATE_N(clknet_4_10_0_clk),
    .RESET_B(net536),
    .Q(net634),
    .Q_N(net633));
 sky130_fd_sc_hd__dlrbp_1 merge864 (.D(net263),
    .GATE(clknet_4_12_0_clk),
    .RESET_B(net377),
    .Q(net636),
    .Q_N(net635));
 sky130_fd_sc_hd__dlrbp_1 merge865 (.D(net239),
    .GATE(clknet_4_13_0_clk),
    .RESET_B(net265),
    .Q(net638),
    .Q_N(net637));
 sky130_fd_sc_hd__dlrtn_2 merge866 (.D(net240),
    .GATE_N(clknet_4_14_0_clk),
    .RESET_B(net584),
    .Q(net639));
 sky130_fd_sc_hd__dlrtn_2 merge867 (.D(net246),
    .GATE_N(clknet_4_15_0_clk),
    .RESET_B(net580),
    .Q(net640));
 sky130_fd_sc_hd__dlrtn_2 merge868 (.D(net617),
    .GATE_N(clknet_4_3_0_clk),
    .RESET_B(net576),
    .Q(net896));
 sky130_fd_sc_hd__dlrtp_2 merge869 (.D(net332),
    .GATE(clknet_4_3_0_clk),
    .RESET_B(net209),
    .Q(net641));
 sky130_fd_sc_hd__dlrtp_4 merge870 (.D(net251),
    .GATE(clknet_4_12_0_clk),
    .RESET_B(net603),
    .Q(net915));
 sky130_fd_sc_hd__dlrtp_2 merge871 (.D(net628),
    .GATE(clknet_4_8_0_clk),
    .RESET_B(net318),
    .Q(net642));
 sky130_fd_sc_hd__edfxbp_1 merge872 (.CLK(clknet_4_3_0_clk),
    .D(net279),
    .DE(net602),
    .Q(net643),
    .Q_N(net891));
 sky130_fd_sc_hd__edfxtp_1 merge873 (.CLK(clknet_4_9_0_clk),
    .D(net498),
    .DE(net619),
    .Q(net644));
 sky130_fd_sc_hd__sdlclkp_1 merge874 (.CLK(clknet_4_6_0_clk),
    .GATE(net206),
    .SCE(net268),
    .GCLK(net933));
 sky130_fd_sc_hd__sdlclkp_2 merge875 (.CLK(clknet_4_14_0_clk),
    .GATE(net356),
    .SCE(net370),
    .GCLK(net645));
 sky130_fd_sc_hd__sdlclkp_4 merge876 (.CLK(clknet_4_15_0_clk),
    .SCE(net461),
    .GCLK(net646));
 sky130_fd_sc_hd__dfrbp_2 merge877 (.CLK(clknet_4_0_0_clk),
    .D(net119),
    .RESET_B(net225),
    .Q(net951),
    .Q_N(net950));
 sky130_fd_sc_hd__dfrbp_2 merge878 (.CLK(clknet_4_0_0_clk),
    .D(net210),
    .RESET_B(net109),
    .Q(net648),
    .Q_N(net647));
 sky130_fd_sc_hd__dfrtn_1 merge879 (.CLK_N(clknet_4_14_0_clk),
    .D(net557),
    .RESET_B(net621),
    .Q(net649));
 sky130_fd_sc_hd__dfrtp_4 merge880 (.CLK(clknet_4_3_0_clk),
    .D(net589),
    .RESET_B(net568),
    .Q(net920));
 sky130_fd_sc_hd__dfrtp_4 merge881 (.CLK(clknet_4_1_0_clk),
    .D(net184),
    .RESET_B(net567),
    .Q(net650));
 sky130_fd_sc_hd__dfrtp_2 merge882 (.CLK(clknet_4_10_0_clk),
    .D(net528),
    .RESET_B(net529),
    .Q(net651));
 sky130_fd_sc_hd__dfsbp_2 merge883 (.CLK(clknet_4_8_0_clk),
    .D(net419),
    .SET_B(net620),
    .Q(net653),
    .Q_N(net652));
 sky130_fd_sc_hd__dfsbp_2 merge884 (.CLK(clknet_4_12_0_clk),
    .D(net343),
    .SET_B(net558),
    .Q(net655),
    .Q_N(net654));
 sky130_fd_sc_hd__dfxbp_1 s885 (.CLK(clknet_4_4_0_clk),
    .D(net67),
    .Q(net657),
    .Q_N(net656));
 sky130_fd_sc_hd__dfxbp_2 s886 (.CLK(clknet_4_4_0_clk),
    .D(net72),
    .Q(net659),
    .Q_N(net658));
 sky130_fd_sc_hd__dfxtp_1 s887 (.CLK(clknet_4_5_0_clk),
    .D(net78),
    .Q(net660));
 sky130_fd_sc_hd__dfxtp_4 s888 (.CLK(clknet_4_4_0_clk),
    .D(net79),
    .Q(net661));
 sky130_fd_sc_hd__dfxtp_2 s889 (.CLK(clknet_4_5_0_clk),
    .D(net80),
    .Q(net662));
 sky130_fd_sc_hd__dlclkp_1 s890 (.CLK(clknet_4_4_0_clk),
    .GATE(net92),
    .GCLK(net924));
 sky130_fd_sc_hd__dlclkp_2 s891 (.CLK(clknet_4_1_0_clk),
    .GATE(net93),
    .GCLK(net663));
 sky130_fd_sc_hd__dlclkp_4 s892 (.CLK(clknet_4_1_0_clk),
    .GATE(net95),
    .GCLK(net664));
 sky130_fd_sc_hd__dlxbn_1 s893 (.D(net98),
    .GATE_N(clknet_4_1_0_clk),
    .Q(net666),
    .Q_N(net665));
 sky130_fd_sc_hd__dlxbn_1 s894 (.D(net143),
    .GATE_N(clknet_4_7_0_clk),
    .Q(net906),
    .Q_N(net667));
 sky130_fd_sc_hd__dlxbp_1 s895 (.D(net166),
    .GATE(clknet_4_5_0_clk),
    .Q(net898),
    .Q_N(net668));
 sky130_fd_sc_hd__dlxtn_2 s896 (.D(net168),
    .GATE_N(clknet_4_6_0_clk),
    .Q(net669));
 sky130_fd_sc_hd__dlxtn_1 s897 (.D(net175),
    .GATE_N(clknet_4_5_0_clk),
    .Q(net670));
 sky130_fd_sc_hd__dlxtn_2 s898 (.D(net176),
    .GATE_N(clknet_4_4_0_clk),
    .Q(net671));
 sky130_fd_sc_hd__dlxtp_1 s899 (.D(net177),
    .GATE(clknet_4_4_0_clk),
    .Q(net672));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s900 (.D(net178),
    .SLEEP_B(clknet_4_5_0_clk),
    .Q(net673));
 sky130_fd_sc_hd__dfxbp_2 s901 (.CLK(clknet_4_1_0_clk),
    .D(net191),
    .Q(net675),
    .Q_N(net674));
 sky130_fd_sc_hd__dfxbp_1 s902 (.CLK(clknet_4_3_0_clk),
    .D(net197),
    .Q(net677),
    .Q_N(net676));
 sky130_fd_sc_hd__dfxtp_2 s903 (.CLK(clknet_4_1_0_clk),
    .D(net201),
    .Q(net916));
 sky130_fd_sc_hd__dfxtp_4 s904 (.CLK(clknet_4_1_0_clk),
    .D(net203),
    .Q(net678));
 sky130_fd_sc_hd__dfxtp_2 s905 (.CLK(clknet_4_1_0_clk),
    .D(net204),
    .Q(net679));
 sky130_fd_sc_hd__dlclkp_1 s906 (.CLK(clknet_4_1_0_clk),
    .GATE(net205),
    .GCLK(net680));
 sky130_fd_sc_hd__dlclkp_2 s907 (.CLK(clknet_4_0_0_clk),
    .GATE(net211),
    .GCLK(net902));
 sky130_fd_sc_hd__dlclkp_4 s908 (.CLK(clknet_4_0_0_clk),
    .GATE(net213),
    .GCLK(net914));
 sky130_fd_sc_hd__dlxbn_2 s909 (.D(net223),
    .GATE_N(clknet_4_2_0_clk),
    .Q(net682),
    .Q_N(net681));
 sky130_fd_sc_hd__dlxbn_1 s910 (.D(net224),
    .GATE_N(clknet_4_2_0_clk),
    .Q(net684),
    .Q_N(net683));
 sky130_fd_sc_hd__dlxbp_1 s911 (.D(net227),
    .GATE(clknet_4_2_0_clk),
    .Q(net686),
    .Q_N(net685));
 sky130_fd_sc_hd__dlxtn_2 s912 (.D(net228),
    .GATE_N(clknet_4_2_0_clk),
    .Q(net687));
 sky130_fd_sc_hd__dlxtn_2 s913 (.D(net230),
    .GATE_N(clknet_4_2_0_clk),
    .Q(net688));
 sky130_fd_sc_hd__dlxtn_1 s914 (.D(net237),
    .GATE_N(clknet_4_7_0_clk),
    .Q(net689));
 sky130_fd_sc_hd__dlxtp_1 s915 (.D(net245),
    .GATE(clknet_4_13_0_clk),
    .Q(net690));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s916 (.D(net247),
    .SLEEP_B(clknet_4_13_0_clk),
    .Q(net691));
 sky130_fd_sc_hd__dfxbp_2 s917 (.CLK(clknet_4_12_0_clk),
    .D(net252),
    .Q(net693),
    .Q_N(net692));
 sky130_fd_sc_hd__dfxbp_1 s918 (.CLK(clknet_4_7_0_clk),
    .D(net255),
    .Q(net695),
    .Q_N(net694));
 sky130_fd_sc_hd__dfxtp_1 s919 (.CLK(clknet_4_7_0_clk),
    .D(net258),
    .Q(net696));
 sky130_fd_sc_hd__dfxtp_1 s920 (.CLK(clknet_4_12_0_clk),
    .D(net264),
    .Q(net697));
 sky130_fd_sc_hd__dfxtp_1 s921 (.CLK(clknet_4_12_0_clk),
    .D(net266),
    .Q(net698));
 sky130_fd_sc_hd__dlclkp_1 s922 (.CLK(clknet_4_12_0_clk),
    .GATE(net267),
    .GCLK(net699));
 sky130_fd_sc_hd__dlclkp_2 s923 (.CLK(clknet_4_6_0_clk),
    .GATE(net270),
    .GCLK(net700));
 sky130_fd_sc_hd__dlclkp_4 s924 (.CLK(clknet_4_6_0_clk),
    .GATE(net272),
    .GCLK(net701));
 sky130_fd_sc_hd__dlxbn_2 s925 (.D(net273),
    .GATE_N(clknet_4_12_0_clk),
    .Q(net703),
    .Q_N(net702));
 sky130_fd_sc_hd__dlxbn_1 s926 (.D(net280),
    .GATE_N(clknet_4_6_0_clk),
    .Q(net705),
    .Q_N(net704));
 sky130_fd_sc_hd__dlxbp_1 s927 (.D(net281),
    .GATE(clknet_4_6_0_clk),
    .Q(net707),
    .Q_N(net706));
 sky130_fd_sc_hd__dlxtn_1 s928 (.D(net282),
    .GATE_N(clknet_4_6_0_clk),
    .Q(net708));
 sky130_fd_sc_hd__dlxtn_2 s929 (.D(net292),
    .GATE_N(clknet_4_9_0_clk),
    .Q(net709));
 sky130_fd_sc_hd__dlxtn_1 s930 (.D(net293),
    .GATE_N(clknet_4_6_0_clk),
    .Q(net710));
 sky130_fd_sc_hd__dlxtp_1 s931 (.D(net295),
    .GATE(clknet_4_6_0_clk),
    .Q(net711));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s932 (.D(net312),
    .SLEEP_B(clknet_4_3_0_clk),
    .Q(net712));
 sky130_fd_sc_hd__dfxbp_1 s933 (.CLK(clknet_4_3_0_clk),
    .D(net314),
    .Q(net714),
    .Q_N(net713));
 sky130_fd_sc_hd__dfxbp_1 s934 (.CLK(clknet_4_2_0_clk),
    .D(net321),
    .Q(net923),
    .Q_N(net715));
 sky130_fd_sc_hd__dfxtp_1 s935 (.CLK(clknet_4_2_0_clk),
    .D(net326),
    .Q(net716));
 sky130_fd_sc_hd__dfxtp_2 s936 (.CLK(clknet_4_2_0_clk),
    .D(net334),
    .Q(net717));
 sky130_fd_sc_hd__dfxtp_2 s937 (.CLK(clknet_4_2_0_clk),
    .D(net335),
    .Q(net718));
 sky130_fd_sc_hd__dlclkp_1 s938 (.CLK(clknet_4_2_0_clk),
    .GATE(net336),
    .GCLK(net719));
 sky130_fd_sc_hd__dlclkp_2 s939 (.CLK(clknet_4_13_0_clk),
    .GATE(net347),
    .GCLK(net720));
 sky130_fd_sc_hd__dlclkp_4 s940 (.CLK(clknet_4_15_0_clk),
    .GATE(net348),
    .GCLK(net721));
 sky130_fd_sc_hd__dlxbn_1 s941 (.D(net349),
    .GATE_N(clknet_4_15_0_clk),
    .Q(net723),
    .Q_N(net722));
 sky130_fd_sc_hd__dlxbn_2 s942 (.D(net352),
    .GATE_N(clknet_4_15_0_clk),
    .Q(net725),
    .Q_N(net724));
 sky130_fd_sc_hd__dlxbp_1 s943 (.D(net353),
    .GATE(clknet_4_15_0_clk),
    .Q(net727),
    .Q_N(net726));
 sky130_fd_sc_hd__dlxtn_1 s944 (.D(net357),
    .GATE_N(clknet_4_13_0_clk),
    .Q(net728));
 sky130_fd_sc_hd__dlxtn_4 s945 (.D(net359),
    .GATE_N(clknet_4_15_0_clk),
    .Q(net904));
 sky130_fd_sc_hd__dlxtn_2 s946 (.D(net363),
    .GATE_N(clknet_4_12_0_clk),
    .Q(net729));
 sky130_fd_sc_hd__dlxtp_1 s947 (.D(net374),
    .GATE(clknet_4_12_0_clk),
    .Q(net730));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s948 (.D(net378),
    .SLEEP_B(clknet_4_14_0_clk),
    .Q(net731));
 sky130_fd_sc_hd__dfxbp_2 s949 (.CLK(clknet_4_14_0_clk),
    .D(net380),
    .Q(net733),
    .Q_N(net732));
 sky130_fd_sc_hd__dfxbp_1 s950 (.CLK(clknet_4_9_0_clk),
    .D(net382),
    .Q(net735),
    .Q_N(net734));
 sky130_fd_sc_hd__dfxtp_2 s951 (.CLK(clknet_4_14_0_clk),
    .D(net383),
    .Q(net736));
 sky130_fd_sc_hd__dfxtp_4 s952 (.CLK(clknet_4_9_0_clk),
    .D(net390),
    .Q(net888));
 sky130_fd_sc_hd__dfxtp_1 s953 (.CLK(clknet_4_9_0_clk),
    .D(net393),
    .Q(net737));
 sky130_fd_sc_hd__dlclkp_1 s954 (.CLK(clknet_4_9_0_clk),
    .GATE(net396),
    .GCLK(net738));
 sky130_fd_sc_hd__dlclkp_2 s955 (.CLK(clknet_4_9_0_clk),
    .GATE(net397),
    .GCLK(net739));
 sky130_fd_sc_hd__dlclkp_4 s956 (.CLK(clknet_4_9_0_clk),
    .GATE(net398),
    .GCLK(net740));
 sky130_fd_sc_hd__dlxbn_1 s957 (.D(net403),
    .GATE_N(clknet_4_9_0_clk),
    .Q(net742),
    .Q_N(net741));
 sky130_fd_sc_hd__dlxbn_1 s958 (.D(net409),
    .GATE_N(clknet_4_8_0_clk),
    .Q(net903),
    .Q_N(net743));
 sky130_fd_sc_hd__dlxbp_1 s959 (.D(net411),
    .GATE(clknet_4_9_0_clk),
    .Q(net745),
    .Q_N(net744));
 sky130_fd_sc_hd__dlxtn_2 s960 (.D(net414),
    .GATE_N(clknet_4_9_0_clk),
    .Q(net746));
 sky130_fd_sc_hd__dlxtn_2 s961 (.D(net416),
    .GATE_N(clknet_4_8_0_clk),
    .Q(net747));
 sky130_fd_sc_hd__dlxtn_1 s962 (.D(net418),
    .GATE_N(clknet_4_8_0_clk),
    .Q(net748));
 sky130_fd_sc_hd__dlxtp_1 s963 (.D(net425),
    .GATE(clknet_4_8_0_clk),
    .Q(net882));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s964 (.D(net427),
    .SLEEP_B(clknet_4_8_0_clk),
    .Q(net886));
 sky130_fd_sc_hd__dfxbp_1 s965 (.CLK(clknet_4_8_0_clk),
    .D(net433),
    .Q(net750),
    .Q_N(net749));
 sky130_fd_sc_hd__dfxbp_1 s966 (.CLK(clknet_4_8_0_clk),
    .D(net434),
    .Q(net752),
    .Q_N(net751));
 sky130_fd_sc_hd__dfxtp_2 s967 (.CLK(clknet_4_14_0_clk),
    .D(net463),
    .Q(net753));
 sky130_fd_sc_hd__dfxtp_1 s968 (.CLK(clknet_4_14_0_clk),
    .D(net471),
    .Q(net754));
 sky130_fd_sc_hd__dfxtp_2 s969 (.CLK(clknet_4_14_0_clk),
    .D(net477),
    .Q(net755));
 sky130_fd_sc_hd__dlclkp_1 s970 (.CLK(clknet_4_11_0_clk),
    .GATE(net478),
    .GCLK(net756));
 sky130_fd_sc_hd__dlclkp_2 s971 (.CLK(clknet_4_14_0_clk),
    .GATE(net480),
    .GCLK(net757));
 sky130_fd_sc_hd__dlclkp_4 s972 (.CLK(clknet_4_14_0_clk),
    .GATE(net482),
    .GCLK(net758));
 sky130_fd_sc_hd__dlxbn_1 s973 (.D(net485),
    .GATE_N(clknet_4_14_0_clk),
    .Q(net760),
    .Q_N(net759));
 sky130_fd_sc_hd__dlxbn_1 s974 (.D(net488),
    .GATE_N(clknet_4_11_0_clk),
    .Q(net762),
    .Q_N(net761));
 sky130_fd_sc_hd__dlxbp_1 s975 (.D(net490),
    .GATE(clknet_4_11_0_clk),
    .Q(net764),
    .Q_N(net763));
 sky130_fd_sc_hd__dlxtn_2 s976 (.D(net492),
    .GATE_N(clknet_4_11_0_clk),
    .Q(net765));
 sky130_fd_sc_hd__dlxtn_2 s977 (.D(net496),
    .GATE_N(clknet_4_11_0_clk),
    .Q(net766));
 sky130_fd_sc_hd__dlxtn_1 s978 (.D(net499),
    .GATE_N(clknet_4_11_0_clk),
    .Q(net767));
 sky130_fd_sc_hd__dlxtp_1 s979 (.D(net501),
    .GATE(clknet_4_11_0_clk),
    .Q(net887));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s980 (.D(net503),
    .SLEEP_B(clknet_4_11_0_clk),
    .Q(net768));
 sky130_fd_sc_hd__dfxbp_2 s981 (.CLK(clknet_4_11_0_clk),
    .D(net509),
    .Q(net878),
    .Q_N(net769));
 sky130_fd_sc_hd__dfxbp_1 s982 (.CLK(clknet_4_11_0_clk),
    .D(net510),
    .Q(net771),
    .Q_N(net770));
 sky130_fd_sc_hd__dfxtp_1 s983 (.CLK(clknet_4_11_0_clk),
    .D(net512),
    .Q(net772));
 sky130_fd_sc_hd__dfxtp_1 s984 (.CLK(clknet_4_10_0_clk),
    .D(net517),
    .Q(net773));
 sky130_fd_sc_hd__dfxtp_2 s985 (.CLK(clknet_4_10_0_clk),
    .D(net520),
    .Q(net774));
 sky130_fd_sc_hd__dlclkp_1 s986 (.CLK(clknet_4_10_0_clk),
    .GATE(net524),
    .GCLK(net945));
 sky130_fd_sc_hd__dlclkp_2 s987 (.CLK(clknet_4_10_0_clk),
    .GATE(net525),
    .GCLK(net883));
 sky130_fd_sc_hd__dlclkp_4 s988 (.CLK(clknet_4_10_0_clk),
    .GATE(net543),
    .GCLK(net775));
 sky130_fd_sc_hd__dlxbn_1 s989 (.D(net546),
    .GATE_N(clknet_4_8_0_clk),
    .Q(net777),
    .Q_N(net776));
 sky130_fd_sc_hd__dlxbn_1 s990 (.D(net554),
    .GATE_N(clknet_4_10_0_clk),
    .Q(net779),
    .Q_N(net778));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Right_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Right_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Right_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Right_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Right_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Right_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Right_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Right_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Right_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Right_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Right_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Right_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Right_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Right_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Right_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Right_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Right_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Right_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Right_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Right_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Right_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_161 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_162 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_163 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_164 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_165 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_166 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_167 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_168 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_169 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_170 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_171 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_172 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_173 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_174 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_175 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_176 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_177 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_178 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_179 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_180 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_181 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_182 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Left_183 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Left_184 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Left_185 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Left_186 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Left_187 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Left_188 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Left_189 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Left_190 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Left_191 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Left_192 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Left_193 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Left_194 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Left_195 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Left_196 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Left_197 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Left_198 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Left_199 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Left_200 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Left_201 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Left_202 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Left_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1347 ();
 sky130_fd_sc_hd__buf_2 input1 (.A(in0),
    .X(net165));
 sky130_fd_sc_hd__dlymetal6s2s_1 input2 (.A(in1),
    .X(net465));
 sky130_fd_sc_hd__clkbuf_2 input3 (.A(in10),
    .X(net780));
 sky130_fd_sc_hd__buf_2 input4 (.A(in11),
    .X(net781));
 sky130_fd_sc_hd__clkbuf_2 input5 (.A(in12),
    .X(net782));
 sky130_fd_sc_hd__buf_1 input6 (.A(in13),
    .X(net783));
 sky130_fd_sc_hd__clkbuf_2 input7 (.A(in14),
    .X(net784));
 sky130_fd_sc_hd__clkbuf_2 input8 (.A(in15),
    .X(net785));
 sky130_fd_sc_hd__buf_2 input9 (.A(in16),
    .X(net786));
 sky130_fd_sc_hd__dlymetal6s2s_1 input10 (.A(in17),
    .X(net787));
 sky130_fd_sc_hd__clkbuf_2 input11 (.A(in18),
    .X(net788));
 sky130_fd_sc_hd__buf_1 input12 (.A(in19),
    .X(net789));
 sky130_fd_sc_hd__buf_8 input13 (.A(in2),
    .X(net790));
 sky130_fd_sc_hd__dlymetal6s2s_1 input14 (.A(in20),
    .X(net791));
 sky130_fd_sc_hd__buf_1 input15 (.A(in21),
    .X(net792));
 sky130_fd_sc_hd__buf_4 input16 (.A(in22),
    .X(net793));
 sky130_fd_sc_hd__buf_1 input17 (.A(in23),
    .X(net794));
 sky130_fd_sc_hd__buf_1 input18 (.A(in24),
    .X(net795));
 sky130_fd_sc_hd__clkbuf_2 input19 (.A(in25),
    .X(net796));
 sky130_fd_sc_hd__buf_1 input20 (.A(in26),
    .X(net797));
 sky130_fd_sc_hd__buf_1 input21 (.A(in27),
    .X(net798));
 sky130_fd_sc_hd__clkbuf_1 input22 (.A(in28),
    .X(net799));
 sky130_fd_sc_hd__buf_1 input23 (.A(in29),
    .X(net800));
 sky130_fd_sc_hd__clkbuf_2 input24 (.A(in3),
    .X(net801));
 sky130_fd_sc_hd__clkbuf_4 input25 (.A(in30),
    .X(net802));
 sky130_fd_sc_hd__buf_1 input26 (.A(in31),
    .X(net803));
 sky130_fd_sc_hd__clkbuf_2 input27 (.A(in32),
    .X(net804));
 sky130_fd_sc_hd__dlymetal6s2s_1 input28 (.A(in33),
    .X(net805));
 sky130_fd_sc_hd__buf_1 input29 (.A(in34),
    .X(net806));
 sky130_fd_sc_hd__clkbuf_2 input30 (.A(in35),
    .X(net807));
 sky130_fd_sc_hd__buf_4 input31 (.A(in36),
    .X(net808));
 sky130_fd_sc_hd__clkbuf_2 input32 (.A(in37),
    .X(net809));
 sky130_fd_sc_hd__clkbuf_4 input33 (.A(in38),
    .X(net810));
 sky130_fd_sc_hd__clkbuf_4 input34 (.A(in39),
    .X(net811));
 sky130_fd_sc_hd__dlymetal6s2s_1 input35 (.A(in4),
    .X(net812));
 sky130_fd_sc_hd__clkbuf_4 input36 (.A(in40),
    .X(net813));
 sky130_fd_sc_hd__clkbuf_2 input37 (.A(in41),
    .X(net814));
 sky130_fd_sc_hd__clkbuf_4 input38 (.A(in42),
    .X(net815));
 sky130_fd_sc_hd__clkbuf_2 input39 (.A(in43),
    .X(net816));
 sky130_fd_sc_hd__buf_2 input40 (.A(in44),
    .X(net817));
 sky130_fd_sc_hd__buf_1 input41 (.A(in45),
    .X(net818));
 sky130_fd_sc_hd__clkbuf_2 input42 (.A(in46),
    .X(net819));
 sky130_fd_sc_hd__clkbuf_4 input43 (.A(in47),
    .X(net820));
 sky130_fd_sc_hd__buf_1 input44 (.A(in48),
    .X(net821));
 sky130_fd_sc_hd__clkbuf_1 input45 (.A(in49),
    .X(net822));
 sky130_fd_sc_hd__clkbuf_2 input46 (.A(in5),
    .X(net823));
 sky130_fd_sc_hd__dlymetal6s2s_1 input47 (.A(in50),
    .X(net824));
 sky130_fd_sc_hd__clkbuf_2 input48 (.A(in51),
    .X(net825));
 sky130_fd_sc_hd__buf_2 input49 (.A(in52),
    .X(net826));
 sky130_fd_sc_hd__clkbuf_4 input50 (.A(in53),
    .X(net827));
 sky130_fd_sc_hd__clkbuf_2 input51 (.A(in54),
    .X(net828));
 sky130_fd_sc_hd__buf_2 input52 (.A(in55),
    .X(net829));
 sky130_fd_sc_hd__clkbuf_1 input53 (.A(in56),
    .X(net830));
 sky130_fd_sc_hd__buf_1 input54 (.A(in57),
    .X(net831));
 sky130_fd_sc_hd__clkbuf_2 input55 (.A(in58),
    .X(net832));
 sky130_fd_sc_hd__clkbuf_2 input56 (.A(in59),
    .X(net833));
 sky130_fd_sc_hd__buf_1 input57 (.A(in6),
    .X(net834));
 sky130_fd_sc_hd__buf_1 input58 (.A(in60),
    .X(net835));
 sky130_fd_sc_hd__clkbuf_1 input59 (.A(in61),
    .X(net836));
 sky130_fd_sc_hd__buf_2 input60 (.A(in62),
    .X(net837));
 sky130_fd_sc_hd__buf_1 input61 (.A(in63),
    .X(net838));
 sky130_fd_sc_hd__buf_2 input62 (.A(in64),
    .X(net839));
 sky130_fd_sc_hd__buf_1 input63 (.A(in65),
    .X(net840));
 sky130_fd_sc_hd__dlymetal6s2s_1 input64 (.A(in66),
    .X(net841));
 sky130_fd_sc_hd__buf_1 input65 (.A(in67),
    .X(net842));
 sky130_fd_sc_hd__buf_2 input66 (.A(in68),
    .X(net843));
 sky130_fd_sc_hd__clkbuf_1 input67 (.A(in69),
    .X(net844));
 sky130_fd_sc_hd__buf_2 input68 (.A(in7),
    .X(net845));
 sky130_fd_sc_hd__clkbuf_2 input69 (.A(in70),
    .X(net846));
 sky130_fd_sc_hd__clkbuf_1 input70 (.A(in71),
    .X(net847));
 sky130_fd_sc_hd__buf_4 input71 (.A(in72),
    .X(net848));
 sky130_fd_sc_hd__clkbuf_4 input72 (.A(in73),
    .X(net849));
 sky130_fd_sc_hd__clkbuf_1 input73 (.A(in74),
    .X(net850));
 sky130_fd_sc_hd__clkbuf_1 input74 (.A(in75),
    .X(net851));
 sky130_fd_sc_hd__clkbuf_1 input75 (.A(in76),
    .X(net852));
 sky130_fd_sc_hd__clkbuf_1 input76 (.A(in77),
    .X(net853));
 sky130_fd_sc_hd__clkbuf_4 input77 (.A(in78),
    .X(net854));
 sky130_fd_sc_hd__clkbuf_4 input78 (.A(in79),
    .X(net855));
 sky130_fd_sc_hd__buf_2 input79 (.A(in8),
    .X(net856));
 sky130_fd_sc_hd__buf_1 input80 (.A(in80),
    .X(net857));
 sky130_fd_sc_hd__clkbuf_1 input81 (.A(in81),
    .X(net858));
 sky130_fd_sc_hd__buf_1 input82 (.A(in82),
    .X(net859));
 sky130_fd_sc_hd__clkbuf_1 input83 (.A(in83),
    .X(net860));
 sky130_fd_sc_hd__buf_1 input84 (.A(in84),
    .X(net861));
 sky130_fd_sc_hd__clkbuf_1 input85 (.A(in85),
    .X(net862));
 sky130_fd_sc_hd__buf_1 input86 (.A(in86),
    .X(net863));
 sky130_fd_sc_hd__clkbuf_4 input87 (.A(in87),
    .X(net864));
 sky130_fd_sc_hd__clkbuf_4 input88 (.A(in88),
    .X(net865));
 sky130_fd_sc_hd__clkbuf_2 input89 (.A(in89),
    .X(net866));
 sky130_fd_sc_hd__buf_6 input90 (.A(in9),
    .X(net867));
 sky130_fd_sc_hd__buf_1 input91 (.A(in90),
    .X(net868));
 sky130_fd_sc_hd__buf_1 input92 (.A(in91),
    .X(net869));
 sky130_fd_sc_hd__buf_1 input93 (.A(in92),
    .X(net870));
 sky130_fd_sc_hd__buf_2 input94 (.A(in93),
    .X(net871));
 sky130_fd_sc_hd__clkbuf_2 input95 (.A(in94),
    .X(net872));
 sky130_fd_sc_hd__buf_1 input96 (.A(in95),
    .X(net873));
 sky130_fd_sc_hd__dlymetal6s2s_1 input97 (.A(in96),
    .X(net874));
 sky130_fd_sc_hd__clkbuf_2 input98 (.A(in97),
    .X(net875));
 sky130_fd_sc_hd__clkbuf_4 input99 (.A(in98),
    .X(net876));
 sky130_fd_sc_hd__buf_1 input100 (.A(in99),
    .X(net877));
 sky130_fd_sc_hd__buf_2 output101 (.A(net878),
    .X(out0));
 sky130_fd_sc_hd__clkbuf_1 output102 (.A(net879),
    .X(out1));
 sky130_fd_sc_hd__buf_2 output103 (.A(net880),
    .X(out10));
 sky130_fd_sc_hd__buf_2 output104 (.A(net881),
    .X(out12));
 sky130_fd_sc_hd__buf_2 output105 (.A(net882),
    .X(out13));
 sky130_fd_sc_hd__clkbuf_1 output106 (.A(clknet_1_1__leaf_net883),
    .X(out14));
 sky130_fd_sc_hd__clkbuf_1 output107 (.A(clknet_1_1__leaf_net884),
    .X(out15));
 sky130_fd_sc_hd__buf_2 output108 (.A(net885),
    .X(out16));
 sky130_fd_sc_hd__buf_2 output109 (.A(net886),
    .X(out17));
 sky130_fd_sc_hd__buf_2 output110 (.A(net887),
    .X(out18));
 sky130_fd_sc_hd__buf_2 output111 (.A(net888),
    .X(out19));
 sky130_fd_sc_hd__buf_2 output112 (.A(net889),
    .X(out2));
 sky130_fd_sc_hd__buf_2 output113 (.A(net890),
    .X(out20));
 sky130_fd_sc_hd__buf_2 output114 (.A(net891),
    .X(out21));
 sky130_fd_sc_hd__clkbuf_1 output115 (.A(clknet_1_0__leaf_net892),
    .X(out22));
 sky130_fd_sc_hd__clkbuf_1 output116 (.A(clknet_1_0__leaf_net893),
    .X(out23));
 sky130_fd_sc_hd__buf_2 output117 (.A(net894),
    .X(out24));
 sky130_fd_sc_hd__buf_2 output118 (.A(net1001),
    .X(out26));
 sky130_fd_sc_hd__buf_2 output119 (.A(net896),
    .X(out27));
 sky130_fd_sc_hd__clkbuf_1 output120 (.A(clknet_1_1__leaf_net897),
    .X(out28));
 sky130_fd_sc_hd__buf_2 output121 (.A(net1021),
    .X(out3));
 sky130_fd_sc_hd__clkbuf_1 output122 (.A(clknet_1_0__leaf_net899),
    .X(out30));
 sky130_fd_sc_hd__buf_2 output123 (.A(net900),
    .X(out31));
 sky130_fd_sc_hd__buf_2 output124 (.A(net901),
    .X(out32));
 sky130_fd_sc_hd__clkbuf_1 output125 (.A(clknet_1_1__leaf_net902),
    .X(out34));
 sky130_fd_sc_hd__buf_2 output126 (.A(net903),
    .X(out35));
 sky130_fd_sc_hd__buf_2 output127 (.A(net904),
    .X(out36));
 sky130_fd_sc_hd__buf_2 output128 (.A(net999),
    .X(out37));
 sky130_fd_sc_hd__buf_2 output129 (.A(net1023),
    .X(out38));
 sky130_fd_sc_hd__clkbuf_1 output130 (.A(clknet_1_1__leaf_net907),
    .X(out39));
 sky130_fd_sc_hd__clkbuf_1 output131 (.A(clknet_1_1__leaf_net908),
    .X(out4));
 sky130_fd_sc_hd__clkbuf_1 output132 (.A(clknet_1_1__leaf_net909),
    .X(out40));
 sky130_fd_sc_hd__buf_2 output133 (.A(net994),
    .X(out41));
 sky130_fd_sc_hd__clkbuf_1 output134 (.A(clknet_1_0__leaf_net911),
    .X(out42));
 sky130_fd_sc_hd__buf_2 output135 (.A(net912),
    .X(out45));
 sky130_fd_sc_hd__buf_2 output136 (.A(net913),
    .X(out46));
 sky130_fd_sc_hd__clkbuf_1 output137 (.A(clknet_1_1__leaf_net914),
    .X(out47));
 sky130_fd_sc_hd__buf_2 output138 (.A(net915),
    .X(out48));
 sky130_fd_sc_hd__buf_2 output139 (.A(net916),
    .X(out49));
 sky130_fd_sc_hd__clkbuf_1 output140 (.A(clknet_1_1__leaf_net917),
    .X(out5));
 sky130_fd_sc_hd__clkbuf_1 output141 (.A(clknet_1_0__leaf_net918),
    .X(out50));
 sky130_fd_sc_hd__clkbuf_1 output142 (.A(clknet_1_0__leaf_net919),
    .X(out51));
 sky130_fd_sc_hd__buf_2 output143 (.A(net920),
    .X(out52));
 sky130_fd_sc_hd__buf_2 output144 (.A(net971),
    .X(out53));
 sky130_fd_sc_hd__clkbuf_1 output145 (.A(clknet_1_0__leaf_net922),
    .X(out54));
 sky130_fd_sc_hd__buf_2 output146 (.A(net923),
    .X(out55));
 sky130_fd_sc_hd__clkbuf_1 output147 (.A(clknet_1_0__leaf_net924),
    .X(out56));
 sky130_fd_sc_hd__clkbuf_1 output148 (.A(clknet_1_1__leaf_net925),
    .X(out58));
 sky130_fd_sc_hd__buf_2 output149 (.A(net926),
    .X(out59));
 sky130_fd_sc_hd__clkbuf_1 output150 (.A(clknet_1_1__leaf_net927),
    .X(out60));
 sky130_fd_sc_hd__clkbuf_1 output151 (.A(clknet_1_1__leaf_net928),
    .X(out61));
 sky130_fd_sc_hd__buf_2 output152 (.A(net1042),
    .X(out62));
 sky130_fd_sc_hd__buf_2 output153 (.A(net930),
    .X(out63));
 sky130_fd_sc_hd__clkbuf_1 output154 (.A(clknet_1_1__leaf_net931),
    .X(out64));
 sky130_fd_sc_hd__buf_2 output155 (.A(net932),
    .X(out65));
 sky130_fd_sc_hd__clkbuf_1 output156 (.A(clknet_1_0__leaf_net933),
    .X(out67));
 sky130_fd_sc_hd__buf_2 output157 (.A(net934),
    .X(out68));
 sky130_fd_sc_hd__buf_2 output158 (.A(net935),
    .X(out7));
 sky130_fd_sc_hd__buf_2 output159 (.A(net936),
    .X(out70));
 sky130_fd_sc_hd__buf_2 output160 (.A(net937),
    .X(out71));
 sky130_fd_sc_hd__clkbuf_1 output161 (.A(clknet_1_0__leaf_net938),
    .X(out72));
 sky130_fd_sc_hd__buf_2 output162 (.A(net939),
    .X(out73));
 sky130_fd_sc_hd__buf_2 output163 (.A(net940),
    .X(out74));
 sky130_fd_sc_hd__buf_2 output164 (.A(net941),
    .X(out75));
 sky130_fd_sc_hd__clkbuf_1 output165 (.A(clknet_1_0__leaf_net942),
    .X(out76));
 sky130_fd_sc_hd__buf_2 output166 (.A(net943),
    .X(out78));
 sky130_fd_sc_hd__clkbuf_1 output167 (.A(clknet_1_0__leaf_net944),
    .X(out79));
 sky130_fd_sc_hd__clkbuf_1 output168 (.A(clknet_1_1__leaf_net945),
    .X(out8));
 sky130_fd_sc_hd__buf_2 output169 (.A(net946),
    .X(out80));
 sky130_fd_sc_hd__buf_2 output170 (.A(net947),
    .X(out81));
 sky130_fd_sc_hd__clkbuf_1 output171 (.A(clknet_1_0__leaf_net948),
    .X(out83));
 sky130_fd_sc_hd__buf_2 output172 (.A(net949),
    .X(out84));
 sky130_fd_sc_hd__buf_2 output173 (.A(net950),
    .X(out85));
 sky130_fd_sc_hd__buf_2 output174 (.A(net951),
    .X(out88));
 sky130_fd_sc_hd__clkbuf_1 output175 (.A(clknet_1_1__leaf_net952),
    .X(out89));
 sky130_fd_sc_hd__buf_2 output176 (.A(net953),
    .X(out90));
 sky130_fd_sc_hd__buf_2 output177 (.A(net954),
    .X(out91));
 sky130_fd_sc_hd__buf_2 output178 (.A(net955),
    .X(out93));
 sky130_fd_sc_hd__buf_2 output179 (.A(net956),
    .X(out94));
 sky130_fd_sc_hd__buf_2 output180 (.A(net957),
    .X(out95));
 sky130_fd_sc_hd__buf_2 output181 (.A(net958),
    .X(out96));
 sky130_fd_sc_hd__buf_2 output182 (.A(net959),
    .X(out98));
 sky130_fd_sc_hd__buf_2 output183 (.A(net960),
    .X(out99));
 sky130_fd_sc_hd__buf_2 fanout184 (.A(net260),
    .X(net961));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout185 (.A(net260),
    .X(net962));
 sky130_fd_sc_hd__clkbuf_2 fanout186 (.A(net248),
    .X(net963));
 sky130_fd_sc_hd__clkbuf_4 fanout187 (.A(net965),
    .X(net964));
 sky130_fd_sc_hd__buf_4 fanout188 (.A(net233),
    .X(net965));
 sky130_fd_sc_hd__buf_4 fanout189 (.A(net160),
    .X(net966));
 sky130_fd_sc_hd__clkbuf_4 fanout190 (.A(net880),
    .X(net967));
 sky130_fd_sc_hd__buf_2 fanout191 (.A(net73),
    .X(net968));
 sky130_fd_sc_hd__clkbuf_4 fanout192 (.A(net1051),
    .X(net969));
 sky130_fd_sc_hd__buf_8 fanout193 (.A(net236),
    .X(net970));
 sky130_fd_sc_hd__buf_4 fanout194 (.A(net921),
    .X(net971));
 sky130_fd_sc_hd__clkbuf_4 fanout195 (.A(net147),
    .X(net972));
 sky130_fd_sc_hd__buf_4 fanout196 (.A(net53),
    .X(net973));
 sky130_fd_sc_hd__buf_2 fanout197 (.A(net53),
    .X(net974));
 sky130_fd_sc_hd__buf_2 fanout198 (.A(net976),
    .X(net975));
 sky130_fd_sc_hd__buf_2 fanout199 (.A(net977),
    .X(net976));
 sky130_fd_sc_hd__buf_2 fanout200 (.A(net232),
    .X(net977));
 sky130_fd_sc_hd__buf_2 fanout201 (.A(net170),
    .X(net978));
 sky130_fd_sc_hd__buf_6 fanout202 (.A(net150),
    .X(net979));
 sky130_fd_sc_hd__buf_1 fanout203 (.A(net150),
    .X(net980));
 sky130_fd_sc_hd__buf_8 fanout204 (.A(net982),
    .X(net981));
 sky130_fd_sc_hd__buf_6 fanout205 (.A(net132),
    .X(net982));
 sky130_fd_sc_hd__buf_8 fanout206 (.A(net984),
    .X(net983));
 sky130_fd_sc_hd__buf_6 fanout207 (.A(net130),
    .X(net984));
 sky130_fd_sc_hd__clkbuf_4 fanout208 (.A(net986),
    .X(net985));
 sky130_fd_sc_hd__buf_4 fanout209 (.A(net48),
    .X(net986));
 sky130_fd_sc_hd__buf_2 fanout210 (.A(net149),
    .X(net987));
 sky130_fd_sc_hd__buf_6 fanout211 (.A(net127),
    .X(net988));
 sky130_fd_sc_hd__clkbuf_4 fanout212 (.A(net65),
    .X(net989));
 sky130_fd_sc_hd__clkbuf_4 fanout213 (.A(net991),
    .X(net990));
 sky130_fd_sc_hd__buf_2 fanout214 (.A(net42),
    .X(net991));
 sky130_fd_sc_hd__buf_12 fanout215 (.A(net994),
    .X(net992));
 sky130_fd_sc_hd__buf_2 fanout216 (.A(net994),
    .X(net993));
 sky130_fd_sc_hd__buf_12 fanout217 (.A(net910),
    .X(net994));
 sky130_fd_sc_hd__clkbuf_4 fanout218 (.A(net996),
    .X(net995));
 sky130_fd_sc_hd__buf_2 fanout219 (.A(net33),
    .X(net996));
 sky130_fd_sc_hd__buf_8 fanout220 (.A(net929),
    .X(net997));
 sky130_fd_sc_hd__clkbuf_2 fanout221 (.A(net929),
    .X(net998));
 sky130_fd_sc_hd__buf_2 fanout222 (.A(net905),
    .X(net999));
 sky130_fd_sc_hd__buf_2 fanout223 (.A(net259),
    .X(net1000));
 sky130_fd_sc_hd__clkbuf_4 fanout224 (.A(net895),
    .X(net1001));
 sky130_fd_sc_hd__clkbuf_4 fanout225 (.A(net460),
    .X(net1002));
 sky130_fd_sc_hd__buf_12 fanout226 (.A(net1004),
    .X(net1003));
 sky130_fd_sc_hd__buf_8 fanout227 (.A(net22),
    .X(net1004));
 sky130_fd_sc_hd__clkbuf_4 fanout228 (.A(net935),
    .X(net1005));
 sky130_fd_sc_hd__clkbuf_4 fanout229 (.A(net345),
    .X(net1006));
 sky130_fd_sc_hd__buf_8 fanout230 (.A(net1008),
    .X(net1007));
 sky130_fd_sc_hd__buf_8 fanout231 (.A(net20),
    .X(net1008));
 sky130_fd_sc_hd__clkbuf_4 fanout232 (.A(net754),
    .X(net1009));
 sky130_fd_sc_hd__buf_4 fanout233 (.A(net731),
    .X(net1010));
 sky130_fd_sc_hd__buf_2 max_cap234 (.A(net711),
    .X(net1011));
 sky130_fd_sc_hd__clkbuf_4 fanout235 (.A(net710),
    .X(net1012));
 sky130_fd_sc_hd__buf_4 fanout236 (.A(net698),
    .X(net1013));
 sky130_fd_sc_hd__clkbuf_4 fanout237 (.A(net691),
    .X(net1014));
 sky130_fd_sc_hd__clkbuf_4 fanout238 (.A(net1016),
    .X(net1015));
 sky130_fd_sc_hd__buf_2 fanout239 (.A(net689),
    .X(net1016));
 sky130_fd_sc_hd__clkbuf_4 fanout240 (.A(net1018),
    .X(net1017));
 sky130_fd_sc_hd__clkbuf_2 fanout241 (.A(net673),
    .X(net1018));
 sky130_fd_sc_hd__clkbuf_2 max_cap242 (.A(net672),
    .X(net1019));
 sky130_fd_sc_hd__clkbuf_4 fanout243 (.A(net670),
    .X(net1020));
 sky130_fd_sc_hd__buf_4 max_cap244 (.A(net898),
    .X(net1021));
 sky130_fd_sc_hd__buf_4 fanout245 (.A(net667),
    .X(net1022));
 sky130_fd_sc_hd__buf_4 fanout246 (.A(net906),
    .X(net1023));
 sky130_fd_sc_hd__buf_12 fanout247 (.A(net867),
    .X(net1024));
 sky130_fd_sc_hd__buf_4 fanout248 (.A(net785),
    .X(net1025));
 sky130_fd_sc_hd__clkbuf_4 fanout249 (.A(net785),
    .X(net1026));
 sky130_fd_sc_hd__buf_4 fanout250 (.A(net1028),
    .X(net1027));
 sky130_fd_sc_hd__buf_2 fanout251 (.A(net856),
    .X(net1028));
 sky130_fd_sc_hd__clkbuf_4 fanout252 (.A(net824),
    .X(net1029));
 sky130_fd_sc_hd__clkbuf_2 fanout253 (.A(net824),
    .X(net1030));
 sky130_fd_sc_hd__clkbuf_8 fanout254 (.A(net823),
    .X(net1031));
 sky130_fd_sc_hd__buf_4 fanout255 (.A(net815),
    .X(net1032));
 sky130_fd_sc_hd__buf_4 fanout256 (.A(net780),
    .X(net1033));
 sky130_fd_sc_hd__clkbuf_4 fanout257 (.A(net796),
    .X(net1034));
 sky130_fd_sc_hd__buf_6 fanout258 (.A(net1036),
    .X(net1035));
 sky130_fd_sc_hd__buf_2 fanout259 (.A(net789),
    .X(net1036));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net775 (.A(net775),
    .X(clknet_0_net775));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net775 (.A(clknet_0_net775),
    .X(clknet_1_0__leaf_net775));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net775 (.A(clknet_0_net775),
    .X(clknet_1_1__leaf_net775));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net883 (.A(net883),
    .X(clknet_0_net883));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net883 (.A(clknet_0_net883),
    .X(clknet_1_0__leaf_net883));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net883 (.A(clknet_0_net883),
    .X(clknet_1_1__leaf_net883));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net533 (.A(net533),
    .X(clknet_0_net533));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net533 (.A(clknet_0_net533),
    .X(clknet_1_0__leaf_net533));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net533 (.A(clknet_0_net533),
    .X(clknet_1_1__leaf_net533));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net945 (.A(net945),
    .X(clknet_0_net945));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net945 (.A(clknet_0_net945),
    .X(clknet_1_0__leaf_net945));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net945 (.A(clknet_0_net945),
    .X(clknet_1_1__leaf_net945));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net758 (.A(net758),
    .X(clknet_0_net758));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net758 (.A(clknet_0_net758),
    .X(clknet_1_0__leaf_net758));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net758 (.A(clknet_0_net758),
    .X(clknet_1_1__leaf_net758));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net489 (.A(net489),
    .X(clknet_0_net489));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net489 (.A(clknet_0_net489),
    .X(clknet_1_0__leaf_net489));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net489 (.A(clknet_0_net489),
    .X(clknet_1_1__leaf_net489));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net487 (.A(net487),
    .X(clknet_0_net487));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net487 (.A(clknet_0_net487),
    .X(clknet_1_0__leaf_net487));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net487 (.A(clknet_0_net487),
    .X(clknet_1_1__leaf_net487));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net757 (.A(net757),
    .X(clknet_0_net757));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net757 (.A(clknet_0_net757),
    .X(clknet_1_0__leaf_net757));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net757 (.A(clknet_0_net757),
    .X(clknet_1_1__leaf_net757));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net484 (.A(net484),
    .X(clknet_0_net484));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net484 (.A(clknet_0_net484),
    .X(clknet_1_0__leaf_net484));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net484 (.A(clknet_0_net484),
    .X(clknet_1_1__leaf_net484));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net504 (.A(net504),
    .X(clknet_0_net504));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net504 (.A(clknet_0_net504),
    .X(clknet_1_0__leaf_net504));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net504 (.A(clknet_0_net504),
    .X(clknet_1_1__leaf_net504));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net506 (.A(net506),
    .X(clknet_0_net506));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net506 (.A(clknet_0_net506),
    .X(clknet_1_0__leaf_net506));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net506 (.A(clknet_0_net506),
    .X(clknet_1_1__leaf_net506));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net511 (.A(net511),
    .X(clknet_0_net511));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net511 (.A(clknet_0_net511),
    .X(clknet_1_0__leaf_net511));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net511 (.A(clknet_0_net511),
    .X(clknet_1_1__leaf_net511));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net481 (.A(net481),
    .X(clknet_0_net481));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net481 (.A(clknet_0_net481),
    .X(clknet_1_0__leaf_net481));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net481 (.A(clknet_0_net481),
    .X(clknet_1_1__leaf_net481));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net502 (.A(net502),
    .X(clknet_0_net502));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net502 (.A(clknet_0_net502),
    .X(clknet_1_0__leaf_net502));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net502 (.A(clknet_0_net502),
    .X(clknet_1_1__leaf_net502));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net497 (.A(net497),
    .X(clknet_0_net497));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net497 (.A(clknet_0_net497),
    .X(clknet_1_0__leaf_net497));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net497 (.A(clknet_0_net497),
    .X(clknet_1_1__leaf_net497));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net756 (.A(net756),
    .X(clknet_0_net756));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net756 (.A(clknet_0_net756),
    .X(clknet_1_0__leaf_net756));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net756 (.A(clknet_0_net756),
    .X(clknet_1_1__leaf_net756));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net527 (.A(net527),
    .X(clknet_0_net527));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net527 (.A(clknet_0_net527),
    .X(clknet_1_0__leaf_net527));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net527 (.A(clknet_0_net527),
    .X(clknet_1_1__leaf_net527));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net740 (.A(net740),
    .X(clknet_0_net740));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net740 (.A(clknet_0_net740),
    .X(clknet_1_0__leaf_net740));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net740 (.A(clknet_0_net740),
    .X(clknet_1_1__leaf_net740));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net399 (.A(net399),
    .X(clknet_0_net399));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net399 (.A(clknet_0_net399),
    .X(clknet_1_0__leaf_net399));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net399 (.A(clknet_0_net399),
    .X(clknet_1_1__leaf_net399));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net899 (.A(net899),
    .X(clknet_0_net899));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net899 (.A(clknet_0_net899),
    .X(clknet_1_0__leaf_net899));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net899 (.A(clknet_0_net899),
    .X(clknet_1_1__leaf_net899));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net428 (.A(net428),
    .X(clknet_0_net428));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net428 (.A(clknet_0_net428),
    .X(clknet_1_0__leaf_net428));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net428 (.A(clknet_0_net428),
    .X(clknet_1_1__leaf_net428));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net420 (.A(net420),
    .X(clknet_0_net420));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net420 (.A(clknet_0_net420),
    .X(clknet_1_0__leaf_net420));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net420 (.A(clknet_0_net420),
    .X(clknet_1_1__leaf_net420));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net421 (.A(net421),
    .X(clknet_0_net421));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net421 (.A(clknet_0_net421),
    .X(clknet_1_0__leaf_net421));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net421 (.A(clknet_0_net421),
    .X(clknet_1_1__leaf_net421));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net400 (.A(net400),
    .X(clknet_0_net400));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net400 (.A(clknet_0_net400),
    .X(clknet_1_0__leaf_net400));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net400 (.A(clknet_0_net400),
    .X(clknet_1_1__leaf_net400));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net739 (.A(net739),
    .X(clknet_0_net739));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net739 (.A(clknet_0_net739),
    .X(clknet_1_0__leaf_net739));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net739 (.A(clknet_0_net739),
    .X(clknet_1_1__leaf_net739));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net405 (.A(net405),
    .X(clknet_0_net405));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net405 (.A(clknet_0_net405),
    .X(clknet_1_0__leaf_net405));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net405 (.A(clknet_0_net405),
    .X(clknet_1_1__leaf_net405));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net404 (.A(net404),
    .X(clknet_0_net404));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net404 (.A(clknet_0_net404),
    .X(clknet_1_0__leaf_net404));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net404 (.A(clknet_0_net404),
    .X(clknet_1_1__leaf_net404));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net884 (.A(net884),
    .X(clknet_0_net884));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net884 (.A(clknet_0_net884),
    .X(clknet_1_0__leaf_net884));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net884 (.A(clknet_0_net884),
    .X(clknet_1_1__leaf_net884));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net495 (.A(net495),
    .X(clknet_0_net495));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net495 (.A(clknet_0_net495),
    .X(clknet_1_0__leaf_net495));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net495 (.A(clknet_0_net495),
    .X(clknet_1_1__leaf_net495));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net494 (.A(net494),
    .X(clknet_0_net494));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net494 (.A(clknet_0_net494),
    .X(clknet_1_0__leaf_net494));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net494 (.A(clknet_0_net494),
    .X(clknet_1_1__leaf_net494));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net446 (.A(net446),
    .X(clknet_0_net446));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net446 (.A(clknet_0_net446),
    .X(clknet_1_0__leaf_net446));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net446 (.A(clknet_0_net446),
    .X(clknet_1_1__leaf_net446));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net908 (.A(net908),
    .X(clknet_0_net908));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net908 (.A(clknet_0_net908),
    .X(clknet_1_0__leaf_net908));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net908 (.A(clknet_0_net908),
    .X(clknet_1_1__leaf_net908));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net892 (.A(net892),
    .X(clknet_0_net892));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net892 (.A(clknet_0_net892),
    .X(clknet_1_0__leaf_net892));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net892 (.A(clknet_0_net892),
    .X(clknet_1_1__leaf_net892));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net402 (.A(net402),
    .X(clknet_0_net402));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net402 (.A(clknet_0_net402),
    .X(clknet_1_0__leaf_net402));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net402 (.A(clknet_0_net402),
    .X(clknet_1_1__leaf_net402));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net738 (.A(net738),
    .X(clknet_0_net738));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net738 (.A(clknet_0_net738),
    .X(clknet_1_0__leaf_net738));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net738 (.A(clknet_0_net738),
    .X(clknet_1_1__leaf_net738));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net721 (.A(net721),
    .X(clknet_0_net721));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net721 (.A(clknet_0_net721),
    .X(clknet_1_0__leaf_net721));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net721 (.A(clknet_0_net721),
    .X(clknet_1_1__leaf_net721));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net355 (.A(net355),
    .X(clknet_0_net355));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net355 (.A(clknet_0_net355),
    .X(clknet_1_0__leaf_net355));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net355 (.A(clknet_0_net355),
    .X(clknet_1_1__leaf_net355));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net361 (.A(net361),
    .X(clknet_0_net361));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net361 (.A(clknet_0_net361),
    .X(clknet_1_0__leaf_net361));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net361 (.A(clknet_0_net361),
    .X(clknet_1_1__leaf_net361));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net486 (.A(net486),
    .X(clknet_0_net486));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net486 (.A(clknet_0_net486),
    .X(clknet_1_0__leaf_net486));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net486 (.A(clknet_0_net486),
    .X(clknet_1_1__leaf_net486));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net394 (.A(net394),
    .X(clknet_0_net394));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net394 (.A(clknet_0_net394),
    .X(clknet_1_0__leaf_net394));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net394 (.A(clknet_0_net394),
    .X(clknet_1_1__leaf_net394));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net365 (.A(net365),
    .X(clknet_0_net365));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net365 (.A(clknet_0_net365),
    .X(clknet_1_0__leaf_net365));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net365 (.A(clknet_0_net365),
    .X(clknet_1_1__leaf_net365));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net645 (.A(net645),
    .X(clknet_0_net645));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net645 (.A(clknet_0_net645),
    .X(clknet_1_0__leaf_net645));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net645 (.A(clknet_0_net645),
    .X(clknet_1_1__leaf_net645));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net391 (.A(net391),
    .X(clknet_0_net391));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net391 (.A(clknet_0_net391),
    .X(clknet_1_0__leaf_net391));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net391 (.A(clknet_0_net391),
    .X(clknet_1_1__leaf_net391));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net376 (.A(net376),
    .X(clknet_0_net376));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net376 (.A(clknet_0_net376),
    .X(clknet_1_0__leaf_net376));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net376 (.A(clknet_0_net376),
    .X(clknet_1_1__leaf_net376));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net375 (.A(net375),
    .X(clknet_0_net375));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net375 (.A(clknet_0_net375),
    .X(clknet_1_0__leaf_net375));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net375 (.A(clknet_0_net375),
    .X(clknet_1_1__leaf_net375));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net473 (.A(net473),
    .X(clknet_0_net473));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net473 (.A(clknet_0_net473),
    .X(clknet_1_0__leaf_net473));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net473 (.A(clknet_0_net473),
    .X(clknet_1_1__leaf_net473));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net476 (.A(net476),
    .X(clknet_0_net476));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net476 (.A(clknet_0_net476),
    .X(clknet_1_0__leaf_net476));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net476 (.A(clknet_0_net476),
    .X(clknet_1_1__leaf_net476));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net612 (.A(net612),
    .X(clknet_0_net612));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net612 (.A(clknet_0_net612),
    .X(clknet_1_0__leaf_net612));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net612 (.A(clknet_0_net612),
    .X(clknet_1_1__leaf_net612));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net387 (.A(net387),
    .X(clknet_0_net387));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net387 (.A(clknet_0_net387),
    .X(clknet_1_0__leaf_net387));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net387 (.A(clknet_0_net387),
    .X(clknet_1_1__leaf_net387));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net389 (.A(net389),
    .X(clknet_0_net389));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net389 (.A(clknet_0_net389),
    .X(clknet_1_0__leaf_net389));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net389 (.A(clknet_0_net389),
    .X(clknet_1_1__leaf_net389));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net366 (.A(net366),
    .X(clknet_0_net366));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net366 (.A(clknet_0_net366),
    .X(clknet_1_0__leaf_net366));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net366 (.A(clknet_0_net366),
    .X(clknet_1_1__leaf_net366));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net388 (.A(net388),
    .X(clknet_0_net388));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net388 (.A(clknet_0_net388),
    .X(clknet_1_0__leaf_net388));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net388 (.A(clknet_0_net388),
    .X(clknet_1_1__leaf_net388));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net909 (.A(net909),
    .X(clknet_0_net909));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net909 (.A(clknet_0_net909),
    .X(clknet_1_0__leaf_net909));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net909 (.A(clknet_0_net909),
    .X(clknet_1_1__leaf_net909));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net379 (.A(net379),
    .X(clknet_0_net379));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net379 (.A(clknet_0_net379),
    .X(clknet_1_0__leaf_net379));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net379 (.A(clknet_0_net379),
    .X(clknet_1_1__leaf_net379));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net368 (.A(net368),
    .X(clknet_0_net368));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net368 (.A(clknet_0_net368),
    .X(clknet_1_0__leaf_net368));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net368 (.A(clknet_0_net368),
    .X(clknet_1_1__leaf_net368));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net369 (.A(net369),
    .X(clknet_0_net369));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net369 (.A(clknet_0_net369),
    .X(clknet_1_0__leaf_net369));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net369 (.A(clknet_0_net369),
    .X(clknet_1_1__leaf_net369));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net358 (.A(net358),
    .X(clknet_0_net358));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net358 (.A(clknet_0_net358),
    .X(clknet_1_0__leaf_net358));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net358 (.A(clknet_0_net358),
    .X(clknet_1_1__leaf_net358));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net450 (.A(net450),
    .X(clknet_0_net450));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net450 (.A(clknet_0_net450),
    .X(clknet_1_0__leaf_net450));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net450 (.A(clknet_0_net450),
    .X(clknet_1_1__leaf_net450));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net720 (.A(net720),
    .X(clknet_0_net720));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net720 (.A(clknet_0_net720),
    .X(clknet_1_0__leaf_net720));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net720 (.A(clknet_0_net720),
    .X(clknet_1_1__leaf_net720));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net354 (.A(net354),
    .X(clknet_0_net354));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net354 (.A(clknet_0_net354),
    .X(clknet_1_0__leaf_net354));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net354 (.A(clknet_0_net354),
    .X(clknet_1_1__leaf_net354));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net392 (.A(net392),
    .X(clknet_0_net392));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net392 (.A(clknet_0_net392),
    .X(clknet_1_0__leaf_net392));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net392 (.A(clknet_0_net392),
    .X(clknet_1_1__leaf_net392));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net386 (.A(net386),
    .X(clknet_0_net386));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net386 (.A(clknet_0_net386),
    .X(clknet_1_0__leaf_net386));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net386 (.A(clknet_0_net386),
    .X(clknet_1_1__leaf_net386));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net351 (.A(net351),
    .X(clknet_0_net351));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net351 (.A(clknet_0_net351),
    .X(clknet_1_0__leaf_net351));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net351 (.A(clknet_0_net351),
    .X(clknet_1_1__leaf_net351));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net719 (.A(net719),
    .X(clknet_0_net719));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net719 (.A(clknet_0_net719),
    .X(clknet_1_0__leaf_net719));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net719 (.A(clknet_0_net719),
    .X(clknet_1_1__leaf_net719));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net701 (.A(net701),
    .X(clknet_0_net701));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net701 (.A(clknet_0_net701),
    .X(clknet_1_0__leaf_net701));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net701 (.A(clknet_0_net701),
    .X(clknet_1_1__leaf_net701));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net385 (.A(net385),
    .X(clknet_0_net385));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net385 (.A(clknet_0_net385),
    .X(clknet_1_0__leaf_net385));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net385 (.A(clknet_0_net385),
    .X(clknet_1_1__leaf_net385));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net925 (.A(net925),
    .X(clknet_0_net925));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net925 (.A(clknet_0_net925),
    .X(clknet_1_0__leaf_net925));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net925 (.A(clknet_0_net925),
    .X(clknet_1_1__leaf_net925));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net301 (.A(net301),
    .X(clknet_0_net301));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net301 (.A(clknet_0_net301),
    .X(clknet_1_0__leaf_net301));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net301 (.A(clknet_0_net301),
    .X(clknet_1_1__leaf_net301));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net700 (.A(net700),
    .X(clknet_0_net700));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net700 (.A(clknet_0_net700),
    .X(clknet_1_0__leaf_net700));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net700 (.A(clknet_0_net700),
    .X(clknet_1_1__leaf_net700));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net275 (.A(net275),
    .X(clknet_0_net275));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net275 (.A(clknet_0_net275),
    .X(clknet_1_0__leaf_net275));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net275 (.A(clknet_0_net275),
    .X(clknet_1_1__leaf_net275));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net271 (.A(net271),
    .X(clknet_0_net271));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net271 (.A(clknet_0_net271),
    .X(clknet_1_0__leaf_net271));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net271 (.A(clknet_0_net271),
    .X(clknet_1_1__leaf_net271));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net305 (.A(net305),
    .X(clknet_0_net305));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net305 (.A(clknet_0_net305),
    .X(clknet_1_0__leaf_net305));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net305 (.A(clknet_0_net305),
    .X(clknet_1_1__leaf_net305));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net299 (.A(net299),
    .X(clknet_0_net299));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net299 (.A(clknet_0_net299),
    .X(clknet_1_0__leaf_net299));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net299 (.A(clknet_0_net299),
    .X(clknet_1_1__leaf_net299));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net917 (.A(net917),
    .X(clknet_0_net917));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net917 (.A(clknet_0_net917),
    .X(clknet_1_0__leaf_net917));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net917 (.A(clknet_0_net917),
    .X(clknet_1_1__leaf_net917));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net283 (.A(net283),
    .X(clknet_0_net283));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net283 (.A(clknet_0_net283),
    .X(clknet_1_0__leaf_net283));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net283 (.A(clknet_0_net283),
    .X(clknet_1_1__leaf_net283));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net277 (.A(net277),
    .X(clknet_0_net277));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net277 (.A(clknet_0_net277),
    .X(clknet_1_0__leaf_net277));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net277 (.A(clknet_0_net277),
    .X(clknet_1_1__leaf_net277));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net699 (.A(net699),
    .X(clknet_0_net699));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net699 (.A(clknet_0_net699),
    .X(clknet_1_0__leaf_net699));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net699 (.A(clknet_0_net699),
    .X(clknet_1_1__leaf_net699));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net269 (.A(net269),
    .X(clknet_0_net269));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net269 (.A(clknet_0_net269),
    .X(clknet_1_0__leaf_net269));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net269 (.A(clknet_0_net269),
    .X(clknet_1_1__leaf_net269));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net933 (.A(net933),
    .X(clknet_0_net933));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net933 (.A(clknet_0_net933),
    .X(clknet_1_0__leaf_net933));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net933 (.A(clknet_0_net933),
    .X(clknet_1_1__leaf_net933));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net288 (.A(net288),
    .X(clknet_0_net288));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net288 (.A(clknet_0_net288),
    .X(clknet_1_0__leaf_net288));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net288 (.A(clknet_0_net288),
    .X(clknet_1_1__leaf_net288));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net291 (.A(net291),
    .X(clknet_0_net291));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net291 (.A(clknet_0_net291),
    .X(clknet_1_0__leaf_net291));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net291 (.A(clknet_0_net291),
    .X(clknet_1_1__leaf_net291));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net220 (.A(net220),
    .X(clknet_0_net220));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net220 (.A(clknet_0_net220),
    .X(clknet_1_0__leaf_net220));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net220 (.A(clknet_0_net220),
    .X(clknet_1_1__leaf_net220));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net942 (.A(net942),
    .X(clknet_0_net942));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net942 (.A(clknet_0_net942),
    .X(clknet_1_0__leaf_net942));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net942 (.A(clknet_0_net942),
    .X(clknet_1_1__leaf_net942));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net226 (.A(net226),
    .X(clknet_0_net226));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net226 (.A(clknet_0_net226),
    .X(clknet_1_0__leaf_net226));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net226 (.A(clknet_0_net226),
    .X(clknet_1_1__leaf_net226));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net222 (.A(net222),
    .X(clknet_0_net222));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net222 (.A(clknet_0_net222),
    .X(clknet_1_0__leaf_net222));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net222 (.A(clknet_0_net222),
    .X(clknet_1_1__leaf_net222));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net208 (.A(net208),
    .X(clknet_0_net208));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net208 (.A(clknet_0_net208),
    .X(clknet_1_0__leaf_net208));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net208 (.A(clknet_0_net208),
    .X(clknet_1_1__leaf_net208));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net914 (.A(net914),
    .X(clknet_0_net914));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net914 (.A(clknet_0_net914),
    .X(clknet_1_0__leaf_net914));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net914 (.A(clknet_0_net914),
    .X(clknet_1_1__leaf_net914));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net328 (.A(net328),
    .X(clknet_0_net328));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net328 (.A(clknet_0_net328),
    .X(clknet_1_0__leaf_net328));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net328 (.A(clknet_0_net328),
    .X(clknet_1_1__leaf_net328));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net320 (.A(net320),
    .X(clknet_0_net320));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net320 (.A(clknet_0_net320),
    .X(clknet_1_0__leaf_net320));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net320 (.A(clknet_0_net320),
    .X(clknet_1_1__leaf_net320));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net216 (.A(net216),
    .X(clknet_0_net216));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net216 (.A(clknet_0_net216),
    .X(clknet_1_0__leaf_net216));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net216 (.A(clknet_0_net216),
    .X(clknet_1_1__leaf_net216));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net214 (.A(net214),
    .X(clknet_0_net214));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net214 (.A(clknet_0_net214),
    .X(clknet_1_0__leaf_net214));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net214 (.A(clknet_0_net214),
    .X(clknet_1_1__leaf_net214));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net922 (.A(net922),
    .X(clknet_0_net922));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net922 (.A(clknet_0_net922),
    .X(clknet_1_0__leaf_net922));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net922 (.A(clknet_0_net922),
    .X(clknet_1_1__leaf_net922));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net330 (.A(net330),
    .X(clknet_0_net330));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net330 (.A(clknet_0_net330),
    .X(clknet_1_0__leaf_net330));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net330 (.A(clknet_0_net330),
    .X(clknet_1_1__leaf_net330));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net331 (.A(net331),
    .X(clknet_0_net331));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net331 (.A(clknet_0_net331),
    .X(clknet_1_0__leaf_net331));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net331 (.A(clknet_0_net331),
    .X(clknet_1_1__leaf_net331));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net918 (.A(net918),
    .X(clknet_0_net918));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net918 (.A(clknet_0_net918),
    .X(clknet_1_0__leaf_net918));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net918 (.A(clknet_0_net918),
    .X(clknet_1_1__leaf_net918));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net902 (.A(net902),
    .X(clknet_0_net902));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net902 (.A(clknet_0_net902),
    .X(clknet_1_0__leaf_net902));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net902 (.A(clknet_0_net902),
    .X(clknet_1_1__leaf_net902));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net680 (.A(net680),
    .X(clknet_0_net680));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net680 (.A(clknet_0_net680),
    .X(clknet_1_0__leaf_net680));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net680 (.A(clknet_0_net680),
    .X(clknet_1_1__leaf_net680));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net907 (.A(net907),
    .X(clknet_0_net907));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net907 (.A(clknet_0_net907),
    .X(clknet_1_0__leaf_net907));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net907 (.A(clknet_0_net907),
    .X(clknet_1_1__leaf_net907));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net911 (.A(net911),
    .X(clknet_0_net911));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net911 (.A(clknet_0_net911),
    .X(clknet_1_0__leaf_net911));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net911 (.A(clknet_0_net911),
    .X(clknet_1_1__leaf_net911));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net938 (.A(net938),
    .X(clknet_0_net938));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net938 (.A(clknet_0_net938),
    .X(clknet_1_0__leaf_net938));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net938 (.A(clknet_0_net938),
    .X(clknet_1_1__leaf_net938));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net664 (.A(net664),
    .X(clknet_0_net664));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net664 (.A(clknet_0_net664),
    .X(clknet_1_0__leaf_net664));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net664 (.A(clknet_0_net664),
    .X(clknet_1_1__leaf_net664));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net105 (.A(net105),
    .X(clknet_0_net105));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net105 (.A(clknet_0_net105),
    .X(clknet_1_0__leaf_net105));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net105 (.A(clknet_0_net105),
    .X(clknet_1_1__leaf_net105));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net325 (.A(net325),
    .X(clknet_0_net325));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net325 (.A(clknet_0_net325),
    .X(clknet_1_0__leaf_net325));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net325 (.A(clknet_0_net325),
    .X(clknet_1_1__leaf_net325));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net218 (.A(net218),
    .X(clknet_0_net218));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net218 (.A(clknet_0_net218),
    .X(clknet_1_0__leaf_net218));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net218 (.A(clknet_0_net218),
    .X(clknet_1_1__leaf_net218));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net114 (.A(net114),
    .X(clknet_0_net114));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net114 (.A(clknet_0_net114),
    .X(clknet_1_0__leaf_net114));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net114 (.A(clknet_0_net114),
    .X(clknet_1_1__leaf_net114));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net111 (.A(net111),
    .X(clknet_0_net111));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net111 (.A(clknet_0_net111),
    .X(clknet_1_0__leaf_net111));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net111 (.A(clknet_0_net111),
    .X(clknet_1_1__leaf_net111));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net948 (.A(net948),
    .X(clknet_0_net948));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net948 (.A(clknet_0_net948),
    .X(clknet_1_0__leaf_net948));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net948 (.A(clknet_0_net948),
    .X(clknet_1_1__leaf_net948));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net952 (.A(net952),
    .X(clknet_0_net952));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net952 (.A(clknet_0_net952),
    .X(clknet_1_0__leaf_net952));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net952 (.A(clknet_0_net952),
    .X(clknet_1_1__leaf_net952));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net928 (.A(net928),
    .X(clknet_0_net928));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net928 (.A(clknet_0_net928),
    .X(clknet_1_0__leaf_net928));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net928 (.A(clknet_0_net928),
    .X(clknet_1_1__leaf_net928));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net927 (.A(net927),
    .X(clknet_0_net927));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net927 (.A(clknet_0_net927),
    .X(clknet_1_0__leaf_net927));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net927 (.A(clknet_0_net927),
    .X(clknet_1_1__leaf_net927));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net897 (.A(net897),
    .X(clknet_0_net897));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net897 (.A(clknet_0_net897),
    .X(clknet_1_0__leaf_net897));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net897 (.A(clknet_0_net897),
    .X(clknet_1_1__leaf_net897));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net110 (.A(net110),
    .X(clknet_0_net110));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net110 (.A(clknet_0_net110),
    .X(clknet_1_0__leaf_net110));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net110 (.A(clknet_0_net110),
    .X(clknet_1_1__leaf_net110));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net96 (.A(net96),
    .X(clknet_0_net96));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net96 (.A(clknet_0_net96),
    .X(clknet_1_0__leaf_net96));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net96 (.A(clknet_0_net96),
    .X(clknet_1_1__leaf_net96));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net315 (.A(net315),
    .X(clknet_0_net315));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net315 (.A(clknet_0_net315),
    .X(clknet_1_0__leaf_net315));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net315 (.A(clknet_0_net315),
    .X(clknet_1_1__leaf_net315));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net893 (.A(net893),
    .X(clknet_0_net893));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net893 (.A(clknet_0_net893),
    .X(clknet_1_0__leaf_net893));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net893 (.A(clknet_0_net893),
    .X(clknet_1_1__leaf_net893));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net412 (.A(net412),
    .X(clknet_0_net412));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net412 (.A(clknet_0_net412),
    .X(clknet_1_0__leaf_net412));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net412 (.A(clknet_0_net412),
    .X(clknet_1_1__leaf_net412));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net193 (.A(net193),
    .X(clknet_0_net193));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net193 (.A(clknet_0_net193),
    .X(clknet_1_0__leaf_net193));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net193 (.A(clknet_0_net193),
    .X(clknet_1_1__leaf_net193));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net99 (.A(net99),
    .X(clknet_0_net99));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net99 (.A(clknet_0_net99),
    .X(clknet_1_0__leaf_net99));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net99 (.A(clknet_0_net99),
    .X(clknet_1_1__leaf_net99));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net614 (.A(net614),
    .X(clknet_0_net614));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net614 (.A(clknet_0_net614),
    .X(clknet_1_0__leaf_net614));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net614 (.A(clknet_0_net614),
    .X(clknet_1_1__leaf_net614));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net190 (.A(net190),
    .X(clknet_0_net190));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net190 (.A(clknet_0_net190),
    .X(clknet_1_0__leaf_net190));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net190 (.A(clknet_0_net190),
    .X(clknet_1_1__leaf_net190));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net196 (.A(net196),
    .X(clknet_0_net196));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net196 (.A(clknet_0_net196),
    .X(clknet_1_0__leaf_net196));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net196 (.A(clknet_0_net196),
    .X(clknet_1_1__leaf_net196));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net919 (.A(net919),
    .X(clknet_0_net919));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net919 (.A(clknet_0_net919),
    .X(clknet_1_0__leaf_net919));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net919 (.A(clknet_0_net919),
    .X(clknet_1_1__leaf_net919));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net944 (.A(net944),
    .X(clknet_0_net944));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net944 (.A(clknet_0_net944),
    .X(clknet_1_0__leaf_net944));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net944 (.A(clknet_0_net944),
    .X(clknet_1_1__leaf_net944));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net199 (.A(net199),
    .X(clknet_0_net199));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net199 (.A(clknet_0_net199),
    .X(clknet_1_0__leaf_net199));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net199 (.A(clknet_0_net199),
    .X(clknet_1_1__leaf_net199));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net200 (.A(net200),
    .X(clknet_0_net200));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net200 (.A(clknet_0_net200),
    .X(clknet_1_0__leaf_net200));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net200 (.A(clknet_0_net200),
    .X(clknet_1_1__leaf_net200));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net100 (.A(net100),
    .X(clknet_0_net100));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net100 (.A(clknet_0_net100),
    .X(clknet_1_0__leaf_net100));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net100 (.A(clknet_0_net100),
    .X(clknet_1_1__leaf_net100));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net663 (.A(net663),
    .X(clknet_0_net663));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net663 (.A(clknet_0_net663),
    .X(clknet_1_0__leaf_net663));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net663 (.A(clknet_0_net663),
    .X(clknet_1_1__leaf_net663));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net931 (.A(net931),
    .X(clknet_0_net931));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net931 (.A(clknet_0_net931),
    .X(clknet_1_0__leaf_net931));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net931 (.A(clknet_0_net931),
    .X(clknet_1_1__leaf_net931));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net924 (.A(net924),
    .X(clknet_0_net924));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net924 (.A(clknet_0_net924),
    .X(clknet_1_0__leaf_net924));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net924 (.A(clknet_0_net924),
    .X(clknet_1_1__leaf_net924));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net646 (.A(net646),
    .X(clknet_0_net646));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net646 (.A(clknet_0_net646),
    .X(clknet_1_0__leaf_net646));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net646 (.A(clknet_0_net646),
    .X(clknet_1_1__leaf_net646));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net468 (.A(net468),
    .X(clknet_0_net468));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net468 (.A(clknet_0_net468),
    .X(clknet_1_0__leaf_net468));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net468 (.A(clknet_0_net468),
    .X(clknet_1_1__leaf_net468));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net474 (.A(net474),
    .X(clknet_0_net474));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net474 (.A(clknet_0_net474),
    .X(clknet_1_0__leaf_net474));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net474 (.A(clknet_0_net474),
    .X(clknet_1_1__leaf_net474));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net467 (.A(net467),
    .X(clknet_0_net467));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net467 (.A(clknet_0_net467),
    .X(clknet_1_0__leaf_net467));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net467 (.A(clknet_0_net467),
    .X(clknet_1_1__leaf_net467));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net462 (.A(net462),
    .X(clknet_0_net462));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net462 (.A(clknet_0_net462),
    .X(clknet_1_0__leaf_net462));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net462 (.A(clknet_0_net462),
    .X(clknet_1_1__leaf_net462));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net613 (.A(net613),
    .X(clknet_0_net613));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net613 (.A(clknet_0_net613),
    .X(clknet_1_0__leaf_net613));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net613 (.A(clknet_0_net613),
    .X(clknet_1_1__leaf_net613));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net189 (.A(net189),
    .X(clknet_0_net189));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net189 (.A(clknet_0_net189),
    .X(clknet_1_0__leaf_net189));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net189 (.A(clknet_0_net189),
    .X(clknet_1_1__leaf_net189));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net169 (.A(net169),
    .X(clknet_0_net169));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net169 (.A(clknet_0_net169),
    .X(clknet_1_0__leaf_net169));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net169 (.A(clknet_0_net169),
    .X(clknet_1_1__leaf_net169));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net198 (.A(net198),
    .X(clknet_0_net198));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net198 (.A(clknet_0_net198),
    .X(clknet_1_0__leaf_net198));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net198 (.A(clknet_0_net198),
    .X(clknet_1_1__leaf_net198));
 sky130_fd_sc_hd__dlygate4sd3_1 rebuffer1 (.A(net1078),
    .X(net1037));
 sky130_fd_sc_hd__a2111o_1 clone2 (.A1(net21),
    .A2(net1025),
    .B1(net1063),
    .C1(net1003),
    .D1(net1039),
    .X(net1038));
 sky130_fd_sc_hd__a2111o_1 clone3 (.A1(net801),
    .A2(net790),
    .B1(net784),
    .C1(net786),
    .D1(net1024),
    .X(net1039));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer4 (.A(net921),
    .X(net1040));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer5 (.A(net1040),
    .X(net1041));
 sky130_fd_sc_hd__clkbuf_1 clone6 (.A(net1043),
    .X(net1042));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer7 (.A(net929),
    .X(net1043));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer8 (.A(net1053),
    .X(net1044));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer9 (.A(net1044),
    .X(net1045));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer10 (.A(net1044),
    .X(net1046));
 sky130_fd_sc_hd__clkbuf_1 clone11 (.A(net127),
    .X(net1047));
 sky130_fd_sc_hd__clkbuf_1 clone12 (.A(net1049),
    .X(net1048));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer13 (.A(net132),
    .X(net1049));
 sky130_fd_sc_hd__clkbuf_1 clone14 (.A(net22),
    .X(net1050));
 sky130_fd_sc_hd__clkbuf_1 clone15 (.A(net236),
    .X(net1051));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer16 (.A(net133),
    .X(net1052));
 sky130_fd_sc_hd__clkbuf_1 clone17 (.A(net867),
    .X(net1053));
 sky130_fd_sc_hd__clkbuf_4 clone18 (.A(net1004),
    .X(net1054));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer19 (.A(net1004),
    .X(net1055));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer20 (.A(net1055),
    .X(net1056));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer21 (.A(net981),
    .X(net1057));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer22 (.A(net1057),
    .X(net1058));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer23 (.A(net981),
    .X(net1059));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer24 (.A(net1059),
    .X(net1060));
 sky130_fd_sc_hd__clkbuf_1 clone25 (.A(net984),
    .X(net1061));
 sky130_fd_sc_hd__clkbuf_1 clone26 (.A(net1063),
    .X(net1062));
 sky130_fd_sc_hd__clkbuf_1 clone27 (.A(net20),
    .X(net1063));
 sky130_fd_sc_hd__clkbuf_1 clone28 (.A(net994),
    .X(net1064));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer29 (.A(net981),
    .X(net1065));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(net657),
    .X(net1066));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(net724),
    .X(net1067));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(net662),
    .X(net1068));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(net951),
    .X(net1069));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(net661),
    .X(net1070));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(net639),
    .X(net1071));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(net145),
    .X(net1072));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(net660),
    .X(net1073));
 sky130_fd_sc_hd__clkbuf_1 fanout1 (.A(net1025),
    .X(net1074));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_A (.DIODE(clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(in0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(in1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(in10));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(in11));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(in12));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(in13));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(in14));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(in15));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(in16));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(in17));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(in18));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(in19));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(in2));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(in20));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(in21));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(in22));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(in23));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(in24));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(in25));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(in26));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(in27));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_A (.DIODE(in28));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_A (.DIODE(in29));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_A (.DIODE(in3));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_A (.DIODE(in30));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_A (.DIODE(in31));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_A (.DIODE(in32));
 sky130_fd_sc_hd__diode_2 ANTENNA_input28_A (.DIODE(in33));
 sky130_fd_sc_hd__diode_2 ANTENNA_input29_A (.DIODE(in34));
 sky130_fd_sc_hd__diode_2 ANTENNA_input30_A (.DIODE(in35));
 sky130_fd_sc_hd__diode_2 ANTENNA_input31_A (.DIODE(in36));
 sky130_fd_sc_hd__diode_2 ANTENNA_input32_A (.DIODE(in37));
 sky130_fd_sc_hd__diode_2 ANTENNA_input33_A (.DIODE(in38));
 sky130_fd_sc_hd__diode_2 ANTENNA_input34_A (.DIODE(in39));
 sky130_fd_sc_hd__diode_2 ANTENNA_input35_A (.DIODE(in4));
 sky130_fd_sc_hd__diode_2 ANTENNA_input36_A (.DIODE(in40));
 sky130_fd_sc_hd__diode_2 ANTENNA_input37_A (.DIODE(in41));
 sky130_fd_sc_hd__diode_2 ANTENNA_input38_A (.DIODE(in42));
 sky130_fd_sc_hd__diode_2 ANTENNA_input39_A (.DIODE(in43));
 sky130_fd_sc_hd__diode_2 ANTENNA_input40_A (.DIODE(in44));
 sky130_fd_sc_hd__diode_2 ANTENNA_input41_A (.DIODE(in45));
 sky130_fd_sc_hd__diode_2 ANTENNA_input42_A (.DIODE(in46));
 sky130_fd_sc_hd__diode_2 ANTENNA_input43_A (.DIODE(in47));
 sky130_fd_sc_hd__diode_2 ANTENNA_input44_A (.DIODE(in48));
 sky130_fd_sc_hd__diode_2 ANTENNA_input45_A (.DIODE(in49));
 sky130_fd_sc_hd__diode_2 ANTENNA_input46_A (.DIODE(in5));
 sky130_fd_sc_hd__diode_2 ANTENNA_input47_A (.DIODE(in50));
 sky130_fd_sc_hd__diode_2 ANTENNA_input48_A (.DIODE(in51));
 sky130_fd_sc_hd__diode_2 ANTENNA_input49_A (.DIODE(in52));
 sky130_fd_sc_hd__diode_2 ANTENNA_input50_A (.DIODE(in53));
 sky130_fd_sc_hd__diode_2 ANTENNA_input51_A (.DIODE(in54));
 sky130_fd_sc_hd__diode_2 ANTENNA_input52_A (.DIODE(in55));
 sky130_fd_sc_hd__diode_2 ANTENNA_input53_A (.DIODE(in56));
 sky130_fd_sc_hd__diode_2 ANTENNA_input54_A (.DIODE(in57));
 sky130_fd_sc_hd__diode_2 ANTENNA_input55_A (.DIODE(in58));
 sky130_fd_sc_hd__diode_2 ANTENNA_input56_A (.DIODE(in59));
 sky130_fd_sc_hd__diode_2 ANTENNA_input57_A (.DIODE(in6));
 sky130_fd_sc_hd__diode_2 ANTENNA_input58_A (.DIODE(in60));
 sky130_fd_sc_hd__diode_2 ANTENNA_input59_A (.DIODE(in61));
 sky130_fd_sc_hd__diode_2 ANTENNA_input60_A (.DIODE(in62));
 sky130_fd_sc_hd__diode_2 ANTENNA_input61_A (.DIODE(in63));
 sky130_fd_sc_hd__diode_2 ANTENNA_input62_A (.DIODE(in64));
 sky130_fd_sc_hd__diode_2 ANTENNA_input63_A (.DIODE(in65));
 sky130_fd_sc_hd__diode_2 ANTENNA_input64_A (.DIODE(in66));
 sky130_fd_sc_hd__diode_2 ANTENNA_input65_A (.DIODE(in67));
 sky130_fd_sc_hd__diode_2 ANTENNA_input66_A (.DIODE(in68));
 sky130_fd_sc_hd__diode_2 ANTENNA_input67_A (.DIODE(in69));
 sky130_fd_sc_hd__diode_2 ANTENNA_input68_A (.DIODE(in7));
 sky130_fd_sc_hd__diode_2 ANTENNA_input69_A (.DIODE(in70));
 sky130_fd_sc_hd__diode_2 ANTENNA_input70_A (.DIODE(in71));
 sky130_fd_sc_hd__diode_2 ANTENNA_input71_A (.DIODE(in72));
 sky130_fd_sc_hd__diode_2 ANTENNA_input72_A (.DIODE(in73));
 sky130_fd_sc_hd__diode_2 ANTENNA_input73_A (.DIODE(in74));
 sky130_fd_sc_hd__diode_2 ANTENNA_input74_A (.DIODE(in75));
 sky130_fd_sc_hd__diode_2 ANTENNA_input75_A (.DIODE(in76));
 sky130_fd_sc_hd__diode_2 ANTENNA_input76_A (.DIODE(in77));
 sky130_fd_sc_hd__diode_2 ANTENNA_input77_A (.DIODE(in78));
 sky130_fd_sc_hd__diode_2 ANTENNA_input78_A (.DIODE(in79));
 sky130_fd_sc_hd__diode_2 ANTENNA_input79_A (.DIODE(in8));
 sky130_fd_sc_hd__diode_2 ANTENNA_input80_A (.DIODE(in80));
 sky130_fd_sc_hd__diode_2 ANTENNA_input81_A (.DIODE(in81));
 sky130_fd_sc_hd__diode_2 ANTENNA_input82_A (.DIODE(in82));
 sky130_fd_sc_hd__diode_2 ANTENNA_input83_A (.DIODE(in83));
 sky130_fd_sc_hd__diode_2 ANTENNA_input84_A (.DIODE(in84));
 sky130_fd_sc_hd__diode_2 ANTENNA_input85_A (.DIODE(in85));
 sky130_fd_sc_hd__diode_2 ANTENNA_input86_A (.DIODE(in86));
 sky130_fd_sc_hd__diode_2 ANTENNA_input87_A (.DIODE(in87));
 sky130_fd_sc_hd__diode_2 ANTENNA_input88_A (.DIODE(in88));
 sky130_fd_sc_hd__diode_2 ANTENNA_input89_A (.DIODE(in89));
 sky130_fd_sc_hd__diode_2 ANTENNA_input90_A (.DIODE(in9));
 sky130_fd_sc_hd__diode_2 ANTENNA_input91_A (.DIODE(in90));
 sky130_fd_sc_hd__diode_2 ANTENNA_input92_A (.DIODE(in91));
 sky130_fd_sc_hd__diode_2 ANTENNA_input93_A (.DIODE(in92));
 sky130_fd_sc_hd__diode_2 ANTENNA_input94_A (.DIODE(in93));
 sky130_fd_sc_hd__diode_2 ANTENNA_input95_A (.DIODE(in94));
 sky130_fd_sc_hd__diode_2 ANTENNA_input96_A (.DIODE(in95));
 sky130_fd_sc_hd__diode_2 ANTENNA_input97_A (.DIODE(in96));
 sky130_fd_sc_hd__diode_2 ANTENNA_input98_A (.DIODE(in97));
 sky130_fd_sc_hd__diode_2 ANTENNA_input99_A (.DIODE(in98));
 sky130_fd_sc_hd__diode_2 ANTENNA_input100_A (.DIODE(in99));
 sky130_fd_sc_hd__diode_2 ANTENNA_c127_S0 (.DIODE(net0));
 sky130_fd_sc_hd__diode_2 ANTENNA_c113_A1 (.DIODE(net0));
 sky130_fd_sc_hd__diode_2 ANTENNA_c110_B1 (.DIODE(net0));
 sky130_fd_sc_hd__diode_2 ANTENNA_c106_S1 (.DIODE(net0));
 sky130_fd_sc_hd__diode_2 ANTENNA_c104_S1 (.DIODE(net0));
 sky130_fd_sc_hd__diode_2 ANTENNA_c103_S0 (.DIODE(net0));
 sky130_fd_sc_hd__diode_2 ANTENNA_c102_A3 (.DIODE(net0));
 sky130_fd_sc_hd__diode_2 ANTENNA_c100_X (.DIODE(net0));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net100_A (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c218_X (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_A0 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_A0 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_A3 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_A0 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c366_S1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c237_Q (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_A0 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_c297_A1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_S0 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_A2 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_A3 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_A3 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_c275_A1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_c271_B1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_c270_C1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_X (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout207_A (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_A3 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_A0 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_c269_X (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_A0 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_S0 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_A2 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_c279_S1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_c277_Q_N (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_A1 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_A0 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_A0 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_A1 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_A0 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_c277_Q (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_c671_A1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_c666_SCD (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_c665_RESET_B (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_c662_A1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_c531_A2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_c529_D (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_c528_SCD (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_c404_A1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_A2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_A1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_c279_X (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout195_A (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_A2 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_X (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_c672_A0 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_c662_B1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_c529_SCD (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_c413_A1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_B1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_X (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout203_A (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout202_A (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_X (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_A0 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_A0 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_B1 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_X (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout189_A (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA_c693_A2 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_X (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_A1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_A0 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_B1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c428_A1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c311_A1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_A0 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_Q (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout201_A (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_A1 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_A1 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_A2 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_A1 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_X (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA_c582_A1 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_A2 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_A1 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_A1 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_A1 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_A0 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_A0 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_X (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_A0 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_A3 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_A1 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_A1 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_A2 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_A1 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_A2 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_X (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone2_A1 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_c138_C1 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_c668_C1 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_c665_D (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_c661_A2 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_c265_B1 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_S0 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_c140_A1 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_c136_A1 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_c134_X (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone14_A (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout227_A (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_X (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone15_A (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout193_A (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c400_X (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_A0 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_A2 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_A1 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_A2 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_C1 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_A2 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_X (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge866_D (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA_c404_X (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_A0 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA_c565_A1 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_D (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_X (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout223_A (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA_c693_A0 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_A2 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_X (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_D1 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_c534_A0 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_c410_A3 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_c404_A2 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_c264_A2 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_S1 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_A1 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_S0 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_A2 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_A0 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_c143_X (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_c127_A0 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c120_A3 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c119_D1 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c110_C1 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c109_S0 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c108_A3 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c106_A1 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c105_X (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge843_SCE (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_X (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_A2 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c184_A1 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c180_A1 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_D1 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_A2 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_A0 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_S0 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_A2 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_A2 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_X (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout229_A (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA_c693_A1 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA_c660_A1 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA_c546_A2 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA_c533_X (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer1_A (.DIODE(net1078));
 sky130_fd_sc_hd__diode_2 ANTENNA_c408_A0 (.DIODE(net1075));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_S0 (.DIODE(net1075));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_A2 (.DIODE(net1075));
 sky130_fd_sc_hd__diode_2 ANTENNA_c267_C1 (.DIODE(net1075));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_A1 (.DIODE(net1075));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_A3 (.DIODE(net1075));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_A3 (.DIODE(net1075));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_X (.DIODE(net1075));
 sky130_fd_sc_hd__diode_2 ANTENNA_c538_A1 (.DIODE(net1077));
 sky130_fd_sc_hd__diode_2 ANTENNA_c530_D (.DIODE(net1077));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_C1 (.DIODE(net1076));
 sky130_fd_sc_hd__diode_2 ANTENNA_c264_B1 (.DIODE(net1077));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_A2 (.DIODE(net1077));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_A0 (.DIODE(net1077));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_X (.DIODE(net1077));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_A0 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_A1 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_c263_A2 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_c108_A1 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_c107_S0 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_c106_X (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_A0 (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_A0 (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_A0 (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA_c611_A0 (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA_c610_A0 (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_A2 (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_A2 (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_X (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_A1 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_A1 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_A0 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA_c676_S0 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA_c673_A2 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA_c672_S0 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA_c663_B1 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA_c661_X (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA_c678_A (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_A2 (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_A2 (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA_c680_A1 (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA_c676_A2 (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA_c670_B1 (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA_c666_Q_N (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A1 (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_A1 (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_A2 (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA_c674_A2 (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA_c671_A2 (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA_c668_A1 (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA_c667_RESET_B (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA_c666_Q (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_A0 (.DIODE(net457));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_A2 (.DIODE(net457));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_A0 (.DIODE(net457));
 sky130_fd_sc_hd__diode_2 ANTENNA_c691_A0 (.DIODE(net457));
 sky130_fd_sc_hd__diode_2 ANTENNA_c681_S0 (.DIODE(net457));
 sky130_fd_sc_hd__diode_2 ANTENNA_c674_A3 (.DIODE(net457));
 sky130_fd_sc_hd__diode_2 ANTENNA_c668_A2 (.DIODE(net457));
 sky130_fd_sc_hd__diode_2 ANTENNA_c667_Q (.DIODE(net457));
 sky130_fd_sc_hd__diode_2 ANTENNA_c321_A1 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_A1 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_A0 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_A1 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_A3 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_c191_A3 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_S0 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_A3 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_A3 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_X (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout225_A (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA_c676_A3 (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA_c702_A1 (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA_c696_A0 (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_A2 (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA_c670_X (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA_c723_A3 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_A0 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_A3 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_A2 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_c559_A2 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_c555_A2 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_A3 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_A0 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_A3 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_A1 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_X (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout197_A (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout196_A (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_X (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge855_RESET_B (.DIODE(net537));
 sky130_fd_sc_hd__diode_2 ANTENNA_c747_X (.DIODE(net537));
 sky130_fd_sc_hd__diode_2 ANTENNA_c562_A0 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_A0 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_c434_A2 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_A0 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_S1 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_S1 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_A1 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_A2 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_X (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_A1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_c693_S0 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_c687_A2 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_A1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_c561_A0 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_S0 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_A2 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_A3 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_c180_A0 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_A2 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_X (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge803_Q (.DIODE(net572));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_S1 (.DIODE(net572));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_A2 (.DIODE(net572));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_A3 (.DIODE(net572));
 sky130_fd_sc_hd__diode_2 ANTENNA_c258_S0 (.DIODE(net572));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_C1 (.DIODE(net572));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge804_Q (.DIODE(net573));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_A2 (.DIODE(net573));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_D1 (.DIODE(net573));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_D1 (.DIODE(net573));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_D1 (.DIODE(net573));
 sky130_fd_sc_hd__diode_2 ANTENNA_c286_D1 (.DIODE(net573));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_S1 (.DIODE(net573));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_S1 (.DIODE(net573));
 sky130_fd_sc_hd__diode_2 ANTENNA_c283_SCE (.DIODE(net573));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_S1 (.DIODE(net573));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge835_Q (.DIODE(net607));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_A3 (.DIODE(net607));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_A2 (.DIODE(net607));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_S0 (.DIODE(net607));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_A2 (.DIODE(net607));
 sky130_fd_sc_hd__diode_2 ANTENNA_c446_A2 (.DIODE(net607));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_A2 (.DIODE(net607));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge838_Q (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA_c540_A2 (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA_c533_A3 (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA_c531_S1 (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_S0 (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_A1 (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge846_Q_N (.DIODE(net615));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_A3 (.DIODE(net615));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_A3 (.DIODE(net615));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_S0 (.DIODE(net615));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_A3 (.DIODE(net615));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_S1 (.DIODE(net615));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge879_RESET_B (.DIODE(net621));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge852_X (.DIODE(net621));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge855_Q (.DIODE(net623));
 sky130_fd_sc_hd__diode_2 ANTENNA_c769_A2 (.DIODE(net623));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_S0 (.DIODE(net623));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_A3 (.DIODE(net623));
 sky130_fd_sc_hd__diode_2 ANTENNA_c701_A3 (.DIODE(net623));
 sky130_fd_sc_hd__diode_2 ANTENNA_c686_A3 (.DIODE(net623));
 sky130_fd_sc_hd__diode_2 ANTENNA_c669_C1 (.DIODE(net623));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge856_Q (.DIODE(net625));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_A2 (.DIODE(net625));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_A1 (.DIODE(net625));
 sky130_fd_sc_hd__diode_2 ANTENNA_c615_A3 (.DIODE(net625));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge860_Q (.DIODE(net629));
 sky130_fd_sc_hd__diode_2 ANTENNA_c502_A3 (.DIODE(net629));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_A2 (.DIODE(net629));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_A3 (.DIODE(net629));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_S0 (.DIODE(net629));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_S1 (.DIODE(net629));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_A3 (.DIODE(net629));
 sky130_fd_sc_hd__diode_2 ANTENNA_c235_C1 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_c234_D1 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_c228_D (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_A2 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_A1 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_A2 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_A0 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_c183_A1 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_X (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge861_Q (.DIODE(net630));
 sky130_fd_sc_hd__diode_2 ANTENNA_c373_A3 (.DIODE(net630));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_S1 (.DIODE(net630));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_S0 (.DIODE(net630));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_A2 (.DIODE(net630));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_S0 (.DIODE(net630));
 sky130_fd_sc_hd__diode_2 ANTENNA_c218_A3 (.DIODE(net630));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_A3 (.DIODE(net630));
 sky130_fd_sc_hd__diode_2 ANTENNA_c216_S1 (.DIODE(net630));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge864_Q (.DIODE(net636));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_S0 (.DIODE(net636));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_S0 (.DIODE(net636));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_C1 (.DIODE(net636));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold35_A (.DIODE(net639));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge866_Q (.DIODE(net639));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_SCE (.DIODE(net639));
 sky130_fd_sc_hd__diode_2 ANTENNA_c698_S1 (.DIODE(net639));
 sky130_fd_sc_hd__diode_2 ANTENNA_c696_S0 (.DIODE(net639));
 sky130_fd_sc_hd__diode_2 ANTENNA_c415_A3 (.DIODE(net639));
 sky130_fd_sc_hd__diode_2 ANTENNA_c413_S0 (.DIODE(net639));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge867_Q (.DIODE(net640));
 sky130_fd_sc_hd__diode_2 ANTENNA_c681_S1 (.DIODE(net640));
 sky130_fd_sc_hd__diode_2 ANTENNA_c680_B1 (.DIODE(net640));
 sky130_fd_sc_hd__diode_2 ANTENNA_c677_B1 (.DIODE(net640));
 sky130_fd_sc_hd__diode_2 ANTENNA_c535_S0 (.DIODE(net640));
 sky130_fd_sc_hd__diode_2 ANTENNA_c412_S0 (.DIODE(net640));
 sky130_fd_sc_hd__diode_2 ANTENNA_c411_S0 (.DIODE(net640));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge869_Q (.DIODE(net641));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_S0 (.DIODE(net641));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_A2 (.DIODE(net641));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_A3 (.DIODE(net641));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_A1 (.DIODE(net641));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_A3 (.DIODE(net641));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_A3 (.DIODE(net641));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_A3 (.DIODE(net641));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_S0 (.DIODE(net641));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge871_Q (.DIODE(net642));
 sky130_fd_sc_hd__diode_2 ANTENNA_c767_A1 (.DIODE(net642));
 sky130_fd_sc_hd__diode_2 ANTENNA_c761_A3 (.DIODE(net642));
 sky130_fd_sc_hd__diode_2 ANTENNA_c633_S0 (.DIODE(net642));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_C1 (.DIODE(net642));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_S0 (.DIODE(net642));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_A3 (.DIODE(net642));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_A2 (.DIODE(net642));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge873_Q (.DIODE(net644));
 sky130_fd_sc_hd__diode_2 ANTENNA_c720_A3 (.DIODE(net644));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_A1 (.DIODE(net644));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_A2 (.DIODE(net644));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_S1 (.DIODE(net644));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_B1 (.DIODE(net644));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_A3 (.DIODE(net644));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_A3 (.DIODE(net644));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_S0 (.DIODE(net644));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge879_Q (.DIODE(net649));
 sky130_fd_sc_hd__diode_2 ANTENNA_c766_A2 (.DIODE(net649));
 sky130_fd_sc_hd__diode_2 ANTENNA_c762_A3 (.DIODE(net649));
 sky130_fd_sc_hd__diode_2 ANTENNA_c747_A3 (.DIODE(net649));
 sky130_fd_sc_hd__diode_2 ANTENNA_c746_B1 (.DIODE(net649));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_A2 (.DIODE(net649));
 sky130_fd_sc_hd__diode_2 ANTENNA_c703_A2 (.DIODE(net649));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_A2 (.DIODE(net649));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_S0 (.DIODE(net649));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout212_A (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_A2 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_A0 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA_c183_X (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge881_Q (.DIODE(net650));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_A2 (.DIODE(net650));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_A3 (.DIODE(net650));
 sky130_fd_sc_hd__diode_2 ANTENNA_c350_A3 (.DIODE(net650));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_A2 (.DIODE(net650));
 sky130_fd_sc_hd__diode_2 ANTENNA_c346_S0 (.DIODE(net650));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_S1 (.DIODE(net650));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_A3 (.DIODE(net650));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_C1 (.DIODE(net650));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_S1 (.DIODE(net650));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_A3 (.DIODE(net650));
 sky130_fd_sc_hd__diode_2 ANTENNA_s886_Q_N (.DIODE(net658));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_A3 (.DIODE(net658));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_S1 (.DIODE(net658));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_S0 (.DIODE(net658));
 sky130_fd_sc_hd__diode_2 ANTENNA_c446_A3 (.DIODE(net658));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_A3 (.DIODE(net658));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_S0 (.DIODE(net658));
 sky130_fd_sc_hd__diode_2 ANTENNA_s886_Q (.DIODE(net659));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_S0 (.DIODE(net659));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_S1 (.DIODE(net659));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_A3 (.DIODE(net659));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_S0 (.DIODE(net659));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_A2 (.DIODE(net659));
 sky130_fd_sc_hd__diode_2 ANTENNA_c206_S1 (.DIODE(net659));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_D1 (.DIODE(net659));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold34_A (.DIODE(net661));
 sky130_fd_sc_hd__diode_2 ANTENNA_s888_Q (.DIODE(net661));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_A2 (.DIODE(net661));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_S0 (.DIODE(net661));
 sky130_fd_sc_hd__diode_2 ANTENNA_c311_S0 (.DIODE(net661));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_S0 (.DIODE(net661));
 sky130_fd_sc_hd__diode_2 ANTENNA_c205_S1 (.DIODE(net661));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_S1 (.DIODE(net661));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout245_A (.DIODE(net667));
 sky130_fd_sc_hd__diode_2 ANTENNA_c685_A2 (.DIODE(net667));
 sky130_fd_sc_hd__diode_2 ANTENNA_s894_Q_N (.DIODE(net667));
 sky130_fd_sc_hd__diode_2 ANTENNA_s895_Q_N (.DIODE(net668));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_A3 (.DIODE(net668));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_S0 (.DIODE(net668));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_A3 (.DIODE(net668));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_S0 (.DIODE(net668));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_S1 (.DIODE(net668));
 sky130_fd_sc_hd__diode_2 ANTENNA_s896_Q (.DIODE(net669));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_A2 (.DIODE(net669));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_S0 (.DIODE(net669));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_S0 (.DIODE(net669));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_A2 (.DIODE(net669));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_S0 (.DIODE(net669));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_S1 (.DIODE(net669));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_S1 (.DIODE(net669));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_S1 (.DIODE(net669));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_S1 (.DIODE(net669));
 sky130_fd_sc_hd__diode_2 ANTENNA_s901_Q_N (.DIODE(net674));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A2 (.DIODE(net674));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_S0 (.DIODE(net674));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_A3 (.DIODE(net674));
 sky130_fd_sc_hd__diode_2 ANTENNA_s901_Q (.DIODE(net675));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_A3 (.DIODE(net675));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_A2 (.DIODE(net675));
 sky130_fd_sc_hd__diode_2 ANTENNA_c615_S1 (.DIODE(net675));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_S1 (.DIODE(net675));
 sky130_fd_sc_hd__diode_2 ANTENNA_s904_Q (.DIODE(net678));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_A3 (.DIODE(net678));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_A1 (.DIODE(net678));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_A1 (.DIODE(net678));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_S1 (.DIODE(net678));
 sky130_fd_sc_hd__diode_2 ANTENNA_c482_S0 (.DIODE(net678));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_A2 (.DIODE(net678));
 sky130_fd_sc_hd__diode_2 ANTENNA_c350_S1 (.DIODE(net678));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_S0 (.DIODE(net678));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_S0 (.DIODE(net678));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_S0 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_A1 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_A3 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c190_A2 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_S1 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_S0 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_Q_N (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_s909_Q_N (.DIODE(net681));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_S1 (.DIODE(net681));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_S0 (.DIODE(net681));
 sky130_fd_sc_hd__diode_2 ANTENNA_c369_S1 (.DIODE(net681));
 sky130_fd_sc_hd__diode_2 ANTENNA_c368_S0 (.DIODE(net681));
 sky130_fd_sc_hd__diode_2 ANTENNA_s909_Q (.DIODE(net682));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_D1 (.DIODE(net682));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_A3 (.DIODE(net682));
 sky130_fd_sc_hd__diode_2 ANTENNA_c496_S0 (.DIODE(net682));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_A3 (.DIODE(net682));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_S1 (.DIODE(net682));
 sky130_fd_sc_hd__diode_2 ANTENNA_s911_Q_N (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_S1 (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_S1 (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA_c372_S0 (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA_c371_S1 (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA_s912_Q (.DIODE(net687));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_S0 (.DIODE(net687));
 sky130_fd_sc_hd__diode_2 ANTENNA_c502_S1 (.DIODE(net687));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_S1 (.DIODE(net687));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_S1 (.DIODE(net687));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_S1 (.DIODE(net687));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_S1 (.DIODE(net687));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_S0 (.DIODE(net687));
 sky130_fd_sc_hd__diode_2 ANTENNA_c373_S1 (.DIODE(net687));
 sky130_fd_sc_hd__diode_2 ANTENNA_c372_S1 (.DIODE(net687));
 sky130_fd_sc_hd__diode_2 ANTENNA_s913_Q (.DIODE(net688));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_A3 (.DIODE(net688));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_S1 (.DIODE(net688));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_S0 (.DIODE(net688));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_S0 (.DIODE(net688));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_S1 (.DIODE(net688));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A1 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_D (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_A1 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_A0 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_A0 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_c198_A1 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_Q (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout237_A (.DIODE(net691));
 sky130_fd_sc_hd__diode_2 ANTENNA_c665_SET_B (.DIODE(net691));
 sky130_fd_sc_hd__diode_2 ANTENNA_c669_D1 (.DIODE(net691));
 sky130_fd_sc_hd__diode_2 ANTENNA_c675_S1 (.DIODE(net691));
 sky130_fd_sc_hd__diode_2 ANTENNA_c539_A3 (.DIODE(net691));
 sky130_fd_sc_hd__diode_2 ANTENNA_s916_Q (.DIODE(net691));
 sky130_fd_sc_hd__diode_2 ANTENNA_s917_Q_N (.DIODE(net692));
 sky130_fd_sc_hd__diode_2 ANTENNA_c577_A3 (.DIODE(net692));
 sky130_fd_sc_hd__diode_2 ANTENNA_c535_S1 (.DIODE(net692));
 sky130_fd_sc_hd__diode_2 ANTENNA_c533_S1 (.DIODE(net692));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_S1 (.DIODE(net692));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_S1 (.DIODE(net692));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_S0 (.DIODE(net692));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_S1 (.DIODE(net692));
 sky130_fd_sc_hd__diode_2 ANTENNA_s917_Q (.DIODE(net693));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_A2 (.DIODE(net693));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_A3 (.DIODE(net693));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_A3 (.DIODE(net693));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_S0 (.DIODE(net693));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_S1 (.DIODE(net693));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_S0 (.DIODE(net693));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_D1 (.DIODE(net693));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_S1 (.DIODE(net693));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout236_A (.DIODE(net698));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_A2 (.DIODE(net698));
 sky130_fd_sc_hd__diode_2 ANTENNA_c691_A3 (.DIODE(net698));
 sky130_fd_sc_hd__diode_2 ANTENNA_s921_Q (.DIODE(net698));
 sky130_fd_sc_hd__diode_2 ANTENNA_c372_A3 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_c365_A3 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_A2 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_A2 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_c260_A0 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_D1 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_c118_A2 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_c111_C1 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_c109_X (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net701_A (.DIODE(net701));
 sky130_fd_sc_hd__diode_2 ANTENNA_s924_GCLK (.DIODE(net701));
 sky130_fd_sc_hd__diode_2 ANTENNA_s925_Q_N (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_A2 (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_S1 (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_A3 (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_S1 (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_D1 (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_S1 (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_S1 (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA_s925_Q (.DIODE(net703));
 sky130_fd_sc_hd__diode_2 ANTENNA_c757_A2 (.DIODE(net703));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A2 (.DIODE(net703));
 sky130_fd_sc_hd__diode_2 ANTENNA_c744_A2 (.DIODE(net703));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_A3 (.DIODE(net703));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_A3 (.DIODE(net703));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_S0 (.DIODE(net703));
 sky130_fd_sc_hd__diode_2 ANTENNA_c437_S1 (.DIODE(net703));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout235_A (.DIODE(net710));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_S0 (.DIODE(net710));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_S1 (.DIODE(net710));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_A3 (.DIODE(net710));
 sky130_fd_sc_hd__diode_2 ANTENNA_s930_Q (.DIODE(net710));
 sky130_fd_sc_hd__diode_2 ANTENNA_s933_Q_N (.DIODE(net713));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_A3 (.DIODE(net713));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_A3 (.DIODE(net713));
 sky130_fd_sc_hd__diode_2 ANTENNA_c482_S1 (.DIODE(net713));
 sky130_fd_sc_hd__diode_2 ANTENNA_s933_Q (.DIODE(net714));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_A2 (.DIODE(net714));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_S1 (.DIODE(net714));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_S1 (.DIODE(net714));
 sky130_fd_sc_hd__diode_2 ANTENNA_s936_Q (.DIODE(net717));
 sky130_fd_sc_hd__diode_2 ANTENNA_c762_S0 (.DIODE(net717));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A3 (.DIODE(net717));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A3 (.DIODE(net717));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_A2 (.DIODE(net717));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_S0 (.DIODE(net717));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_S1 (.DIODE(net717));
 sky130_fd_sc_hd__diode_2 ANTENNA_s943_Q_N (.DIODE(net726));
 sky130_fd_sc_hd__diode_2 ANTENNA_c702_A3 (.DIODE(net726));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_A3 (.DIODE(net726));
 sky130_fd_sc_hd__diode_2 ANTENNA_c663_D1 (.DIODE(net726));
 sky130_fd_sc_hd__diode_2 ANTENNA_c544_S1 (.DIODE(net726));
 sky130_fd_sc_hd__diode_2 ANTENNA_c542_S1 (.DIODE(net726));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout191_A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_c344_A1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_A3 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_c190_X (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_s949_Q_N (.DIODE(net732));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_S0 (.DIODE(net732));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_A3 (.DIODE(net732));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_A3 (.DIODE(net732));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_S0 (.DIODE(net732));
 sky130_fd_sc_hd__diode_2 ANTENNA_c587_A3 (.DIODE(net732));
 sky130_fd_sc_hd__diode_2 ANTENNA_c577_S1 (.DIODE(net732));
 sky130_fd_sc_hd__diode_2 ANTENNA_s949_Q (.DIODE(net733));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_S0 (.DIODE(net733));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_S0 (.DIODE(net733));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_S0 (.DIODE(net733));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_S1 (.DIODE(net733));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_S1 (.DIODE(net733));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_S1 (.DIODE(net733));
 sky130_fd_sc_hd__diode_2 ANTENNA_s950_Q_N (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_S1 (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_S1 (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA_c571_S1 (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA_s957_Q (.DIODE(net742));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_S1 (.DIODE(net742));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_S1 (.DIODE(net742));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_S0 (.DIODE(net742));
 sky130_fd_sc_hd__diode_2 ANTENNA_s960_Q (.DIODE(net746));
 sky130_fd_sc_hd__diode_2 ANTENNA_c766_A3 (.DIODE(net746));
 sky130_fd_sc_hd__diode_2 ANTENNA_c614_S0 (.DIODE(net746));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_S0 (.DIODE(net746));
 sky130_fd_sc_hd__diode_2 ANTENNA_c611_S1 (.DIODE(net746));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_S0 (.DIODE(net746));
 sky130_fd_sc_hd__diode_2 ANTENNA_s961_Q (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_A2 (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_A3 (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA_c610_S1 (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_S1 (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_S1 (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_S1 (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA_c677_C1 (.DIODE(net753));
 sky130_fd_sc_hd__diode_2 ANTENNA_s967_Q (.DIODE(net753));
 sky130_fd_sc_hd__diode_2 ANTENNA_c764_S0 (.DIODE(net753));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_S0 (.DIODE(net753));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_S1 (.DIODE(net753));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_S1 (.DIODE(net753));
 sky130_fd_sc_hd__diode_2 ANTENNA_c680_D1 (.DIODE(net753));
 sky130_fd_sc_hd__diode_2 ANTENNA_c676_S1 (.DIODE(net753));
 sky130_fd_sc_hd__diode_2 ANTENNA_s969_Q (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA_c724_A3 (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_A3 (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_S0 (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_S1 (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_S1 (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA_c703_A3 (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_A3 (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_S0 (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA_s976_Q (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_c744_A3 (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_S1 (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_S0 (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_S0 (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_S0 (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_s977_Q (.DIODE(net766));
 sky130_fd_sc_hd__diode_2 ANTENNA_c768_S0 (.DIODE(net766));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_A3 (.DIODE(net766));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_S0 (.DIODE(net766));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_S1 (.DIODE(net766));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_S1 (.DIODE(net766));
 sky130_fd_sc_hd__diode_2 ANTENNA_s981_Q_N (.DIODE(net769));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_S1 (.DIODE(net769));
 sky130_fd_sc_hd__diode_2 ANTENNA_c742_D1 (.DIODE(net769));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_S1 (.DIODE(net769));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_SET_B (.DIODE(net769));
 sky130_fd_sc_hd__diode_2 ANTENNA_s985_Q (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_c767_S0 (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_c763_S1 (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_S1 (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_S1 (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_S1 (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_S1 (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_c230_D1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c220_A1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c215_A2 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_A2 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_S0 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c206_A1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_A3 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_X (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_A0 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_A2 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_S1 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_A1 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_c216_A1 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_A2 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_c208_S1 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_A0 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_X (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_c257_A0 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_B1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_A0 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_c208_A2 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_A3 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_c206_X (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_X (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA_c669_B1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA_c529_SCE (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA_c398_C1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA_c267_D1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_A1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_X (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_S1 (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_A1 (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout256_A (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_X (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA_c661_B1 (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA_c530_RESET_B (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_X (.DIODE(net781));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_A2 (.DIODE(net781));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_A3 (.DIODE(net781));
 sky130_fd_sc_hd__diode_2 ANTENNA_c138_A1 (.DIODE(net781));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_X (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_A1 (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_S1 (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_C1 (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout249_A (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout248_A (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_X (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone3_C1 (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_C1 (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_X (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_S0 (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_c148_A2 (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_c140_A0 (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_c138_A2 (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_A1 (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_X (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c203_A0 (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_A3 (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_A2 (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_X (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA_c532_A2 (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA_c531_A0 (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_B1 (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone3_A2 (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_X (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_A3 (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_A2 (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA_c143_B1 (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_B1 (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_A1 (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_A2 (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_A2 (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_X (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_c274_A1 (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_c265_A1 (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_c134_C1 (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_X (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_A1 (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_A1 (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_X (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c235_B1 (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_A2 (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c194_A3 (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c191_A2 (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_D1 (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c159_S0 (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_D1 (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c130_S0 (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c117_A2 (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_X (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_c430_A0 (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_c427_A0 (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout257_A (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_X (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_A1 (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA_c203_A2 (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_A3 (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_X (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_D1 (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_A1 (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone3_A1 (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_X (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_c148_A0 (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_A1 (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_X (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_c563_A0 (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_A2 (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_A2 (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_A3 (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_c295_C1 (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_c286_C1 (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_A2 (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_X (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_A1 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_S0 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c158_B1 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_input30_X (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_A0 (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_A1 (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_input31_X (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_A0 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_A3 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_B1 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_D (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_A0 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_S0 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_B1 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_A3 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_A3 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_A2 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_input32_X (.DIODE(net809));
 sky130_fd_sc_hd__diode_2 ANTENNA_c431_A0 (.DIODE(net809));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_A1 (.DIODE(net809));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_A2 (.DIODE(net809));
 sky130_fd_sc_hd__diode_2 ANTENNA_input33_X (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_A0 (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_A1 (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_c311_A0 (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_c221_A0 (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_c220_D1 (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_c183_S1 (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_A1 (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_C1 (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_input34_X (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_A0 (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_A1 (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_A2 (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_c286_B1 (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_A2 (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_S0 (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_B1 (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_input35_X (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_A0 (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_c272_B1 (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_c264_D1 (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_input36_X (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_A1 (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c555_A0 (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_A1 (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_A3 (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_B1 (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_A1 (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_A3 (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c158_C1 (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_input37_X (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_A0 (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_A0 (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_A0 (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout255_A (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_input38_X (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_c765_A1 (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_A1 (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_A3 (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_input39_X (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_A1 (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_A2 (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_input40_X (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c218_A0 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c203_A1 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_A2 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_S0 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_B1 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_input41_X (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c222_A0 (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c220_B1 (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_input42_X (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_A0 (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_c183_S0 (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_input43_X (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_c263_A1 (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_c221_S0 (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_c205_A2 (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_c180_A2 (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_C1 (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_c107_A3 (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_input44_X (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_c183_A2 (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_A0 (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_A1 (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout254_A (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_input46_X (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_A3 (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout253_A (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout252_A (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_input47_X (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_input48_X (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_A1 (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_A1 (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_input49_X (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_A0 (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_c182_A2 (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_c180_S0 (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_A2 (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_input50_X (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_A3 (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_A1 (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_A3 (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_c182_A3 (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_c180_A3 (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_c128_A3 (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_input51_X (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_S0 (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_A1 (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_input52_X (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_S0 (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_A3 (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_A1 (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_A1 (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_A2 (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_input55_X (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_A0 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_A3 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_C1 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_input56_X (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_A2 (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_c120_S1 (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_c118_D1 (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_input57_X (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_A0 (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_A3 (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_input60_X (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c212_A0 (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_S0 (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_RESET_B (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_C1 (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_input61_X (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_c256_A0 (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_A3 (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_input62_X (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c241_A1 (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_A2 (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c194_S0 (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_A2 (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c184_A2 (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_A3 (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c100_A3 (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_input64_X (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_A0 (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_A3 (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_c208_A3 (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_input65_X (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_A0 (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_S0 (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_input66_X (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_A3 (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_A3 (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_S0 (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c259_S0 (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_A1 (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c120_S0 (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c105_A3 (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c272_D1 (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_input68_X (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_c416_A0 (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_c407_A2 (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_c397_B1 (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_c266_B1 (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_c265_C1 (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_c148_S1 (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_c138_B1 (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_input69_X (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_c229_B1 (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_A1 (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_A2 (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_c222_A2 (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_c198_S1 (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_input71_X (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_A0 (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_c494_A2 (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_A1 (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_A0 (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_A2 (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_A3 (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_c128_S0 (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_c126_A2 (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_c123_A2 (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_c110_A2 (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_input72_X (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_A1 (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_A1 (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c119_C1 (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c111_A1 (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c109_S1 (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c102_A2 (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c101_S0 (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c100_S0 (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_input77_X (.DIODE(net854));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_A3 (.DIODE(net854));
 sky130_fd_sc_hd__diode_2 ANTENNA_c215_A3 (.DIODE(net854));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_A3 (.DIODE(net854));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_A1 (.DIODE(net854));
 sky130_fd_sc_hd__diode_2 ANTENNA_c205_S0 (.DIODE(net854));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_S1 (.DIODE(net854));
 sky130_fd_sc_hd__diode_2 ANTENNA_c198_A2 (.DIODE(net854));
 sky130_fd_sc_hd__diode_2 ANTENNA_c128_A2 (.DIODE(net854));
 sky130_fd_sc_hd__diode_2 ANTENNA_c115_A2 (.DIODE(net854));
 sky130_fd_sc_hd__diode_2 ANTENNA_input78_X (.DIODE(net855));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_A1 (.DIODE(net855));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_A0 (.DIODE(net855));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_A2 (.DIODE(net855));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_A2 (.DIODE(net855));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_A3 (.DIODE(net855));
 sky130_fd_sc_hd__diode_2 ANTENNA_c366_A1 (.DIODE(net855));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_A3 (.DIODE(net855));
 sky130_fd_sc_hd__diode_2 ANTENNA_c231_A3 (.DIODE(net855));
 sky130_fd_sc_hd__diode_2 ANTENNA_c104_S0 (.DIODE(net855));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout251_A (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_input79_X (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_A1 (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_A1 (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_input87_X (.DIODE(net864));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_A0 (.DIODE(net864));
 sky130_fd_sc_hd__diode_2 ANTENNA_c346_A1 (.DIODE(net864));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_A2 (.DIODE(net864));
 sky130_fd_sc_hd__diode_2 ANTENNA_c208_S0 (.DIODE(net864));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_S0 (.DIODE(net864));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_A1 (.DIODE(net864));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_S0 (.DIODE(net864));
 sky130_fd_sc_hd__diode_2 ANTENNA_c198_S0 (.DIODE(net864));
 sky130_fd_sc_hd__diode_2 ANTENNA_input88_X (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_A1 (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_A0 (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_A1 (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_A1 (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_A3 (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_A0 (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c222_S1 (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c220_C1 (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c103_A2 (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c100_S1 (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone17_A (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout247_A (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_input90_X (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_A0 (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_input95_X (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_c370_A3 (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_A1 (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_c261_A1 (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_c101_S1 (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_input99_X (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_A0 (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_A1 (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_A2 (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_A2 (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA_c222_S0 (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA_c220_A2 (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA_c105_S1 (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA_c103_S1 (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA_c101_A3 (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA_c100_A0 (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout190_A (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_output103_A (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c768_A1 (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c759_A2 (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_X (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_output105_A (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_s963_Q (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_A2 (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_S1 (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_S0 (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_A3 (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_output108_A (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge840_Q (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_c764_A3 (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_A3 (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_A3 (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_output109_A (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_s964_Q (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_c767_A2 (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_S0 (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_S0 (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_S0 (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_S1 (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_S1 (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_output110_A (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_s979_Q (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_c767_A3 (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_c764_S1 (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_c763_S0 (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_S0 (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_output111_A (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_s952_Q (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_c762_S1 (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_S1 (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_S0 (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_A2 (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_S0 (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_S1 (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_S1 (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_S1 (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_S1 (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_output113_A (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge851_Q (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c633_A3 (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_S0 (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_S1 (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_output114_A (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge872_Q_N (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_S0 (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_A1 (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c482_A3 (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_output117_A (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge826_Q (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c763_A1 (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c614_A1 (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout224_A (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_A0 (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_c222_X (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_output119_A (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge868_Q (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_A3 (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_A3 (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_S0 (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_S0 (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_S1 (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_S1 (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap244_A (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_s895_Q (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_S0 (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_S0 (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_output126_A (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_s958_Q (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_S1 (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_c614_A3 (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_c610_S0 (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_output127_A (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_s945_Q (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c614_A2 (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_A2 (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_S0 (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_S0 (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c557_C1 (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c556_S1 (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c549_S1 (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout246_A (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_s894_Q (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_S0 (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_A3 (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net909_A (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_c561_X (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_output135_A (.DIODE(net912));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_A1 (.DIODE(net912));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_A1 (.DIODE(net912));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_S0 (.DIODE(net912));
 sky130_fd_sc_hd__diode_2 ANTENNA_c257_S1 (.DIODE(net912));
 sky130_fd_sc_hd__diode_2 ANTENNA_c229_D1 (.DIODE(net912));
 sky130_fd_sc_hd__diode_2 ANTENNA_c112_D1 (.DIODE(net912));
 sky130_fd_sc_hd__diode_2 ANTENNA_c109_A2 (.DIODE(net912));
 sky130_fd_sc_hd__diode_2 ANTENNA_c103_X (.DIODE(net912));
 sky130_fd_sc_hd__diode_2 ANTENNA_output138_A (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge870_Q (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_A2 (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_A2 (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_S0 (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_A3 (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_A3 (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_S0 (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_c416_S0 (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_output139_A (.DIODE(net916));
 sky130_fd_sc_hd__diode_2 ANTENNA_s903_Q (.DIODE(net916));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_A3 (.DIODE(net916));
 sky130_fd_sc_hd__diode_2 ANTENNA_c502_S0 (.DIODE(net916));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_S0 (.DIODE(net916));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_A3 (.DIODE(net916));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_S0 (.DIODE(net916));
 sky130_fd_sc_hd__diode_2 ANTENNA_c344_S1 (.DIODE(net916));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net917_A (.DIODE(net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_X (.DIODE(net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_output143_A (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge880_Q (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_A3 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_A2 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_S0 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_S0 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_C1 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_A2 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_output149_A (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_c260_A2 (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_c131_B1 (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_c130_X (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer7_A (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout221_A (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout220_A (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c138_X (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_output157_A (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge839_Q (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_S0 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c350_A2 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_A0 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c231_S1 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c216_S0 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout228_A (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_output158_A (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c104_X (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_output163_A (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_A1 (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_A1 (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_S1 (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_A0 (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_A3 (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_SCD (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_A1 (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_c182_X (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_output164_A (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c258_A0 (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c131_A2 (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c124_A2 (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c122_A1 (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c121_A2 (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c118_X (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_output166_A (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_A0 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c258_A1 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c190_A0 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_S1 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_A2 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c184_S0 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c182_A1 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c180_X (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_output170_A (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge854_Q (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_A1 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_A3 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_B1 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_A2 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_A3 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_S0 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_output179_A (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge818_Q (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_S0 (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_A1 (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_c323_A1 (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_c241_D1 (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_output180_A (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c263_A3 (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c228_SET_B (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_S0 (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c221_A2 (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_A0 (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c216_A2 (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_A3 (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_X (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout184_X (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_A1 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_A1 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_A2 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c424_A2 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c437_A2 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_A3 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_A1 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_A1 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_A1 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_A3 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout186_X (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c538_A2 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c536_A1 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c537_A0 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c530_SCE (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c413_A2 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c416_A1 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_A3 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c415_A0 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c414_A0 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c528_SCE (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout187_X (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_A0 (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_A1 (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c681_A3 (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_A1 (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c410_A0 (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c403_A3 (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c402_S0 (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c401_A2 (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c399_SCD (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c409_A2 (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout188_X (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c665_SCD (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_A3 (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout187_A (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c747_A1 (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_A1 (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c613_A1 (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_A1 (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_A1 (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_SCD (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout189_X (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c687_A1 (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_A2 (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_A3 (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c427_S1 (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_A2 (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_A0 (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_A2 (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_A1 (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_SCE (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_RESET_B (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout190_X (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_A3 (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_A3 (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_A2 (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_A0 (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c430_A1 (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c366_A3 (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_A3 (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c313_A3 (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_A1 (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_S1 (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout191_X (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_A0 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_A3 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c216_A3 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_A1 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c212_A3 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_A2 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_S0 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c194_A2 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_S1 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_A2 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c660_D1 (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout193_X (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_c664_A1 (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_A1 (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_A2 (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_c691_A2 (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout194_X (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_C1 (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_c297_A3 (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_C1 (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_C1 (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_output144_A (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_A2 (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_A1 (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_A0 (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_A1 (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_A2 (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout195_X (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_A1 (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_A1 (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c402_A2 (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_A0 (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_A0 (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_A1 (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_A0 (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_A1 (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_A2 (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_A1 (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout196_X (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_A1 (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_A2 (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_A1 (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_S0 (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_A0 (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_A1 (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_A2 (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_D1 (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_B1 (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_S1 (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout197_X (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_c745_A1 (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_A2 (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_A0 (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A2 (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_A3 (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_c611_A3 (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_A0 (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_A2 (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout199_X (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_c410_S0 (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout198_A (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_A3 (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_c558_A2 (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_A2 (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout200_X (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout199_A (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_A0 (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_A0 (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_A2 (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_A2 (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_A2 (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_A0 (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout201_X (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_A2 (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_A0 (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_A3 (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_A2 (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_A1 (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_A2 (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_A2 (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_A2 (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_A2 (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_c313_A2 (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout202_X (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c555_A1 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_S0 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_B1 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c434_A0 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_A2 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_A1 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_C1 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c297_S0 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_D1 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_B1 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout205_X (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c397_A1 (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout204_A (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_A2 (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_A1 (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_D1 (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout208_X (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c368_A1 (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c372_A0 (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_A3 (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c340_A3 (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_A0 (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c203_S0 (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_A1 (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c235_A2 (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_A3 (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_S0 (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_A1 (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout209_X (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_A2 (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_S1 (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_S1 (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_c313_S0 (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_A3 (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_A3 (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_A3 (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_A3 (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout208_A (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout212_X (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_A2 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_A1 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_S0 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c191_A1 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c190_A1 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_A3 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_S0 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c184_A3 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_SCE (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c208_A1 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout213_X (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_A2 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_A0 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_A2 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_B1 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_A3 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_S1 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_S1 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_S1 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c159_S1 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c182_S0 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout214_X (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_A2 (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_A2 (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c286_A1 (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_S0 (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout213_A (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_C1 (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout215_X (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_B1 (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_A2 (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_A3 (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_A3 (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout216_X (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c427_A1 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c400_D1 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c311_A2 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c297_A2 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c265_D1 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c264_C1 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_S1 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_A0 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone28_A (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout217_X (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_output133_A (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_A1 (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_S0 (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c587_A1 (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout215_A (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout216_A (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c269_D1 (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout218_X (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_A0 (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c400_B1 (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_A3 (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_A3 (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_S0 (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_C1 (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_S1 (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_D1 (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_A0 (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout219_X (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c700_A2 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c686_A0 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c560_SCD (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_A1 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c265_A2 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout218_A (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout220_X (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_A0 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_A3 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c143_C1 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_B1 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c140_S1 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout221_X (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_A2 (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c582_A2 (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c560_RESET_B (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_A2 (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_A2 (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout223_X (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_A1 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c685_A0 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_A2 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_D1 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c431_A1 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c427_A3 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_A1 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c434_A3 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_A3 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_S0 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout224_X (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_A1 (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_A2 (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_A2 (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_output118_A (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c364_A3 (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_A2 (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c231_A2 (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c228_RESET_B (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_S1 (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_A3 (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout225_X (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c671_C1 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c673_S0 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c674_S1 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c675_A2 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_A2 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c766_A0 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_A1 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_S0 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_A3 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_A0 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer19_A (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone18_A (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout227_X (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_A3 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_A2 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout226_A (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout228_X (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_c761_A1 (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_A1 (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_A3 (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_A2 (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_A1 (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_A1 (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_c236_B1 (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_c121_B1 (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_c110_D1 (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_c108_S1 (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout229_X (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c543_A0 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c539_A2 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c535_A3 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c536_A2 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c537_A2 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_A0 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_A2 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_A0 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c587_A2 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_A2 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout232_X (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_A3 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c691_S0 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_S1 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c686_S1 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_S1 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c685_S1 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_S1 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_A3 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A3 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_S0 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout233_X (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_S0 (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_A2 (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_c700_S0 (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_S0 (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_S1 (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_S1 (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_S0 (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_S0 (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_c685_S0 (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_S0 (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap234_X (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_A3 (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_S0 (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_S1 (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_S1 (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_S0 (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_S0 (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout235_X (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_A3 (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_S0 (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_S1 (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_S0 (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_S0 (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_S1 (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_S1 (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_D1 (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_S1 (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c458_S1 (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout236_X (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_c560_SET_B (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_A3 (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_c430_S1 (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_c431_S0 (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_c555_S0 (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_S0 (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_S0 (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_S0 (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_c561_S1 (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_c563_S0 (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout237_X (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c660_C1 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c662_D1 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c668_D1 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c661_D1 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c416_S1 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c530_SET_B (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c415_S1 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c414_S1 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c413_S1 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c412_S1 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout239_X (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c542_A2 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c545_S1 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout238_A (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_S0 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_S1 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_S0 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_S1 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout240_X (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_D1 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_S1 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_S1 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_S1 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c321_S1 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_S1 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_S1 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_S0 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_S1 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_S0 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout241_X (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_A3 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_S0 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_A3 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_S0 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout240_A (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout243_X (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_S1 (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_S0 (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_A3 (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_S1 (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_c323_A3 (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_A3 (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_S0 (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_A3 (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_S0 (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_S1 (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap244_X (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_output121_A (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_S0 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A1 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_A3 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout245_X (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c665_SCE (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c662_C1 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c661_C1 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c557_B1 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_D1 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c532_S1 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c398_D1 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c283_SET_B (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_A1 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_S1 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout246_X (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c554_C1 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_S1 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_SCE (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_output129_A (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A2 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_A3 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_S0 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_A3 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_S0 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_A2 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone3_D1 (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_D1 (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout247_X (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_c664_A2 (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_A0 (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_c148_A3 (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout249_X (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c760_A2 (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c660_A2 (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_S0 (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c554_A1 (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_A3 (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_B1 (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_B1 (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout250_X (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_A1 (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_A3 (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_S1 (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c134_D1 (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_S0 (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_D1 (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_A0 (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c158_D1 (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_D1 (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout251_X (.DIODE(net1028));
 sky130_fd_sc_hd__diode_2 ANTENNA_c685_A1 (.DIODE(net1028));
 sky130_fd_sc_hd__diode_2 ANTENNA_c542_A0 (.DIODE(net1028));
 sky130_fd_sc_hd__diode_2 ANTENNA_c408_A1 (.DIODE(net1028));
 sky130_fd_sc_hd__diode_2 ANTENNA_c274_S1 (.DIODE(net1028));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout250_A (.DIODE(net1028));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout252_X (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_A2 (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_A2 (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_A1 (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_A1 (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_A0 (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_S0 (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_A1 (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_A1 (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_A1 (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_c101_A2 (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout253_X (.DIODE(net1030));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_A2 (.DIODE(net1030));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_A0 (.DIODE(net1030));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_A2 (.DIODE(net1030));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_S1 (.DIODE(net1030));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_A0 (.DIODE(net1030));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout254_X (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_c686_A2 (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_c633_A2 (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_SCD (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_B1 (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_S1 (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_c222_A3 (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_A0 (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_C1 (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_c140_S0 (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_A2 (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout255_X (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A0 (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_A1 (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_c723_A0 (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_A0 (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_c698_A3 (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_A3 (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_A2 (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_A2 (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_c232_C1 (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_c112_B1 (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout256_X (.DIODE(net1033));
 sky130_fd_sc_hd__diode_2 ANTENNA_c399_RESET_B (.DIODE(net1033));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_A3 (.DIODE(net1033));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_S1 (.DIODE(net1033));
 sky130_fd_sc_hd__diode_2 ANTENNA_c266_C1 (.DIODE(net1033));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_A0 (.DIODE(net1033));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_S0 (.DIODE(net1033));
 sky130_fd_sc_hd__diode_2 ANTENNA_c148_S0 (.DIODE(net1033));
 sky130_fd_sc_hd__diode_2 ANTENNA_c134_A1 (.DIODE(net1033));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_A0 (.DIODE(net1033));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_A3 (.DIODE(net1033));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout257_X (.DIODE(net1034));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_A3 (.DIODE(net1034));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_A1 (.DIODE(net1034));
 sky130_fd_sc_hd__diode_2 ANTENNA_c159_A1 (.DIODE(net1034));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_A1 (.DIODE(net1034));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_A2 (.DIODE(net1034));
 sky130_fd_sc_hd__diode_2 ANTENNA_c262_A2 (.DIODE(net1034));
 sky130_fd_sc_hd__diode_2 ANTENNA_c256_S1 (.DIODE(net1034));
 sky130_fd_sc_hd__diode_2 ANTENNA_c226_A3 (.DIODE(net1034));
 sky130_fd_sc_hd__diode_2 ANTENNA_c111_D1 (.DIODE(net1034));
 sky130_fd_sc_hd__diode_2 ANTENNA_c107_S1 (.DIODE(net1034));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout258_X (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_A2 (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_B1 (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA_c267_B1 (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_B1 (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_S0 (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_A2 (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_A2 (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_A3 (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_D (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA_c101_A1 (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout259_X (.DIODE(net1036));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_A1 (.DIODE(net1036));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_A2 (.DIODE(net1036));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_A1 (.DIODE(net1036));
 sky130_fd_sc_hd__diode_2 ANTENNA_c613_A2 (.DIODE(net1036));
 sky130_fd_sc_hd__diode_2 ANTENNA_c528_RESET_B (.DIODE(net1036));
 sky130_fd_sc_hd__diode_2 ANTENNA_c430_A2 (.DIODE(net1036));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout258_A (.DIODE(net1036));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_15_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_14_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_13_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_12_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_11_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_10_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_9_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_8_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_7_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_6_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_5_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_4_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_3_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_2_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_1_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_0_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_X (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c228_CLK_N (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c237_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge813_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge837_GATE_N (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge842_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge858_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge877_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge878_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s907_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s908_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_0_0_clk_X (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge818_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge839_GATE (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge845_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge861_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge881_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s891_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s892_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s893_GATE_N (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s901_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s903_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s904_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s905_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s906_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_1_0_clk_X (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge848_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s909_GATE_N (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s910_GATE_N (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s911_GATE (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s912_GATE_N (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s913_GATE_N (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s934_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s935_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s936_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s937_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s938_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_2_0_clk_X (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge828_GATE_N (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge856_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge860_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge868_GATE_N (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge869_GATE (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge872_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge880_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s902_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s932_SLEEP_B (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s933_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_3_0_clk_X (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_CLK_N (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge803_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge829_GATE_N (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge854_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s885_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s886_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s888_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s890_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s898_GATE_N (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s899_GATE (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_4_0_clk_X (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge797_CLK_N (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge846_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s887_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s889_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s895_GATE (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s897_GATE_N (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s900_SLEEP_B (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_5_0_clk_X (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge835_GATE_N (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge844_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge874_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s896_GATE_N (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s923_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s924_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s926_GATE_N (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s927_GATE (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s928_GATE_N (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s930_GATE_N (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s931_GATE (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_6_0_clk_X (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c277_CLK_N (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c283_CLK_N (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c399_CLK_N (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_CLK_N (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge804_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge816_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge836_GATE_N (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s894_GATE_N (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s914_GATE_N (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s918_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s919_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_7_0_clk_X (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge826_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge840_GATE (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge843_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge851_CLK_N (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge857_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge862_GATE_N (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge871_GATE (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge883_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s958_GATE_N (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s961_GATE_N (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s962_GATE_N (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s963_GATE (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s964_SLEEP_B (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s965_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s966_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s989_GATE_N (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_8_0_clk_X (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge792_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge873_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s929_GATE_N (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s950_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s952_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s953_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s954_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s955_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s956_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s957_GATE_N (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s959_GATE (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s960_GATE_N (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_9_0_clk_X (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_CLK_N (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge827_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s970_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s974_GATE_N (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s975_GATE (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s976_GATE_N (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s977_GATE_N (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s978_GATE_N (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s979_GATE (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s980_SLEEP_B (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s981_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s982_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s983_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_11_0_clk_X (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge805_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge838_GATE (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge864_GATE (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge870_GATE (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge884_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s917_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s920_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s921_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s922_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s925_GATE_N (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s946_GATE_N (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s947_GATE (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_12_0_clk_X (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c560_CLK_N (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge841_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge866_GATE_N (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge875_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge879_CLK_N (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s948_SLEEP_B (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s949_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s951_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s967_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s968_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s969_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s971_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s972_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s973_GATE_N (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_14_0_clk_X (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c665_CLK_N (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c666_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c667_CLK_N (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge855_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge867_GATE_N (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge876_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s940_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s941_GATE_N (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s942_GATE_N (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s943_GATE (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s945_GATE_N (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_15_0_clk_X (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c703_S0 (.DIODE(clknet_1_1__leaf_net756));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_S0 (.DIODE(clknet_1_1__leaf_net756));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_S1 (.DIODE(clknet_1_1__leaf_net756));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net756_X (.DIODE(clknet_1_1__leaf_net756));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_A1 (.DIODE(clknet_1_0__leaf_net404));
 sky130_fd_sc_hd__diode_2 ANTENNA_c742_A2 (.DIODE(clknet_1_0__leaf_net404));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A0 (.DIODE(clknet_1_0__leaf_net404));
 sky130_fd_sc_hd__diode_2 ANTENNA_c763_A0 (.DIODE(clknet_1_0__leaf_net404));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net404_X (.DIODE(clknet_1_0__leaf_net404));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_A0 (.DIODE(clknet_1_1__leaf_net404));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_A1 (.DIODE(clknet_1_1__leaf_net404));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_A1 (.DIODE(clknet_1_1__leaf_net404));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_A0 (.DIODE(clknet_1_1__leaf_net404));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net404_X (.DIODE(clknet_1_1__leaf_net404));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_A2 (.DIODE(clknet_1_0__leaf_net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_A2 (.DIODE(clknet_1_0__leaf_net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_A3 (.DIODE(clknet_1_0__leaf_net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c615_A1 (.DIODE(clknet_1_0__leaf_net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A1 (.DIODE(clknet_1_0__leaf_net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net908_X (.DIODE(clknet_1_0__leaf_net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_A3 (.DIODE(clknet_1_0__leaf_net402));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_A0 (.DIODE(clknet_1_0__leaf_net402));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_A1 (.DIODE(clknet_1_0__leaf_net402));
 sky130_fd_sc_hd__diode_2 ANTENNA_c765_A2 (.DIODE(clknet_1_0__leaf_net402));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net402_X (.DIODE(clknet_1_0__leaf_net402));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_A1 (.DIODE(clknet_1_1__leaf_net402));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_A1 (.DIODE(clknet_1_1__leaf_net402));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_A1 (.DIODE(clknet_1_1__leaf_net402));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_A1 (.DIODE(clknet_1_1__leaf_net402));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net402_X (.DIODE(clknet_1_1__leaf_net402));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_A1 (.DIODE(clknet_1_0__leaf_net361));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_A0 (.DIODE(clknet_1_0__leaf_net361));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_A3 (.DIODE(clknet_1_0__leaf_net361));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_A1 (.DIODE(clknet_1_0__leaf_net361));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_A2 (.DIODE(clknet_1_0__leaf_net361));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net361_X (.DIODE(clknet_1_0__leaf_net361));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_C1 (.DIODE(clknet_1_1__leaf_net361));
 sky130_fd_sc_hd__diode_2 ANTENNA_c566_A2 (.DIODE(clknet_1_1__leaf_net361));
 sky130_fd_sc_hd__diode_2 ANTENNA_c582_A0 (.DIODE(clknet_1_1__leaf_net361));
 sky130_fd_sc_hd__diode_2 ANTENNA_c696_A2 (.DIODE(clknet_1_1__leaf_net361));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net361_X (.DIODE(clknet_1_1__leaf_net361));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_A3 (.DIODE(clknet_1_0__leaf_net476));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_A2 (.DIODE(clknet_1_0__leaf_net476));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_A0 (.DIODE(clknet_1_0__leaf_net476));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_A0 (.DIODE(clknet_1_0__leaf_net476));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_A1 (.DIODE(clknet_1_0__leaf_net476));
 sky130_fd_sc_hd__diode_2 ANTENNA_c768_A0 (.DIODE(clknet_1_0__leaf_net476));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net476_X (.DIODE(clknet_1_0__leaf_net476));
 sky130_fd_sc_hd__diode_2 ANTENNA_c562_A3 (.DIODE(clknet_1_0__leaf_net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_c564_A2 (.DIODE(clknet_1_0__leaf_net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_A1 (.DIODE(clknet_1_0__leaf_net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_A1 (.DIODE(clknet_1_0__leaf_net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_A2 (.DIODE(clknet_1_0__leaf_net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net909_X (.DIODE(clknet_1_0__leaf_net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_A2 (.DIODE(clknet_1_1__leaf_net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_output132_A (.DIODE(clknet_1_1__leaf_net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net909_X (.DIODE(clknet_1_1__leaf_net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_S0 (.DIODE(clknet_1_0__leaf_net701));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_S1 (.DIODE(clknet_1_0__leaf_net701));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_A3 (.DIODE(clknet_1_0__leaf_net701));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_S0 (.DIODE(clknet_1_0__leaf_net701));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_S0 (.DIODE(clknet_1_0__leaf_net701));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_S0 (.DIODE(clknet_1_0__leaf_net701));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net701_X (.DIODE(clknet_1_0__leaf_net701));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_A3 (.DIODE(clknet_1_1__leaf_net701));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_A3 (.DIODE(clknet_1_1__leaf_net701));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_S0 (.DIODE(clknet_1_1__leaf_net701));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_A3 (.DIODE(clknet_1_1__leaf_net701));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_A2 (.DIODE(clknet_1_1__leaf_net701));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_A3 (.DIODE(clknet_1_1__leaf_net701));
 sky130_fd_sc_hd__diode_2 ANTENNA_c739_A3 (.DIODE(clknet_1_1__leaf_net701));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_A1 (.DIODE(clknet_1_1__leaf_net701));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net701_X (.DIODE(clknet_1_1__leaf_net701));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_A2 (.DIODE(clknet_1_0__leaf_net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_c458_A3 (.DIODE(clknet_1_0__leaf_net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_A1 (.DIODE(clknet_1_0__leaf_net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_A2 (.DIODE(clknet_1_0__leaf_net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_A1 (.DIODE(clknet_1_0__leaf_net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_SCD (.DIODE(clknet_1_0__leaf_net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_A0 (.DIODE(clknet_1_0__leaf_net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net917_X (.DIODE(clknet_1_0__leaf_net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_A3 (.DIODE(clknet_1_1__leaf_net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_A2 (.DIODE(clknet_1_1__leaf_net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_A2 (.DIODE(clknet_1_1__leaf_net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_A2 (.DIODE(clknet_1_1__leaf_net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_A0 (.DIODE(clknet_1_1__leaf_net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_A1 (.DIODE(clknet_1_1__leaf_net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_c762_A2 (.DIODE(clknet_1_1__leaf_net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_c764_A1 (.DIODE(clknet_1_1__leaf_net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_c768_A2 (.DIODE(clknet_1_1__leaf_net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_output140_A (.DIODE(clknet_1_1__leaf_net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net917_X (.DIODE(clknet_1_1__leaf_net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_S0 (.DIODE(clknet_1_0__leaf_net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_A1 (.DIODE(clknet_1_0__leaf_net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_A3 (.DIODE(clknet_1_0__leaf_net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_output156_A (.DIODE(clknet_1_0__leaf_net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net933_X (.DIODE(clknet_1_0__leaf_net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c372_A1 (.DIODE(clknet_1_0__leaf_net226));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_A1 (.DIODE(clknet_1_0__leaf_net226));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_A1 (.DIODE(clknet_1_0__leaf_net226));
 sky130_fd_sc_hd__diode_2 ANTENNA_c761_A2 (.DIODE(clknet_1_0__leaf_net226));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net226_X (.DIODE(clknet_1_0__leaf_net226));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_A3 (.DIODE(clknet_1_1__leaf_net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_A1 (.DIODE(clknet_1_1__leaf_net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_A1 (.DIODE(clknet_1_1__leaf_net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_A1 (.DIODE(clknet_1_1__leaf_net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_output120_A (.DIODE(clknet_1_1__leaf_net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net897_X (.DIODE(clknet_1_1__leaf_net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_A1 (.DIODE(clknet_1_0__leaf_net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_A1 (.DIODE(clknet_1_0__leaf_net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_A3 (.DIODE(clknet_1_0__leaf_net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_B1 (.DIODE(clknet_1_0__leaf_net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_output116_A (.DIODE(clknet_1_0__leaf_net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net893_X (.DIODE(clknet_1_0__leaf_net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c231_A0 (.DIODE(clknet_1_0__leaf_net99));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_A0 (.DIODE(clknet_1_0__leaf_net99));
 sky130_fd_sc_hd__diode_2 ANTENNA_c364_A2 (.DIODE(clknet_1_0__leaf_net99));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_A0 (.DIODE(clknet_1_0__leaf_net99));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_A3 (.DIODE(clknet_1_0__leaf_net99));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net99_X (.DIODE(clknet_1_0__leaf_net99));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_A2 (.DIODE(clknet_1_0__leaf_net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_A3 (.DIODE(clknet_1_0__leaf_net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_A2 (.DIODE(clknet_1_0__leaf_net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_output142_A (.DIODE(clknet_1_0__leaf_net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net919_X (.DIODE(clknet_1_0__leaf_net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net100_A (.DIODE(clknet_0_net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net100_A (.DIODE(clknet_0_net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net100_X (.DIODE(clknet_0_net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c236_A2 (.DIODE(clknet_1_0__leaf_net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_A3 (.DIODE(clknet_1_0__leaf_net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_A0 (.DIODE(clknet_1_0__leaf_net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_A1 (.DIODE(clknet_1_0__leaf_net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_S0 (.DIODE(clknet_1_0__leaf_net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_A0 (.DIODE(clknet_1_0__leaf_net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_A2 (.DIODE(clknet_1_0__leaf_net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net100_X (.DIODE(clknet_1_0__leaf_net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_A2 (.DIODE(clknet_1_1__leaf_net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_S0 (.DIODE(clknet_1_1__leaf_net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_A1 (.DIODE(clknet_1_1__leaf_net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c743_A0 (.DIODE(clknet_1_1__leaf_net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net100_X (.DIODE(clknet_1_1__leaf_net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_S0 (.DIODE(clknet_1_0__leaf_net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_S0 (.DIODE(clknet_1_0__leaf_net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_A1 (.DIODE(clknet_1_0__leaf_net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_c371_S0 (.DIODE(clknet_1_0__leaf_net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net931_X (.DIODE(clknet_1_0__leaf_net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_c212_A2 (.DIODE(clknet_1_1__leaf_net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_A1 (.DIODE(clknet_1_1__leaf_net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_A2 (.DIODE(clknet_1_1__leaf_net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_A1 (.DIODE(clknet_1_1__leaf_net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_output154_A (.DIODE(clknet_1_1__leaf_net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net931_X (.DIODE(clknet_1_1__leaf_net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_S0 (.DIODE(clknet_1_0__leaf_net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_c226_S1 (.DIODE(clknet_1_0__leaf_net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_c240_S1 (.DIODE(clknet_1_0__leaf_net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_S1 (.DIODE(clknet_1_0__leaf_net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_output147_A (.DIODE(clknet_1_0__leaf_net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net924_X (.DIODE(clknet_1_0__leaf_net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_c239_D_N (.DIODE(clknet_1_1__leaf_net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_S0 (.DIODE(clknet_1_1__leaf_net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_c350_S0 (.DIODE(clknet_1_1__leaf_net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_S1 (.DIODE(clknet_1_1__leaf_net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_S1 (.DIODE(clknet_1_1__leaf_net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_A2 (.DIODE(clknet_1_1__leaf_net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net924_X (.DIODE(clknet_1_1__leaf_net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_A2 (.DIODE(clknet_1_0__leaf_net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_A1 (.DIODE(clknet_1_0__leaf_net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_A0 (.DIODE(clknet_1_0__leaf_net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_c346_A0 (.DIODE(clknet_1_0__leaf_net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_A3 (.DIODE(clknet_1_0__leaf_net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_A0 (.DIODE(clknet_1_0__leaf_net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_A3 (.DIODE(clknet_1_0__leaf_net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_A3 (.DIODE(clknet_1_0__leaf_net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net169_X (.DIODE(clknet_1_0__leaf_net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_A1 (.DIODE(clknet_1_1__leaf_net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_c558_A3 (.DIODE(clknet_1_1__leaf_net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_A2 (.DIODE(clknet_1_1__leaf_net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_A0 (.DIODE(clknet_1_1__leaf_net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_c613_A3 (.DIODE(clknet_1_1__leaf_net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net169_X (.DIODE(clknet_1_1__leaf_net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_c218_A1 (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_output152_A (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_c216_A0 (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_A3 (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_A1 (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone6_X (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_A1 (.DIODE(net1048));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_A1 (.DIODE(net1048));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_A2 (.DIODE(net1048));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_A2 (.DIODE(net1048));
 sky130_fd_sc_hd__diode_2 ANTENNA_c399_SET_B (.DIODE(net1048));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone12_X (.DIODE(net1048));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_A0 (.DIODE(net1050));
 sky130_fd_sc_hd__diode_2 ANTENNA_c571_A1 (.DIODE(net1050));
 sky130_fd_sc_hd__diode_2 ANTENNA_c666_RESET_B (.DIODE(net1050));
 sky130_fd_sc_hd__diode_2 ANTENNA_c428_A0 (.DIODE(net1050));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone14_X (.DIODE(net1050));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout192_A (.DIODE(net1051));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_A3 (.DIODE(net1051));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_A0 (.DIODE(net1051));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_A3 (.DIODE(net1051));
 sky130_fd_sc_hd__diode_2 ANTENNA_c724_A0 (.DIODE(net1051));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone15_X (.DIODE(net1051));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A0 (.DIODE(net1053));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_A2 (.DIODE(net1053));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer8_A (.DIODE(net1053));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_A1 (.DIODE(net1053));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone17_X (.DIODE(net1053));
 sky130_fd_sc_hd__diode_2 ANTENNA_c398_B1 (.DIODE(net1054));
 sky130_fd_sc_hd__diode_2 ANTENNA_c228_SCD (.DIODE(net1054));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_S0 (.DIODE(net1054));
 sky130_fd_sc_hd__diode_2 ANTENNA_c234_A2 (.DIODE(net1054));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_A2 (.DIODE(net1054));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone18_X (.DIODE(net1054));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer20_A (.DIODE(net1055));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_A0 (.DIODE(net1055));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer19_X (.DIODE(net1055));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_S0 (.DIODE(net1064));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_A2 (.DIODE(net1064));
 sky130_fd_sc_hd__diode_2 ANTENNA_c366_S0 (.DIODE(net1064));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_S1 (.DIODE(net1064));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_A2 (.DIODE(net1064));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone28_X (.DIODE(net1064));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1_X (.DIODE(net1074));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_C1 (.DIODE(net1074));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_C1 (.DIODE(net1074));
 sky130_fd_sc_hd__diode_2 ANTENNA_c270_D1 (.DIODE(net1074));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_A1 (.DIODE(net1074));
 sky130_fd_sc_hd__diode_2 ANTENNA_c136_A2 (.DIODE(net1074));
 sky130_fd_sc_hd__diode_2 ANTENNA_c134_A2 (.DIODE(net1074));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_A2 (.DIODE(net1074));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_A0 (.DIODE(net1074));
 sky130_fd_sc_hd__diode_2 ANTENNA_c198_A3 (.DIODE(net1074));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_A2 (.DIODE(net1074));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(net556));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(clknet_1_1__leaf_net486));
 sky130_fd_sc_hd__mux4_1 clone1 (.A0(net34),
    .A1(net32),
    .A2(net1062),
    .A3(net790),
    .S0(net31),
    .S1(net995),
    .X(net1075));
 sky130_fd_sc_hd__clkbuf_1 rebuffer2 (.A(net36),
    .X(net1076));
 sky130_fd_sc_hd__mux4_1 clone4 (.A0(net31),
    .A1(net792),
    .A2(net25),
    .A3(net34),
    .S0(net1033),
    .S1(net30),
    .X(net1077));
 sky130_fd_sc_hd__mux4_1 clone5 (.A0(net34),
    .A1(net32),
    .A2(net1062),
    .A3(net790),
    .S0(net31),
    .S1(net995),
    .X(net1078));
 sky130_fd_sc_hd__decap_8 FILLER_0_0_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_67 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_90 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_228 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_59 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_71 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_283 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_24 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_60 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_275 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_20 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_143 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_282 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_451 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_495 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_90 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_308 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_355 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_22 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_595 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_616 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_496 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_87 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_170 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_31 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_423 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_535 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_19 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_422 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_588 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_143 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_340 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_619 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_71 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_499 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_563 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_10 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_395 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_612 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_476 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_143 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_479 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_553 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_284 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_67 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_423 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_535 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_507 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_518 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_116 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_163 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_451 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_527 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_17 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_252 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_518 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_10 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_469 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_172 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_471 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_588 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_366 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_32 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_283 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_5 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_168 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_354 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_103 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_463 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_242 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_227 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_308 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_10 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_5 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_5 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_499 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_617 ();
endmodule
